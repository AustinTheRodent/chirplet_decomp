
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity exponential_rom is
  port
  (
    clk       : in  std_logic;
    address   : in  std_logic_vector(15 downto 0);
    data_out  : out std_logic_vector(31 downto 0)
  );
end entity;

architecture rtl of exponential_rom is

  constant C_DATA_WIDTH  : integer := 32;
  constant C_ADDR_WIDTH  : integer := 16;

  constant RAM_DEPTH :integer := 2**C_ADDR_WIDTH;

  type RAM is array (integer range <>) of std_logic_vector (C_DATA_WIDTH-1 downto 0);
  signal mem : RAM (0 to RAM_DEPTH-1) :=
  (
    x"3F800000",
    x"3F7FE002",
    x"3F7FC008",
    x"3F7FA012",
    x"3F7F8020",
    x"3F7F6032",
    x"3F7F4048",
    x"3F7F2062",
    x"3F7F0080",
    x"3F7EE0A2",
    x"3F7EC0C8",
    x"3F7EA0F2",
    x"3F7E811F",
    x"3F7E6151",
    x"3F7E4187",
    x"3F7E21C1",
    x"3F7E01FF",
    x"3F7DE240",
    x"3F7DC286",
    x"3F7DA2D0",
    x"3F7D831D",
    x"3F7D636F",
    x"3F7D43C5",
    x"3F7D241E",
    x"3F7D047C",
    x"3F7CE4DD",
    x"3F7CC542",
    x"3F7CA5AC",
    x"3F7C8619",
    x"3F7C668A",
    x"3F7C46FF",
    x"3F7C2778",
    x"3F7C07F5",
    x"3F7BE876",
    x"3F7BC8FB",
    x"3F7BA984",
    x"3F7B8A11",
    x"3F7B6AA2",
    x"3F7B4B36",
    x"3F7B2BCF",
    x"3F7B0C6B",
    x"3F7AED0C",
    x"3F7ACDB0",
    x"3F7AAE58",
    x"3F7A8F04",
    x"3F7A6FB4",
    x"3F7A5068",
    x"3F7A3120",
    x"3F7A11DC",
    x"3F79F29C",
    x"3F79D360",
    x"3F79B427",
    x"3F7994F3",
    x"3F7975C2",
    x"3F795695",
    x"3F79376C",
    x"3F791847",
    x"3F78F926",
    x"3F78DA09",
    x"3F78BAF0",
    x"3F789BDA",
    x"3F787CC9",
    x"3F785DBB",
    x"3F783EB1",
    x"3F781FAB",
    x"3F7800A9",
    x"3F77E1AB",
    x"3F77C2B1",
    x"3F77A3BA",
    x"3F7784C8",
    x"3F7765D9",
    x"3F7746EE",
    x"3F772808",
    x"3F770924",
    x"3F76EA45",
    x"3F76CB6A",
    x"3F76AC92",
    x"3F768DBF",
    x"3F766EEF",
    x"3F765023",
    x"3F76315B",
    x"3F761297",
    x"3F75F3D6",
    x"3F75D51A",
    x"3F75B661",
    x"3F7597AC",
    x"3F7578FB",
    x"3F755A4E",
    x"3F753BA5",
    x"3F751CFF",
    x"3F74FE5D",
    x"3F74DFBF",
    x"3F74C125",
    x"3F74A28F",
    x"3F7483FD",
    x"3F74656E",
    x"3F7446E3",
    x"3F74285C",
    x"3F7409D9",
    x"3F73EB5A",
    x"3F73CCDE",
    x"3F73AE67",
    x"3F738FF3",
    x"3F737183",
    x"3F735316",
    x"3F7334AE",
    x"3F731649",
    x"3F72F7E8",
    x"3F72D98B",
    x"3F72BB32",
    x"3F729CDC",
    x"3F727E8B",
    x"3F72603D",
    x"3F7241F3",
    x"3F7223AC",
    x"3F72056A",
    x"3F71E72B",
    x"3F71C8F0",
    x"3F71AAB9",
    x"3F718C85",
    x"3F716E56",
    x"3F71502A",
    x"3F713202",
    x"3F7113DD",
    x"3F70F5BD",
    x"3F70D7A0",
    x"3F70B987",
    x"3F709B71",
    x"3F707D60",
    x"3F705F52",
    x"3F704148",
    x"3F702342",
    x"3F70053F",
    x"3F6FE740",
    x"3F6FC945",
    x"3F6FAB4E",
    x"3F6F8D5B",
    x"3F6F6F6B",
    x"3F6F517F",
    x"3F6F3396",
    x"3F6F15B2",
    x"3F6EF7D1",
    x"3F6ED9F4",
    x"3F6EBC1A",
    x"3F6E9E45",
    x"3F6E8073",
    x"3F6E62A5",
    x"3F6E44DA",
    x"3F6E2714",
    x"3F6E0950",
    x"3F6DEB91",
    x"3F6DCDD6",
    x"3F6DB01E",
    x"3F6D926A",
    x"3F6D74B9",
    x"3F6D570C",
    x"3F6D3963",
    x"3F6D1BBE",
    x"3F6CFE1C",
    x"3F6CE07F",
    x"3F6CC2E4",
    x"3F6CA54E",
    x"3F6C87BB",
    x"3F6C6A2C",
    x"3F6C4CA0",
    x"3F6C2F19",
    x"3F6C1195",
    x"3F6BF414",
    x"3F6BD698",
    x"3F6BB91F",
    x"3F6B9BA9",
    x"3F6B7E38",
    x"3F6B60CA",
    x"3F6B4360",
    x"3F6B25F9",
    x"3F6B0896",
    x"3F6AEB37",
    x"3F6ACDDB",
    x"3F6AB083",
    x"3F6A932F",
    x"3F6A75DF",
    x"3F6A5892",
    x"3F6A3B48",
    x"3F6A1E03",
    x"3F6A00C1",
    x"3F69E383",
    x"3F69C648",
    x"3F69A911",
    x"3F698BDE",
    x"3F696EAE",
    x"3F695182",
    x"3F69345A",
    x"3F691735",
    x"3F68FA14",
    x"3F68DCF6",
    x"3F68BFDD",
    x"3F68A2C7",
    x"3F6885B4",
    x"3F6868A5",
    x"3F684B9A",
    x"3F682E92",
    x"3F68118E",
    x"3F67F48E",
    x"3F67D791",
    x"3F67BA98",
    x"3F679DA2",
    x"3F6780B0",
    x"3F6763C2",
    x"3F6746D8",
    x"3F6729F1",
    x"3F670D0D",
    x"3F66F02D",
    x"3F66D351",
    x"3F66B678",
    x"3F6699A3",
    x"3F667CD2",
    x"3F666004",
    x"3F66433A",
    x"3F662673",
    x"3F6609B0",
    x"3F65ECF1",
    x"3F65D035",
    x"3F65B37D",
    x"3F6596C8",
    x"3F657A17",
    x"3F655D6A",
    x"3F6540C0",
    x"3F65241A",
    x"3F650777",
    x"3F64EAD8",
    x"3F64CE3C",
    x"3F64B1A4",
    x"3F649510",
    x"3F64787F",
    x"3F645BF2",
    x"3F643F68",
    x"3F6422E2",
    x"3F64065F",
    x"3F63E9E0",
    x"3F63CD65",
    x"3F63B0ED",
    x"3F639478",
    x"3F637808",
    x"3F635B9A",
    x"3F633F31",
    x"3F6322CB",
    x"3F630668",
    x"3F62EA09",
    x"3F62CDAE",
    x"3F62B156",
    x"3F629501",
    x"3F6278B0",
    x"3F625C63",
    x"3F624019",
    x"3F6223D3",
    x"3F620790",
    x"3F61EB51",
    x"3F61CF16",
    x"3F61B2DD",
    x"3F6196A9",
    x"3F617A78",
    x"3F615E4A",
    x"3F614220",
    x"3F6125FA",
    x"3F6109D7",
    x"3F60EDB7",
    x"3F60D19B",
    x"3F60B583",
    x"3F60996E",
    x"3F607D5C",
    x"3F60614F",
    x"3F604544",
    x"3F60293D",
    x"3F600D3A",
    x"3F5FF13A",
    x"3F5FD53D",
    x"3F5FB945",
    x"3F5F9D4F",
    x"3F5F815D",
    x"3F5F656F",
    x"3F5F4984",
    x"3F5F2D9C",
    x"3F5F11B8",
    x"3F5EF5D8",
    x"3F5ED9FB",
    x"3F5EBE22",
    x"3F5EA24B",
    x"3F5E8679",
    x"3F5E6AAA",
    x"3F5E4EDE",
    x"3F5E3316",
    x"3F5E1751",
    x"3F5DFB90",
    x"3F5DDFD3",
    x"3F5DC418",
    x"3F5DA862",
    x"3F5D8CAE",
    x"3F5D70FE",
    x"3F5D5552",
    x"3F5D39A9",
    x"3F5D1E04",
    x"3F5D0262",
    x"3F5CE6C3",
    x"3F5CCB28",
    x"3F5CAF90",
    x"3F5C93FC",
    x"3F5C786B",
    x"3F5C5CDE",
    x"3F5C4154",
    x"3F5C25CE",
    x"3F5C0A4B",
    x"3F5BEECB",
    x"3F5BD34F",
    x"3F5BB7D6",
    x"3F5B9C61",
    x"3F5B80EF",
    x"3F5B6581",
    x"3F5B4A16",
    x"3F5B2EAE",
    x"3F5B134A",
    x"3F5AF7E9",
    x"3F5ADC8C",
    x"3F5AC132",
    x"3F5AA5DC",
    x"3F5A8A89",
    x"3F5A6F39",
    x"3F5A53ED",
    x"3F5A38A4",
    x"3F5A1D5F",
    x"3F5A021D",
    x"3F59E6DE",
    x"3F59CBA3",
    x"3F59B06B",
    x"3F599537",
    x"3F597A06",
    x"3F595ED8",
    x"3F5943AE",
    x"3F592888",
    x"3F590D64",
    x"3F58F244",
    x"3F58D728",
    x"3F58BC0E",
    x"3F58A0F9",
    x"3F5885E6",
    x"3F586AD7",
    x"3F584FCB",
    x"3F5834C3",
    x"3F5819BE",
    x"3F57FEBD",
    x"3F57E3BF",
    x"3F57C8C4",
    x"3F57ADCC",
    x"3F5792D8",
    x"3F5777E8",
    x"3F575CFA",
    x"3F574210",
    x"3F57272A",
    x"3F570C47",
    x"3F56F167",
    x"3F56D68A",
    x"3F56BBB1",
    x"3F56A0DB",
    x"3F568609",
    x"3F566B3A",
    x"3F56506E",
    x"3F5635A6",
    x"3F561AE1",
    x"3F56001F",
    x"3F55E561",
    x"3F55CAA6",
    x"3F55AFEE",
    x"3F55953A",
    x"3F557A89",
    x"3F555FDB",
    x"3F554531",
    x"3F552A8A",
    x"3F550FE6",
    x"3F54F546",
    x"3F54DAA9",
    x"3F54C00F",
    x"3F54A579",
    x"3F548AE6",
    x"3F547056",
    x"3F5455CA",
    x"3F543B41",
    x"3F5420BB",
    x"3F540638",
    x"3F53EBB9",
    x"3F53D13D",
    x"3F53B6C5",
    x"3F539C50",
    x"3F5381DE",
    x"3F53676F",
    x"3F534D04",
    x"3F53329C",
    x"3F531837",
    x"3F52FDD6",
    x"3F52E378",
    x"3F52C91D",
    x"3F52AEC6",
    x"3F529471",
    x"3F527A21",
    x"3F525FD3",
    x"3F524589",
    x"3F522B42",
    x"3F5210FE",
    x"3F51F6BD",
    x"3F51DC80",
    x"3F51C246",
    x"3F51A810",
    x"3F518DDC",
    x"3F5173AC",
    x"3F51597F",
    x"3F513F56",
    x"3F51252F",
    x"3F510B0C",
    x"3F50F0ED",
    x"3F50D6D0",
    x"3F50BCB7",
    x"3F50A2A1",
    x"3F50888E",
    x"3F506E7F",
    x"3F505473",
    x"3F503A6A",
    x"3F502064",
    x"3F500662",
    x"3F4FEC62",
    x"3F4FD267",
    x"3F4FB86E",
    x"3F4F9E78",
    x"3F4F8486",
    x"3F4F6A97",
    x"3F4F50AC",
    x"3F4F36C3",
    x"3F4F1CDE",
    x"3F4F02FC",
    x"3F4EE91D",
    x"3F4ECF42",
    x"3F4EB569",
    x"3F4E9B94",
    x"3F4E81C2",
    x"3F4E67F4",
    x"3F4E4E28",
    x"3F4E3460",
    x"3F4E1A9B",
    x"3F4E00DA",
    x"3F4DE71B",
    x"3F4DCD60",
    x"3F4DB3A8",
    x"3F4D99F3",
    x"3F4D8041",
    x"3F4D6693",
    x"3F4D4CE8",
    x"3F4D3340",
    x"3F4D199B",
    x"3F4CFFF9",
    x"3F4CE65B",
    x"3F4CCCC0",
    x"3F4CB328",
    x"3F4C9993",
    x"3F4C8001",
    x"3F4C6673",
    x"3F4C4CE8",
    x"3F4C3360",
    x"3F4C19DB",
    x"3F4C0059",
    x"3F4BE6DB",
    x"3F4BCD5F",
    x"3F4BB3E7",
    x"3F4B9A72",
    x"3F4B8101",
    x"3F4B6792",
    x"3F4B4E27",
    x"3F4B34BF",
    x"3F4B1B5A",
    x"3F4B01F8",
    x"3F4AE899",
    x"3F4ACF3E",
    x"3F4AB5E5",
    x"3F4A9C90",
    x"3F4A833E",
    x"3F4A69EF",
    x"3F4A50A4",
    x"3F4A375B",
    x"3F4A1E16",
    x"3F4A04D4",
    x"3F49EB95",
    x"3F49D259",
    x"3F49B920",
    x"3F499FEB",
    x"3F4986B8",
    x"3F496D89",
    x"3F49545D",
    x"3F493B34",
    x"3F49220E",
    x"3F4908EB",
    x"3F48EFCC",
    x"3F48D6AF",
    x"3F48BD96",
    x"3F48A480",
    x"3F488B6D",
    x"3F48725D",
    x"3F485950",
    x"3F484047",
    x"3F482740",
    x"3F480E3D",
    x"3F47F53D",
    x"3F47DC40",
    x"3F47C346",
    x"3F47AA4F",
    x"3F47915B",
    x"3F47786A",
    x"3F475F7D",
    x"3F474693",
    x"3F472DAB",
    x"3F4714C7",
    x"3F46FBE6",
    x"3F46E308",
    x"3F46CA2D",
    x"3F46B156",
    x"3F469881",
    x"3F467FB0",
    x"3F4666E1",
    x"3F464E16",
    x"3F46354E",
    x"3F461C88",
    x"3F4603C6",
    x"3F45EB08",
    x"3F45D24C",
    x"3F45B993",
    x"3F45A0DD",
    x"3F45882B",
    x"3F456F7B",
    x"3F4556CF",
    x"3F453E26",
    x"3F45257F",
    x"3F450CDC",
    x"3F44F43C",
    x"3F44DB9F",
    x"3F44C305",
    x"3F44AA6E",
    x"3F4491DB",
    x"3F44794A",
    x"3F4460BC",
    x"3F444832",
    x"3F442FAA",
    x"3F441726",
    x"3F43FEA4",
    x"3F43E626",
    x"3F43CDAB",
    x"3F43B533",
    x"3F439CBE",
    x"3F43844C",
    x"3F436BDD",
    x"3F435371",
    x"3F433B08",
    x"3F4322A2",
    x"3F430A3F",
    x"3F42F1DF",
    x"3F42D983",
    x"3F42C129",
    x"3F42A8D2",
    x"3F42907F",
    x"3F42782E",
    x"3F425FE1",
    x"3F424796",
    x"3F422F4F",
    x"3F42170A",
    x"3F41FEC9",
    x"3F41E68B",
    x"3F41CE4F",
    x"3F41B617",
    x"3F419DE2",
    x"3F4185B0",
    x"3F416D80",
    x"3F415554",
    x"3F413D2B",
    x"3F412505",
    x"3F410CE2",
    x"3F40F4C2",
    x"3F40DCA5",
    x"3F40C48B",
    x"3F40AC73",
    x"3F40945F",
    x"3F407C4E",
    x"3F406440",
    x"3F404C35",
    x"3F40342D",
    x"3F401C28",
    x"3F400426",
    x"3F3FEC27",
    x"3F3FD42B",
    x"3F3FBC32",
    x"3F3FA43C",
    x"3F3F8C49",
    x"3F3F7459",
    x"3F3F5C6C",
    x"3F3F4482",
    x"3F3F2C9B",
    x"3F3F14B7",
    x"3F3EFCD6",
    x"3F3EE4F8",
    x"3F3ECD1C",
    x"3F3EB544",
    x"3F3E9D6F",
    x"3F3E859D",
    x"3F3E6DCE",
    x"3F3E5602",
    x"3F3E3E38",
    x"3F3E2672",
    x"3F3E0EAF",
    x"3F3DF6EE",
    x"3F3DDF31",
    x"3F3DC777",
    x"3F3DAFBF",
    x"3F3D980B",
    x"3F3D8059",
    x"3F3D68AA",
    x"3F3D50FF",
    x"3F3D3956",
    x"3F3D21B1",
    x"3F3D0A0E",
    x"3F3CF26E",
    x"3F3CDAD1",
    x"3F3CC337",
    x"3F3CABA0",
    x"3F3C940C",
    x"3F3C7C7B",
    x"3F3C64ED",
    x"3F3C4D62",
    x"3F3C35DA",
    x"3F3C1E55",
    x"3F3C06D2",
    x"3F3BEF53",
    x"3F3BD7D7",
    x"3F3BC05D",
    x"3F3BA8E6",
    x"3F3B9173",
    x"3F3B7A02",
    x"3F3B6294",
    x"3F3B4B29",
    x"3F3B33C2",
    x"3F3B1C5C",
    x"3F3B04FA",
    x"3F3AED9B",
    x"3F3AD63F",
    x"3F3ABEE6",
    x"3F3AA78F",
    x"3F3A903C",
    x"3F3A78EB",
    x"3F3A619E",
    x"3F3A4A53",
    x"3F3A330B",
    x"3F3A1BC6",
    x"3F3A0484",
    x"3F39ED45",
    x"3F39D609",
    x"3F39BECF",
    x"3F39A799",
    x"3F399066",
    x"3F397935",
    x"3F396207",
    x"3F394ADC",
    x"3F3933B5",
    x"3F391C8F",
    x"3F39056D",
    x"3F38EE4E",
    x"3F38D732",
    x"3F38C018",
    x"3F38A902",
    x"3F3891EE",
    x"3F387ADD",
    x"3F3863CF",
    x"3F384CC4",
    x"3F3835BC",
    x"3F381EB7",
    x"3F3807B4",
    x"3F37F0B5",
    x"3F37D9B8",
    x"3F37C2BF",
    x"3F37ABC8",
    x"3F3794D4",
    x"3F377DE2",
    x"3F3766F4",
    x"3F375009",
    x"3F373920",
    x"3F37223A",
    x"3F370B58",
    x"3F36F478",
    x"3F36DD9A",
    x"3F36C6C0",
    x"3F36AFE9",
    x"3F369914",
    x"3F368242",
    x"3F366B74",
    x"3F3654A8",
    x"3F363DDE",
    x"3F362718",
    x"3F361055",
    x"3F35F994",
    x"3F35E2D6",
    x"3F35CC1B",
    x"3F35B563",
    x"3F359EAE",
    x"3F3587FC",
    x"3F35714C",
    x"3F355A9F",
    x"3F3543F5",
    x"3F352D4E",
    x"3F3516AA",
    x"3F350009",
    x"3F34E96A",
    x"3F34D2CE",
    x"3F34BC35",
    x"3F34A59F",
    x"3F348F0C",
    x"3F34787B",
    x"3F3461EE",
    x"3F344B63",
    x"3F3434DB",
    x"3F341E56",
    x"3F3407D3",
    x"3F33F154",
    x"3F33DAD7",
    x"3F33C45D",
    x"3F33ADE6",
    x"3F339772",
    x"3F338100",
    x"3F336A91",
    x"3F335425",
    x"3F333DBC",
    x"3F332756",
    x"3F3310F2",
    x"3F32FA92",
    x"3F32E434",
    x"3F32CDD9",
    x"3F32B780",
    x"3F32A12B",
    x"3F328AD8",
    x"3F327488",
    x"3F325E3B",
    x"3F3247F1",
    x"3F3231A9",
    x"3F321B64",
    x"3F320522",
    x"3F31EEE3",
    x"3F31D8A6",
    x"3F31C26D",
    x"3F31AC36",
    x"3F319602",
    x"3F317FD0",
    x"3F3169A2",
    x"3F315376",
    x"3F313D4D",
    x"3F312727",
    x"3F311103",
    x"3F30FAE2",
    x"3F30E4C4",
    x"3F30CEA9",
    x"3F30B891",
    x"3F30A27B",
    x"3F308C68",
    x"3F307658",
    x"3F30604A",
    x"3F304A40",
    x"3F303438",
    x"3F301E33",
    x"3F300830",
    x"3F2FF231",
    x"3F2FDC34",
    x"3F2FC63A",
    x"3F2FB042",
    x"3F2F9A4E",
    x"3F2F845C",
    x"3F2F6E6C",
    x"3F2F5880",
    x"3F2F4296",
    x"3F2F2CAF",
    x"3F2F16CB",
    x"3F2F00EA",
    x"3F2EEB0B",
    x"3F2ED52F",
    x"3F2EBF56",
    x"3F2EA97F",
    x"3F2E93AB",
    x"3F2E7DDA",
    x"3F2E680C",
    x"3F2E5240",
    x"3F2E3C77",
    x"3F2E26B1",
    x"3F2E10EE",
    x"3F2DFB2D",
    x"3F2DE56F",
    x"3F2DCFB3",
    x"3F2DB9FB",
    x"3F2DA445",
    x"3F2D8E92",
    x"3F2D78E1",
    x"3F2D6334",
    x"3F2D4D89",
    x"3F2D37E0",
    x"3F2D223B",
    x"3F2D0C98",
    x"3F2CF6F7",
    x"3F2CE15A",
    x"3F2CCBBF",
    x"3F2CB627",
    x"3F2CA092",
    x"3F2C8AFF",
    x"3F2C756F",
    x"3F2C5FE1",
    x"3F2C4A57",
    x"3F2C34CF",
    x"3F2C1F4A",
    x"3F2C09C7",
    x"3F2BF447",
    x"3F2BDECA",
    x"3F2BC94F",
    x"3F2BB3D8",
    x"3F2B9E63",
    x"3F2B88F0",
    x"3F2B7380",
    x"3F2B5E13",
    x"3F2B48A9",
    x"3F2B3341",
    x"3F2B1DDC",
    x"3F2B087A",
    x"3F2AF31A",
    x"3F2ADDBD",
    x"3F2AC862",
    x"3F2AB30B",
    x"3F2A9DB6",
    x"3F2A8863",
    x"3F2A7314",
    x"3F2A5DC6",
    x"3F2A487C",
    x"3F2A3334",
    x"3F2A1DEF",
    x"3F2A08AD",
    x"3F29F36D",
    x"3F29DE30",
    x"3F29C8F6",
    x"3F29B3BE",
    x"3F299E89",
    x"3F298956",
    x"3F297426",
    x"3F295EF9",
    x"3F2949CF",
    x"3F2934A7",
    x"3F291F81",
    x"3F290A5F",
    x"3F28F53F",
    x"3F28E021",
    x"3F28CB07",
    x"3F28B5EF",
    x"3F28A0D9",
    x"3F288BC6",
    x"3F2876B6",
    x"3F2861A9",
    x"3F284C9E",
    x"3F283796",
    x"3F282290",
    x"3F280D8D",
    x"3F27F88D",
    x"3F27E38F",
    x"3F27CE94",
    x"3F27B99B",
    x"3F27A4A5",
    x"3F278FB2",
    x"3F277AC1",
    x"3F2765D3",
    x"3F2750E8",
    x"3F273BFF",
    x"3F272719",
    x"3F271235",
    x"3F26FD54",
    x"3F26E876",
    x"3F26D39A",
    x"3F26BEC1",
    x"3F26A9EB",
    x"3F269517",
    x"3F268045",
    x"3F266B77",
    x"3F2656AA",
    x"3F2641E1",
    x"3F262D1A",
    x"3F261856",
    x"3F260394",
    x"3F25EED5",
    x"3F25DA18",
    x"3F25C55E",
    x"3F25B0A7",
    x"3F259BF2",
    x"3F258740",
    x"3F257290",
    x"3F255DE3",
    x"3F254939",
    x"3F253491",
    x"3F251FEC",
    x"3F250B49",
    x"3F24F6A9",
    x"3F24E20B",
    x"3F24CD70",
    x"3F24B8D8",
    x"3F24A442",
    x"3F248FAF",
    x"3F247B1E",
    x"3F246690",
    x"3F245205",
    x"3F243D7C",
    x"3F2428F5",
    x"3F241471",
    x"3F23FFF0",
    x"3F23EB71",
    x"3F23D6F5",
    x"3F23C27C",
    x"3F23AE05",
    x"3F239990",
    x"3F23851E",
    x"3F2370AF",
    x"3F235C42",
    x"3F2347D8",
    x"3F233370",
    x"3F231F0B",
    x"3F230AA8",
    x"3F22F648",
    x"3F22E1EB",
    x"3F22CD90",
    x"3F22B937",
    x"3F22A4E1",
    x"3F22908E",
    x"3F227C3D",
    x"3F2267EF",
    x"3F2253A3",
    x"3F223F5A",
    x"3F222B13",
    x"3F2216CF",
    x"3F22028E",
    x"3F21EE4F",
    x"3F21DA12",
    x"3F21C5D8",
    x"3F21B1A1",
    x"3F219D6C",
    x"3F218939",
    x"3F217509",
    x"3F2160DC",
    x"3F214CB1",
    x"3F213889",
    x"3F212463",
    x"3F211040",
    x"3F20FC1F",
    x"3F20E801",
    x"3F20D3E5",
    x"3F20BFCC",
    x"3F20ABB5",
    x"3F2097A1",
    x"3F20838F",
    x"3F206F80",
    x"3F205B73",
    x"3F204769",
    x"3F203361",
    x"3F201F5C",
    x"3F200B5A",
    x"3F1FF759",
    x"3F1FE35C",
    x"3F1FCF61",
    x"3F1FBB68",
    x"3F1FA772",
    x"3F1F937E",
    x"3F1F7F8D",
    x"3F1F6B9E",
    x"3F1F57B2",
    x"3F1F43C8",
    x"3F1F2FE1",
    x"3F1F1BFC",
    x"3F1F081A",
    x"3F1EF43A",
    x"3F1EE05D",
    x"3F1ECC82",
    x"3F1EB8AA",
    x"3F1EA4D4",
    x"3F1E9101",
    x"3F1E7D30",
    x"3F1E6961",
    x"3F1E5595",
    x"3F1E41CC",
    x"3F1E2E05",
    x"3F1E1A40",
    x"3F1E067E",
    x"3F1DF2BF",
    x"3F1DDF02",
    x"3F1DCB47",
    x"3F1DB78F",
    x"3F1DA3D9",
    x"3F1D9026",
    x"3F1D7C75",
    x"3F1D68C7",
    x"3F1D551B",
    x"3F1D4172",
    x"3F1D2DCB",
    x"3F1D1A26",
    x"3F1D0684",
    x"3F1CF2E4",
    x"3F1CDF47",
    x"3F1CCBAD",
    x"3F1CB814",
    x"3F1CA47F",
    x"3F1C90EB",
    x"3F1C7D5A",
    x"3F1C69CC",
    x"3F1C5640",
    x"3F1C42B6",
    x"3F1C2F2F",
    x"3F1C1BAB",
    x"3F1C0828",
    x"3F1BF4A9",
    x"3F1BE12B",
    x"3F1BCDB0",
    x"3F1BBA38",
    x"3F1BA6C2",
    x"3F1B934E",
    x"3F1B7FDD",
    x"3F1B6C6E",
    x"3F1B5902",
    x"3F1B4598",
    x"3F1B3230",
    x"3F1B1ECB",
    x"3F1B0B69",
    x"3F1AF808",
    x"3F1AE4AB",
    x"3F1AD14F",
    x"3F1ABDF6",
    x"3F1AAAA0",
    x"3F1A974C",
    x"3F1A83FA",
    x"3F1A70AB",
    x"3F1A5D5E",
    x"3F1A4A13",
    x"3F1A36CB",
    x"3F1A2386",
    x"3F1A1042",
    x"3F19FD02",
    x"3F19E9C3",
    x"3F19D687",
    x"3F19C34E",
    x"3F19B016",
    x"3F199CE2",
    x"3F1989AF",
    x"3F19767F",
    x"3F196351",
    x"3F195026",
    x"3F193CFD",
    x"3F1929D7",
    x"3F1916B3",
    x"3F190391",
    x"3F18F072",
    x"3F18DD55",
    x"3F18CA3B",
    x"3F18B723",
    x"3F18A40D",
    x"3F1890FA",
    x"3F187DE9",
    x"3F186ADA",
    x"3F1857CE",
    x"3F1844C4",
    x"3F1831BD",
    x"3F181EB8",
    x"3F180BB5",
    x"3F17F8B5",
    x"3F17E5B7",
    x"3F17D2BB",
    x"3F17BFC2",
    x"3F17ACCC",
    x"3F1799D7",
    x"3F1786E5",
    x"3F1773F5",
    x"3F176108",
    x"3F174E1D",
    x"3F173B35",
    x"3F17284E",
    x"3F17156A",
    x"3F170289",
    x"3F16EFAA",
    x"3F16DCCD",
    x"3F16C9F3",
    x"3F16B71B",
    x"3F16A445",
    x"3F169171",
    x"3F167EA0",
    x"3F166BD2",
    x"3F165906",
    x"3F16463C",
    x"3F163374",
    x"3F1620AF",
    x"3F160DEC",
    x"3F15FB2B",
    x"3F15E86D",
    x"3F15D5B1",
    x"3F15C2F8",
    x"3F15B040",
    x"3F159D8C",
    x"3F158AD9",
    x"3F157829",
    x"3F15657B",
    x"3F1552CF",
    x"3F154026",
    x"3F152D7F",
    x"3F151ADB",
    x"3F150839",
    x"3F14F599",
    x"3F14E2FB",
    x"3F14D060",
    x"3F14BDC7",
    x"3F14AB31",
    x"3F14989C",
    x"3F14860A",
    x"3F14737B",
    x"3F1460EE",
    x"3F144E63",
    x"3F143BDA",
    x"3F142954",
    x"3F1416D0",
    x"3F14044E",
    x"3F13F1CF",
    x"3F13DF52",
    x"3F13CCD7",
    x"3F13BA5E",
    x"3F13A7E8",
    x"3F139574",
    x"3F138303",
    x"3F137094",
    x"3F135E27",
    x"3F134BBC",
    x"3F133954",
    x"3F1326EE",
    x"3F13148A",
    x"3F130229",
    x"3F12EFC9",
    x"3F12DD6D",
    x"3F12CB12",
    x"3F12B8BA",
    x"3F12A664",
    x"3F129410",
    x"3F1281BF",
    x"3F126F70",
    x"3F125D23",
    x"3F124AD9",
    x"3F123890",
    x"3F12264A",
    x"3F121407",
    x"3F1201C5",
    x"3F11EF86",
    x"3F11DD4A",
    x"3F11CB0F",
    x"3F11B8D7",
    x"3F11A6A1",
    x"3F11946D",
    x"3F11823C",
    x"3F11700D",
    x"3F115DE0",
    x"3F114BB5",
    x"3F11398D",
    x"3F112767",
    x"3F111543",
    x"3F110321",
    x"3F10F102",
    x"3F10DEE5",
    x"3F10CCCA",
    x"3F10BAB2",
    x"3F10A89C",
    x"3F109688",
    x"3F108476",
    x"3F107267",
    x"3F106059",
    x"3F104E4F",
    x"3F103C46",
    x"3F102A3F",
    x"3F10183B",
    x"3F100639",
    x"3F0FF43A",
    x"3F0FE23C",
    x"3F0FD041",
    x"3F0FBE48",
    x"3F0FAC52",
    x"3F0F9A5D",
    x"3F0F886B",
    x"3F0F767B",
    x"3F0F648D",
    x"3F0F52A2",
    x"3F0F40B9",
    x"3F0F2ED2",
    x"3F0F1CED",
    x"3F0F0B0B",
    x"3F0EF92A",
    x"3F0EE74C",
    x"3F0ED570",
    x"3F0EC397",
    x"3F0EB1C0",
    x"3F0E9FEA",
    x"3F0E8E18",
    x"3F0E7C47",
    x"3F0E6A79",
    x"3F0E58AC",
    x"3F0E46E2",
    x"3F0E351B",
    x"3F0E2355",
    x"3F0E1192",
    x"3F0DFFD1",
    x"3F0DEE12",
    x"3F0DDC55",
    x"3F0DCA9B",
    x"3F0DB8E3",
    x"3F0DA72D",
    x"3F0D9579",
    x"3F0D83C7",
    x"3F0D7218",
    x"3F0D606B",
    x"3F0D4EC0",
    x"3F0D3D17",
    x"3F0D2B70",
    x"3F0D19CC",
    x"3F0D082A",
    x"3F0CF68A",
    x"3F0CE4EC",
    x"3F0CD351",
    x"3F0CC1B8",
    x"3F0CB020",
    x"3F0C9E8B",
    x"3F0C8CF9",
    x"3F0C7B68",
    x"3F0C69DA",
    x"3F0C584E",
    x"3F0C46C4",
    x"3F0C353C",
    x"3F0C23B7",
    x"3F0C1233",
    x"3F0C00B2",
    x"3F0BEF33",
    x"3F0BDDB6",
    x"3F0BCC3C",
    x"3F0BBAC3",
    x"3F0BA94D",
    x"3F0B97D9",
    x"3F0B8667",
    x"3F0B74F7",
    x"3F0B638A",
    x"3F0B521E",
    x"3F0B40B5",
    x"3F0B2F4E",
    x"3F0B1DE9",
    x"3F0B0C87",
    x"3F0AFB26",
    x"3F0AE9C8",
    x"3F0AD86C",
    x"3F0AC712",
    x"3F0AB5BA",
    x"3F0AA464",
    x"3F0A9311",
    x"3F0A81C0",
    x"3F0A7070",
    x"3F0A5F23",
    x"3F0A4DD9",
    x"3F0A3C90",
    x"3F0A2B49",
    x"3F0A1A05",
    x"3F0A08C3",
    x"3F09F783",
    x"3F09E645",
    x"3F09D509",
    x"3F09C3D0",
    x"3F09B298",
    x"3F09A163",
    x"3F099030",
    x"3F097EFF",
    x"3F096DD0",
    x"3F095CA4",
    x"3F094B79",
    x"3F093A51",
    x"3F09292B",
    x"3F091807",
    x"3F0906E5",
    x"3F08F5C5",
    x"3F08E4A7",
    x"3F08D38C",
    x"3F08C272",
    x"3F08B15B",
    x"3F08A046",
    x"3F088F33",
    x"3F087E22",
    x"3F086D13",
    x"3F085C07",
    x"3F084AFC",
    x"3F0839F4",
    x"3F0828EE",
    x"3F0817EA",
    x"3F0806E8",
    x"3F07F5E8",
    x"3F07E4EA",
    x"3F07D3EF",
    x"3F07C2F5",
    x"3F07B1FE",
    x"3F07A109",
    x"3F079016",
    x"3F077F25",
    x"3F076E36",
    x"3F075D49",
    x"3F074C5F",
    x"3F073B76",
    x"3F072A90",
    x"3F0719AC",
    x"3F0708CA",
    x"3F06F7E9",
    x"3F06E70C",
    x"3F06D630",
    x"3F06C556",
    x"3F06B47E",
    x"3F06A3A9",
    x"3F0692D5",
    x"3F068204",
    x"3F067135",
    x"3F066068",
    x"3F064F9D",
    x"3F063ED4",
    x"3F062E0D",
    x"3F061D48",
    x"3F060C86",
    x"3F05FBC5",
    x"3F05EB07",
    x"3F05DA4B",
    x"3F05C990",
    x"3F05B8D8",
    x"3F05A822",
    x"3F05976E",
    x"3F0586BC",
    x"3F05760C",
    x"3F05655F",
    x"3F0554B3",
    x"3F05440A",
    x"3F053362",
    x"3F0522BD",
    x"3F051219",
    x"3F050178",
    x"3F04F0D9",
    x"3F04E03C",
    x"3F04CFA1",
    x"3F04BF08",
    x"3F04AE71",
    x"3F049DDC",
    x"3F048D4A",
    x"3F047CB9",
    x"3F046C2B",
    x"3F045B9E",
    x"3F044B14",
    x"3F043A8B",
    x"3F042A05",
    x"3F041981",
    x"3F0408FF",
    x"3F03F87F",
    x"3F03E801",
    x"3F03D785",
    x"3F03C70B",
    x"3F03B693",
    x"3F03A61D",
    x"3F0395A9",
    x"3F038538",
    x"3F0374C8",
    x"3F03645A",
    x"3F0353EF",
    x"3F034385",
    x"3F03331E",
    x"3F0322B9",
    x"3F031255",
    x"3F0301F4",
    x"3F02F195",
    x"3F02E138",
    x"3F02D0DD",
    x"3F02C083",
    x"3F02B02C",
    x"3F029FD7",
    x"3F028F84",
    x"3F027F34",
    x"3F026EE5",
    x"3F025E98",
    x"3F024E4D",
    x"3F023E04",
    x"3F022DBE",
    x"3F021D79",
    x"3F020D36",
    x"3F01FCF5",
    x"3F01ECB7",
    x"3F01DC7A",
    x"3F01CC40",
    x"3F01BC07",
    x"3F01ABD1",
    x"3F019B9C",
    x"3F018B6A",
    x"3F017B39",
    x"3F016B0B",
    x"3F015ADF",
    x"3F014AB4",
    x"3F013A8C",
    x"3F012A66",
    x"3F011A41",
    x"3F010A1F",
    x"3F00F9FF",
    x"3F00E9E1",
    x"3F00D9C4",
    x"3F00C9AA",
    x"3F00B992",
    x"3F00A97C",
    x"3F009968",
    x"3F008955",
    x"3F007945",
    x"3F006937",
    x"3F00592B",
    x"3F004921",
    x"3F003919",
    x"3F002913",
    x"3F00190E",
    x"3F00090C",
    x"3EFFF218",
    x"3EFFD21C",
    x"3EFFB224",
    x"3EFF9230",
    x"3EFF723F",
    x"3EFF5253",
    x"3EFF326B",
    x"3EFF1286",
    x"3EFEF2A6",
    x"3EFED2CA",
    x"3EFEB2F1",
    x"3EFE931D",
    x"3EFE734D",
    x"3EFE5380",
    x"3EFE33B8",
    x"3EFE13F3",
    x"3EFDF433",
    x"3EFDD476",
    x"3EFDB4BE",
    x"3EFD9509",
    x"3EFD7558",
    x"3EFD55AC",
    x"3EFD3603",
    x"3EFD165E",
    x"3EFCF6BD",
    x"3EFCD720",
    x"3EFCB788",
    x"3EFC97F3",
    x"3EFC7862",
    x"3EFC58D4",
    x"3EFC394B",
    x"3EFC19C6",
    x"3EFBFA45",
    x"3EFBDAC8",
    x"3EFBBB4E",
    x"3EFB9BD9",
    x"3EFB7C67",
    x"3EFB5CFA",
    x"3EFB3D90",
    x"3EFB1E2A",
    x"3EFAFEC8",
    x"3EFADF6B",
    x"3EFAC011",
    x"3EFAA0BB",
    x"3EFA8168",
    x"3EFA621A",
    x"3EFA42D0",
    x"3EFA238A",
    x"3EFA0447",
    x"3EF9E508",
    x"3EF9C5CE",
    x"3EF9A697",
    x"3EF98764",
    x"3EF96835",
    x"3EF9490A",
    x"3EF929E3",
    x"3EF90AC0",
    x"3EF8EBA0",
    x"3EF8CC85",
    x"3EF8AD6D",
    x"3EF88E59",
    x"3EF86F49",
    x"3EF8503D",
    x"3EF83135",
    x"3EF81231",
    x"3EF7F331",
    x"3EF7D434",
    x"3EF7B53C",
    x"3EF79647",
    x"3EF77756",
    x"3EF75869",
    x"3EF73980",
    x"3EF71A9B",
    x"3EF6FBB9",
    x"3EF6DCDC",
    x"3EF6BE02",
    x"3EF69F2C",
    x"3EF6805A",
    x"3EF6618C",
    x"3EF642C2",
    x"3EF623FC",
    x"3EF60539",
    x"3EF5E67A",
    x"3EF5C7BF",
    x"3EF5A908",
    x"3EF58A55",
    x"3EF56BA6",
    x"3EF54CFA",
    x"3EF52E53",
    x"3EF50FAF",
    x"3EF4F10F",
    x"3EF4D272",
    x"3EF4B3DA",
    x"3EF49545",
    x"3EF476B5",
    x"3EF45828",
    x"3EF4399F",
    x"3EF41B19",
    x"3EF3FC98",
    x"3EF3DE1A",
    x"3EF3BFA0",
    x"3EF3A12A",
    x"3EF382B8",
    x"3EF3644A",
    x"3EF345DF",
    x"3EF32778",
    x"3EF30915",
    x"3EF2EAB6",
    x"3EF2CC5A",
    x"3EF2AE03",
    x"3EF28FAF",
    x"3EF2715F",
    x"3EF25313",
    x"3EF234CA",
    x"3EF21685",
    x"3EF1F845",
    x"3EF1DA07",
    x"3EF1BBCE",
    x"3EF19D98",
    x"3EF17F67",
    x"3EF16139",
    x"3EF1430E",
    x"3EF124E8",
    x"3EF106C5",
    x"3EF0E8A6",
    x"3EF0CA8B",
    x"3EF0AC73",
    x"3EF08E60",
    x"3EF07050",
    x"3EF05244",
    x"3EF0343B",
    x"3EF01637",
    x"3EEFF836",
    x"3EEFDA39",
    x"3EEFBC3F",
    x"3EEF9E4A",
    x"3EEF8058",
    x"3EEF6269",
    x"3EEF447F",
    x"3EEF2698",
    x"3EEF08B5",
    x"3EEEEAD6",
    x"3EEECCFB",
    x"3EEEAF23",
    x"3EEE914F",
    x"3EEE737F",
    x"3EEE55B2",
    x"3EEE37E9",
    x"3EEE1A24",
    x"3EEDFC63",
    x"3EEDDEA5",
    x"3EEDC0EB",
    x"3EEDA335",
    x"3EED8582",
    x"3EED67D3",
    x"3EED4A28",
    x"3EED2C81",
    x"3EED0EDD",
    x"3EECF13D",
    x"3EECD3A1",
    x"3EECB608",
    x"3EEC9873",
    x"3EEC7AE2",
    x"3EEC5D55",
    x"3EEC3FCB",
    x"3EEC2245",
    x"3EEC04C2",
    x"3EEBE743",
    x"3EEBC9C8",
    x"3EEBAC51",
    x"3EEB8EDD",
    x"3EEB716D",
    x"3EEB5401",
    x"3EEB3698",
    x"3EEB1933",
    x"3EEAFBD2",
    x"3EEADE74",
    x"3EEAC11A",
    x"3EEAA3C4",
    x"3EEA8671",
    x"3EEA6922",
    x"3EEA4BD7",
    x"3EEA2E8F",
    x"3EEA114B",
    x"3EE9F40B",
    x"3EE9D6CE",
    x"3EE9B995",
    x"3EE99C60",
    x"3EE97F2E",
    x"3EE96200",
    x"3EE944D6",
    x"3EE927AF",
    x"3EE90A8C",
    x"3EE8ED6C",
    x"3EE8D051",
    x"3EE8B338",
    x"3EE89624",
    x"3EE87913",
    x"3EE85C05",
    x"3EE83EFC",
    x"3EE821F6",
    x"3EE804F3",
    x"3EE7E7F4",
    x"3EE7CAF9",
    x"3EE7AE02",
    x"3EE7910E",
    x"3EE7741D",
    x"3EE75731",
    x"3EE73A48",
    x"3EE71D62",
    x"3EE70080",
    x"3EE6E3A2",
    x"3EE6C6C7",
    x"3EE6A9F0",
    x"3EE68D1D",
    x"3EE6704D",
    x"3EE65381",
    x"3EE636B8",
    x"3EE619F3",
    x"3EE5FD32",
    x"3EE5E074",
    x"3EE5C3BA",
    x"3EE5A703",
    x"3EE58A50",
    x"3EE56DA0",
    x"3EE550F4",
    x"3EE5344C",
    x"3EE517A7",
    x"3EE4FB06",
    x"3EE4DE69",
    x"3EE4C1CF",
    x"3EE4A538",
    x"3EE488A5",
    x"3EE46C16",
    x"3EE44F8A",
    x"3EE43302",
    x"3EE4167E",
    x"3EE3F9FD",
    x"3EE3DD7F",
    x"3EE3C105",
    x"3EE3A48F",
    x"3EE3881C",
    x"3EE36BAD",
    x"3EE34F41",
    x"3EE332D9",
    x"3EE31674",
    x"3EE2FA13",
    x"3EE2DDB6",
    x"3EE2C15C",
    x"3EE2A506",
    x"3EE288B3",
    x"3EE26C63",
    x"3EE25018",
    x"3EE233CF",
    x"3EE2178B",
    x"3EE1FB49",
    x"3EE1DF0C",
    x"3EE1C2D2",
    x"3EE1A69B",
    x"3EE18A68",
    x"3EE16E38",
    x"3EE1520C",
    x"3EE135E4",
    x"3EE119BF",
    x"3EE0FD9E",
    x"3EE0E180",
    x"3EE0C565",
    x"3EE0A94E",
    x"3EE08D3B",
    x"3EE0712B",
    x"3EE0551F",
    x"3EE03916",
    x"3EE01D10",
    x"3EE0010E",
    x"3EDFE510",
    x"3EDFC915",
    x"3EDFAD1E",
    x"3EDF912A",
    x"3EDF7539",
    x"3EDF594D",
    x"3EDF3D63",
    x"3EDF217D",
    x"3EDF059B",
    x"3EDEE9BC",
    x"3EDECDE0",
    x"3EDEB208",
    x"3EDE9634",
    x"3EDE7A63",
    x"3EDE5E95",
    x"3EDE42CB",
    x"3EDE2704",
    x"3EDE0B41",
    x"3EDDEF82",
    x"3EDDD3C5",
    x"3EDDB80D",
    x"3EDD9C57",
    x"3EDD80A6",
    x"3EDD64F7",
    x"3EDD494C",
    x"3EDD2DA5",
    x"3EDD1201",
    x"3EDCF660",
    x"3EDCDAC3",
    x"3EDCBF2A",
    x"3EDCA394",
    x"3EDC8801",
    x"3EDC6C72",
    x"3EDC50E6",
    x"3EDC355D",
    x"3EDC19D8",
    x"3EDBFE57",
    x"3EDBE2D9",
    x"3EDBC75E",
    x"3EDBABE7",
    x"3EDB9073",
    x"3EDB7503",
    x"3EDB5996",
    x"3EDB3E2C",
    x"3EDB22C6",
    x"3EDB0764",
    x"3EDAEC05",
    x"3EDAD0A9",
    x"3EDAB550",
    x"3EDA99FB",
    x"3EDA7EAA",
    x"3EDA635C",
    x"3EDA4811",
    x"3EDA2CCA",
    x"3EDA1186",
    x"3ED9F645",
    x"3ED9DB08",
    x"3ED9BFCF",
    x"3ED9A498",
    x"3ED98965",
    x"3ED96E36",
    x"3ED9530A",
    x"3ED937E1",
    x"3ED91CBC",
    x"3ED9019A",
    x"3ED8E67C",
    x"3ED8CB60",
    x"3ED8B049",
    x"3ED89534",
    x"3ED87A23",
    x"3ED85F16",
    x"3ED8440C",
    x"3ED82905",
    x"3ED80E01",
    x"3ED7F301",
    x"3ED7D805",
    x"3ED7BD0B",
    x"3ED7A215",
    x"3ED78723",
    x"3ED76C34",
    x"3ED75148",
    x"3ED7365F",
    x"3ED71B7A",
    x"3ED70098",
    x"3ED6E5BA",
    x"3ED6CADF",
    x"3ED6B007",
    x"3ED69533",
    x"3ED67A62",
    x"3ED65F94",
    x"3ED644CA",
    x"3ED62A03",
    x"3ED60F40",
    x"3ED5F47F",
    x"3ED5D9C2",
    x"3ED5BF09",
    x"3ED5A453",
    x"3ED589A0",
    x"3ED56EF0",
    x"3ED55444",
    x"3ED5399B",
    x"3ED51EF6",
    x"3ED50453",
    x"3ED4E9B5",
    x"3ED4CF19",
    x"3ED4B481",
    x"3ED499EC",
    x"3ED47F5A",
    x"3ED464CC",
    x"3ED44A41",
    x"3ED42FBA",
    x"3ED41535",
    x"3ED3FAB4",
    x"3ED3E037",
    x"3ED3C5BC",
    x"3ED3AB45",
    x"3ED390D1",
    x"3ED37661",
    x"3ED35BF4",
    x"3ED3418A",
    x"3ED32723",
    x"3ED30CC0",
    x"3ED2F260",
    x"3ED2D804",
    x"3ED2BDAA",
    x"3ED2A354",
    x"3ED28901",
    x"3ED26EB2",
    x"3ED25466",
    x"3ED23A1D",
    x"3ED21FD7",
    x"3ED20595",
    x"3ED1EB56",
    x"3ED1D11A",
    x"3ED1B6E1",
    x"3ED19CAC",
    x"3ED1827A",
    x"3ED1684C",
    x"3ED14E20",
    x"3ED133F8",
    x"3ED119D3",
    x"3ED0FFB2",
    x"3ED0E593",
    x"3ED0CB78",
    x"3ED0B160",
    x"3ED0974C",
    x"3ED07D3B",
    x"3ED0632D",
    x"3ED04922",
    x"3ED02F1A",
    x"3ED01516",
    x"3ECFFB15",
    x"3ECFE117",
    x"3ECFC71D",
    x"3ECFAD26",
    x"3ECF9331",
    x"3ECF7941",
    x"3ECF5F53",
    x"3ECF4569",
    x"3ECF2B82",
    x"3ECF119E",
    x"3ECEF7BD",
    x"3ECEDDE0",
    x"3ECEC406",
    x"3ECEAA2F",
    x"3ECE905B",
    x"3ECE768B",
    x"3ECE5CBE",
    x"3ECE42F4",
    x"3ECE292D",
    x"3ECE0F69",
    x"3ECDF5A9",
    x"3ECDDBEC",
    x"3ECDC232",
    x"3ECDA87C",
    x"3ECD8EC8",
    x"3ECD7518",
    x"3ECD5B6B",
    x"3ECD41C1",
    x"3ECD281A",
    x"3ECD0E77",
    x"3ECCF4D7",
    x"3ECCDB3A",
    x"3ECCC1A0",
    x"3ECCA809",
    x"3ECC8E76",
    x"3ECC74E6",
    x"3ECC5B59",
    x"3ECC41CF",
    x"3ECC2848",
    x"3ECC0EC5",
    x"3ECBF545",
    x"3ECBDBC7",
    x"3ECBC24E",
    x"3ECBA8D7",
    x"3ECB8F63",
    x"3ECB75F3",
    x"3ECB5C86",
    x"3ECB431C",
    x"3ECB29B5",
    x"3ECB1051",
    x"3ECAF6F1",
    x"3ECADD94",
    x"3ECAC43A",
    x"3ECAAAE3",
    x"3ECA918F",
    x"3ECA783E",
    x"3ECA5EF1",
    x"3ECA45A7",
    x"3ECA2C5F",
    x"3ECA131B",
    x"3EC9F9DB",
    x"3EC9E09D",
    x"3EC9C763",
    x"3EC9AE2B",
    x"3EC994F7",
    x"3EC97BC6",
    x"3EC96298",
    x"3EC9496D",
    x"3EC93046",
    x"3EC91721",
    x"3EC8FE00",
    x"3EC8E4E2",
    x"3EC8CBC7",
    x"3EC8B2AF",
    x"3EC8999A",
    x"3EC88088",
    x"3EC8677A",
    x"3EC84E6F",
    x"3EC83566",
    x"3EC81C61",
    x"3EC8035F",
    x"3EC7EA60",
    x"3EC7D165",
    x"3EC7B86C",
    x"3EC79F76",
    x"3EC78684",
    x"3EC76D95",
    x"3EC754A9",
    x"3EC73BC0",
    x"3EC722DA",
    x"3EC709F7",
    x"3EC6F117",
    x"3EC6D83B",
    x"3EC6BF61",
    x"3EC6A68B",
    x"3EC68DB8",
    x"3EC674E7",
    x"3EC65C1A",
    x"3EC64350",
    x"3EC62A8A",
    x"3EC611C6",
    x"3EC5F905",
    x"3EC5E047",
    x"3EC5C78D",
    x"3EC5AED6",
    x"3EC59621",
    x"3EC57D70",
    x"3EC564C2",
    x"3EC54C17",
    x"3EC5336F",
    x"3EC51ACA",
    x"3EC50228",
    x"3EC4E989",
    x"3EC4D0EE",
    x"3EC4B855",
    x"3EC49FC0",
    x"3EC4872D",
    x"3EC46E9E",
    x"3EC45612",
    x"3EC43D88",
    x"3EC42502",
    x"3EC40C7F",
    x"3EC3F3FF",
    x"3EC3DB82",
    x"3EC3C308",
    x"3EC3AA91",
    x"3EC3921E",
    x"3EC379AD",
    x"3EC3613F",
    x"3EC348D5",
    x"3EC3306D",
    x"3EC31808",
    x"3EC2FFA7",
    x"3EC2E749",
    x"3EC2CEED",
    x"3EC2B695",
    x"3EC29E40",
    x"3EC285ED",
    x"3EC26D9E",
    x"3EC25552",
    x"3EC23D09",
    x"3EC224C3",
    x"3EC20C80",
    x"3EC1F43F",
    x"3EC1DC02",
    x"3EC1C3C8",
    x"3EC1AB92",
    x"3EC1935E",
    x"3EC17B2D",
    x"3EC162FF",
    x"3EC14AD4",
    x"3EC132AC",
    x"3EC11A87",
    x"3EC10265",
    x"3EC0EA47",
    x"3EC0D22B",
    x"3EC0BA12",
    x"3EC0A1FC",
    x"3EC089EA",
    x"3EC071DA",
    x"3EC059CD",
    x"3EC041C3",
    x"3EC029BD",
    x"3EC011B9",
    x"3EBFF9B8",
    x"3EBFE1BB",
    x"3EBFC9C0",
    x"3EBFB1C8",
    x"3EBF99D3",
    x"3EBF81E2",
    x"3EBF69F3",
    x"3EBF5207",
    x"3EBF3A1E",
    x"3EBF2239",
    x"3EBF0A56",
    x"3EBEF276",
    x"3EBEDA99",
    x"3EBEC2BF",
    x"3EBEAAE9",
    x"3EBE9315",
    x"3EBE7B44",
    x"3EBE6376",
    x"3EBE4BAB",
    x"3EBE33E3",
    x"3EBE1C1E",
    x"3EBE045C",
    x"3EBDEC9D",
    x"3EBDD4E1",
    x"3EBDBD28",
    x"3EBDA571",
    x"3EBD8DBE",
    x"3EBD760E",
    x"3EBD5E61",
    x"3EBD46B6",
    x"3EBD2F0F",
    x"3EBD176B",
    x"3EBCFFC9",
    x"3EBCE82B",
    x"3EBCD08F",
    x"3EBCB8F7",
    x"3EBCA161",
    x"3EBC89CE",
    x"3EBC723F",
    x"3EBC5AB2",
    x"3EBC4328",
    x"3EBC2BA1",
    x"3EBC141D",
    x"3EBBFC9C",
    x"3EBBE51E",
    x"3EBBCDA3",
    x"3EBBB62A",
    x"3EBB9EB5",
    x"3EBB8743",
    x"3EBB6FD3",
    x"3EBB5867",
    x"3EBB40FD",
    x"3EBB2996",
    x"3EBB1233",
    x"3EBAFAD2",
    x"3EBAE374",
    x"3EBACC19",
    x"3EBAB4C1",
    x"3EBA9D6C",
    x"3EBA861A",
    x"3EBA6ECA",
    x"3EBA577E",
    x"3EBA4034",
    x"3EBA28EE",
    x"3EBA11AA",
    x"3EB9FA69",
    x"3EB9E32C",
    x"3EB9CBF1",
    x"3EB9B4B9",
    x"3EB99D84",
    x"3EB98651",
    x"3EB96F22",
    x"3EB957F5",
    x"3EB940CC",
    x"3EB929A5",
    x"3EB91282",
    x"3EB8FB61",
    x"3EB8E443",
    x"3EB8CD28",
    x"3EB8B60F",
    x"3EB89EFA",
    x"3EB887E8",
    x"3EB870D8",
    x"3EB859CB",
    x"3EB842C2",
    x"3EB82BBB",
    x"3EB814B7",
    x"3EB7FDB6",
    x"3EB7E6B7",
    x"3EB7CFBC",
    x"3EB7B8C3",
    x"3EB7A1CE",
    x"3EB78ADB",
    x"3EB773EB",
    x"3EB75CFE",
    x"3EB74614",
    x"3EB72F2C",
    x"3EB71848",
    x"3EB70166",
    x"3EB6EA88",
    x"3EB6D3AC",
    x"3EB6BCD3",
    x"3EB6A5FD",
    x"3EB68F29",
    x"3EB67859",
    x"3EB6618B",
    x"3EB64AC0",
    x"3EB633F8",
    x"3EB61D33",
    x"3EB60671",
    x"3EB5EFB2",
    x"3EB5D8F5",
    x"3EB5C23B",
    x"3EB5AB85",
    x"3EB594D1",
    x"3EB57E1F",
    x"3EB56771",
    x"3EB550C6",
    x"3EB53A1D",
    x"3EB52377",
    x"3EB50CD4",
    x"3EB4F634",
    x"3EB4DF96",
    x"3EB4C8FC",
    x"3EB4B264",
    x"3EB49BCF",
    x"3EB4853D",
    x"3EB46EAE",
    x"3EB45822",
    x"3EB44198",
    x"3EB42B11",
    x"3EB4148D",
    x"3EB3FE0C",
    x"3EB3E78E",
    x"3EB3D112",
    x"3EB3BA99",
    x"3EB3A424",
    x"3EB38DB0",
    x"3EB37740",
    x"3EB360D3",
    x"3EB34A68",
    x"3EB33400",
    x"3EB31D9B",
    x"3EB30739",
    x"3EB2F0D9",
    x"3EB2DA7C",
    x"3EB2C422",
    x"3EB2ADCB",
    x"3EB29777",
    x"3EB28125",
    x"3EB26AD7",
    x"3EB2548B",
    x"3EB23E42",
    x"3EB227FB",
    x"3EB211B8",
    x"3EB1FB77",
    x"3EB1E539",
    x"3EB1CEFD",
    x"3EB1B8C5",
    x"3EB1A28F",
    x"3EB18C5C",
    x"3EB1762C",
    x"3EB15FFF",
    x"3EB149D4",
    x"3EB133AC",
    x"3EB11D87",
    x"3EB10765",
    x"3EB0F145",
    x"3EB0DB29",
    x"3EB0C50F",
    x"3EB0AEF7",
    x"3EB098E3",
    x"3EB082D1",
    x"3EB06CC2",
    x"3EB056B6",
    x"3EB040AC",
    x"3EB02AA6",
    x"3EB014A2",
    x"3EAFFEA1",
    x"3EAFE8A2",
    x"3EAFD2A6",
    x"3EAFBCAE",
    x"3EAFA6B7",
    x"3EAF90C4",
    x"3EAF7AD3",
    x"3EAF64E5",
    x"3EAF4EFA",
    x"3EAF3911",
    x"3EAF232C",
    x"3EAF0D49",
    x"3EAEF768",
    x"3EAEE18B",
    x"3EAECBB0",
    x"3EAEB5D8",
    x"3EAEA002",
    x"3EAE8A30",
    x"3EAE7460",
    x"3EAE5E93",
    x"3EAE48C8",
    x"3EAE3301",
    x"3EAE1D3C",
    x"3EAE0779",
    x"3EADF1BA",
    x"3EADDBFD",
    x"3EADC643",
    x"3EADB08B",
    x"3EAD9AD7",
    x"3EAD8525",
    x"3EAD6F75",
    x"3EAD59C9",
    x"3EAD441F",
    x"3EAD2E78",
    x"3EAD18D3",
    x"3EAD0331",
    x"3EACED92",
    x"3EACD7F6",
    x"3EACC25C",
    x"3EACACC5",
    x"3EAC9731",
    x"3EAC81A0",
    x"3EAC6C11",
    x"3EAC5685",
    x"3EAC40FB",
    x"3EAC2B74",
    x"3EAC15F0",
    x"3EAC006F",
    x"3EABEAF0",
    x"3EABD574",
    x"3EABBFFB",
    x"3EABAA84",
    x"3EAB9510",
    x"3EAB7F9F",
    x"3EAB6A30",
    x"3EAB54C4",
    x"3EAB3F5B",
    x"3EAB29F4",
    x"3EAB1491",
    x"3EAAFF2F",
    x"3EAAE9D1",
    x"3EAAD475",
    x"3EAABF1C",
    x"3EAAA9C5",
    x"3EAA9471",
    x"3EAA7F20",
    x"3EAA69D1",
    x"3EAA5486",
    x"3EAA3F3C",
    x"3EAA29F6",
    x"3EAA14B2",
    x"3EA9FF71",
    x"3EA9EA32",
    x"3EA9D4F6",
    x"3EA9BFBD",
    x"3EA9AA86",
    x"3EA99552",
    x"3EA98021",
    x"3EA96AF2",
    x"3EA955C6",
    x"3EA9409D",
    x"3EA92B76",
    x"3EA91652",
    x"3EA90130",
    x"3EA8EC11",
    x"3EA8D6F5",
    x"3EA8C1DC",
    x"3EA8ACC5",
    x"3EA897B1",
    x"3EA8829F",
    x"3EA86D90",
    x"3EA85883",
    x"3EA8437A",
    x"3EA82E73",
    x"3EA8196E",
    x"3EA8046C",
    x"3EA7EF6D",
    x"3EA7DA70",
    x"3EA7C576",
    x"3EA7B07F",
    x"3EA79B8A",
    x"3EA78698",
    x"3EA771A9",
    x"3EA75CBC",
    x"3EA747D1",
    x"3EA732EA",
    x"3EA71E05",
    x"3EA70922",
    x"3EA6F442",
    x"3EA6DF65",
    x"3EA6CA8B",
    x"3EA6B5B3",
    x"3EA6A0DD",
    x"3EA68C0A",
    x"3EA6773A",
    x"3EA6626D",
    x"3EA64DA2",
    x"3EA638D9",
    x"3EA62413",
    x"3EA60F50",
    x"3EA5FA90",
    x"3EA5E5D1",
    x"3EA5D116",
    x"3EA5BC5D",
    x"3EA5A7A7",
    x"3EA592F3",
    x"3EA57E42",
    x"3EA56994",
    x"3EA554E8",
    x"3EA5403F",
    x"3EA52B98",
    x"3EA516F4",
    x"3EA50252",
    x"3EA4EDB3",
    x"3EA4D917",
    x"3EA4C47D",
    x"3EA4AFE5",
    x"3EA49B51",
    x"3EA486BF",
    x"3EA4722F",
    x"3EA45DA2",
    x"3EA44918",
    x"3EA43490",
    x"3EA4200B",
    x"3EA40B88",
    x"3EA3F708",
    x"3EA3E28A",
    x"3EA3CE0F",
    x"3EA3B997",
    x"3EA3A521",
    x"3EA390AD",
    x"3EA37C3C",
    x"3EA367CE",
    x"3EA35363",
    x"3EA33EF9",
    x"3EA32A93",
    x"3EA3162F",
    x"3EA301CD",
    x"3EA2ED6E",
    x"3EA2D912",
    x"3EA2C4B8",
    x"3EA2B061",
    x"3EA29C0C",
    x"3EA287BA",
    x"3EA2736A",
    x"3EA25F1D",
    x"3EA24AD2",
    x"3EA2368A",
    x"3EA22245",
    x"3EA20E02",
    x"3EA1F9C1",
    x"3EA1E583",
    x"3EA1D148",
    x"3EA1BD0F",
    x"3EA1A8D8",
    x"3EA194A5",
    x"3EA18073",
    x"3EA16C44",
    x"3EA15818",
    x"3EA143EE",
    x"3EA12FC7",
    x"3EA11BA2",
    x"3EA10780",
    x"3EA0F361",
    x"3EA0DF43",
    x"3EA0CB29",
    x"3EA0B711",
    x"3EA0A2FB",
    x"3EA08EE8",
    x"3EA07AD7",
    x"3EA066C9",
    x"3EA052BE",
    x"3EA03EB5",
    x"3EA02AAE",
    x"3EA016AA",
    x"3EA002A8",
    x"3E9FEEA9",
    x"3E9FDAAD",
    x"3E9FC6B3",
    x"3E9FB2BB",
    x"3E9F9EC6",
    x"3E9F8AD3",
    x"3E9F76E3",
    x"3E9F62F6",
    x"3E9F4F0A",
    x"3E9F3B22",
    x"3E9F273C",
    x"3E9F1358",
    x"3E9EFF77",
    x"3E9EEB98",
    x"3E9ED7BC",
    x"3E9EC3E2",
    x"3E9EB00B",
    x"3E9E9C36",
    x"3E9E8864",
    x"3E9E7494",
    x"3E9E60C7",
    x"3E9E4CFC",
    x"3E9E3933",
    x"3E9E256E",
    x"3E9E11AA",
    x"3E9DFDE9",
    x"3E9DEA2B",
    x"3E9DD66F",
    x"3E9DC2B5",
    x"3E9DAEFE",
    x"3E9D9B49",
    x"3E9D8797",
    x"3E9D73E7",
    x"3E9D603A",
    x"3E9D4C8F",
    x"3E9D38E7",
    x"3E9D2541",
    x"3E9D119E",
    x"3E9CFDFD",
    x"3E9CEA5E",
    x"3E9CD6C2",
    x"3E9CC328",
    x"3E9CAF91",
    x"3E9C9BFD",
    x"3E9C886A",
    x"3E9C74DA",
    x"3E9C614D",
    x"3E9C4DC2",
    x"3E9C3A3A",
    x"3E9C26B4",
    x"3E9C1330",
    x"3E9BFFAF",
    x"3E9BEC30",
    x"3E9BD8B4",
    x"3E9BC53A",
    x"3E9BB1C2",
    x"3E9B9E4D",
    x"3E9B8ADB",
    x"3E9B776B",
    x"3E9B63FD",
    x"3E9B5092",
    x"3E9B3D29",
    x"3E9B29C2",
    x"3E9B165E",
    x"3E9B02FD",
    x"3E9AEF9E",
    x"3E9ADC41",
    x"3E9AC8E7",
    x"3E9AB58F",
    x"3E9AA239",
    x"3E9A8EE6",
    x"3E9A7B95",
    x"3E9A6847",
    x"3E9A54FB",
    x"3E9A41B2",
    x"3E9A2E6B",
    x"3E9A1B26",
    x"3E9A07E4",
    x"3E99F4A4",
    x"3E99E167",
    x"3E99CE2C",
    x"3E99BAF3",
    x"3E99A7BD",
    x"3E99948A",
    x"3E998158",
    x"3E996E29",
    x"3E995AFD",
    x"3E9947D2",
    x"3E9934AB",
    x"3E992185",
    x"3E990E62",
    x"3E98FB42",
    x"3E98E824",
    x"3E98D508",
    x"3E98C1EE",
    x"3E98AED7",
    x"3E989BC3",
    x"3E9888B0",
    x"3E9875A0",
    x"3E986293",
    x"3E984F88",
    x"3E983C7F",
    x"3E982979",
    x"3E981675",
    x"3E980373",
    x"3E97F074",
    x"3E97DD77",
    x"3E97CA7C",
    x"3E97B784",
    x"3E97A48E",
    x"3E97919B",
    x"3E977EAA",
    x"3E976BBB",
    x"3E9758CF",
    x"3E9745E5",
    x"3E9732FE",
    x"3E972018",
    x"3E970D36",
    x"3E96FA55",
    x"3E96E777",
    x"3E96D49B",
    x"3E96C1C2",
    x"3E96AEEB",
    x"3E969C16",
    x"3E968944",
    x"3E967674",
    x"3E9663A6",
    x"3E9650DB",
    x"3E963E12",
    x"3E962B4B",
    x"3E961887",
    x"3E9605C5",
    x"3E95F306",
    x"3E95E049",
    x"3E95CD8E",
    x"3E95BAD5",
    x"3E95A81F",
    x"3E95956B",
    x"3E9582BA",
    x"3E95700A",
    x"3E955D5E",
    x"3E954AB3",
    x"3E95380B",
    x"3E952565",
    x"3E9512C2",
    x"3E950020",
    x"3E94ED82",
    x"3E94DAE5",
    x"3E94C84B",
    x"3E94B5B3",
    x"3E94A31D",
    x"3E94908A",
    x"3E947DF9",
    x"3E946B6B",
    x"3E9458DE",
    x"3E944654",
    x"3E9433CD",
    x"3E942148",
    x"3E940EC5",
    x"3E93FC44",
    x"3E93E9C5",
    x"3E93D749",
    x"3E93C4D0",
    x"3E93B258",
    x"3E939FE3",
    x"3E938D70",
    x"3E937B00",
    x"3E936891",
    x"3E935626",
    x"3E9343BC",
    x"3E933155",
    x"3E931EF0",
    x"3E930C8D",
    x"3E92FA2C",
    x"3E92E7CE",
    x"3E92D572",
    x"3E92C319",
    x"3E92B0C2",
    x"3E929E6D",
    x"3E928C1A",
    x"3E9279CA",
    x"3E92677C",
    x"3E925530",
    x"3E9242E6",
    x"3E92309F",
    x"3E921E5A",
    x"3E920C18",
    x"3E91F9D7",
    x"3E91E799",
    x"3E91D55D",
    x"3E91C324",
    x"3E91B0ED",
    x"3E919EB8",
    x"3E918C85",
    x"3E917A54",
    x"3E916826",
    x"3E9155FA",
    x"3E9143D1",
    x"3E9131A9",
    x"3E911F84",
    x"3E910D62",
    x"3E90FB41",
    x"3E90E923",
    x"3E90D707",
    x"3E90C4ED",
    x"3E90B2D5",
    x"3E90A0C0",
    x"3E908EAD",
    x"3E907C9D",
    x"3E906A8E",
    x"3E905882",
    x"3E904678",
    x"3E903470",
    x"3E90226B",
    x"3E901068",
    x"3E8FFE67",
    x"3E8FEC68",
    x"3E8FDA6C",
    x"3E8FC872",
    x"3E8FB67A",
    x"3E8FA484",
    x"3E8F9290",
    x"3E8F809F",
    x"3E8F6EB0",
    x"3E8F5CC4",
    x"3E8F4AD9",
    x"3E8F38F1",
    x"3E8F270B",
    x"3E8F1527",
    x"3E8F0346",
    x"3E8EF166",
    x"3E8EDF89",
    x"3E8ECDAE",
    x"3E8EBBD6",
    x"3E8EA9FF",
    x"3E8E982B",
    x"3E8E8659",
    x"3E8E748A",
    x"3E8E62BC",
    x"3E8E50F1",
    x"3E8E3F28",
    x"3E8E2D61",
    x"3E8E1B9D",
    x"3E8E09DA",
    x"3E8DF81A",
    x"3E8DE65C",
    x"3E8DD4A1",
    x"3E8DC2E7",
    x"3E8DB130",
    x"3E8D9F7B",
    x"3E8D8DC8",
    x"3E8D7C17",
    x"3E8D6A69",
    x"3E8D58BD",
    x"3E8D4713",
    x"3E8D356B",
    x"3E8D23C5",
    x"3E8D1222",
    x"3E8D0081",
    x"3E8CEEE2",
    x"3E8CDD45",
    x"3E8CCBAB",
    x"3E8CBA12",
    x"3E8CA87C",
    x"3E8C96E8",
    x"3E8C8556",
    x"3E8C73C7",
    x"3E8C6239",
    x"3E8C50AE",
    x"3E8C3F25",
    x"3E8C2D9F",
    x"3E8C1C1A",
    x"3E8C0A97",
    x"3E8BF917",
    x"3E8BE799",
    x"3E8BD61D",
    x"3E8BC4A4",
    x"3E8BB32C",
    x"3E8BA1B7",
    x"3E8B9044",
    x"3E8B7ED3",
    x"3E8B6D64",
    x"3E8B5BF7",
    x"3E8B4A8D",
    x"3E8B3925",
    x"3E8B27BF",
    x"3E8B165B",
    x"3E8B04F9",
    x"3E8AF39A",
    x"3E8AE23C",
    x"3E8AD0E1",
    x"3E8ABF88",
    x"3E8AAE31",
    x"3E8A9CDD",
    x"3E8A8B8A",
    x"3E8A7A3A",
    x"3E8A68EB",
    x"3E8A579F",
    x"3E8A4656",
    x"3E8A350E",
    x"3E8A23C8",
    x"3E8A1285",
    x"3E8A0144",
    x"3E89F005",
    x"3E89DEC8",
    x"3E89CD8D",
    x"3E89BC54",
    x"3E89AB1E",
    x"3E8999E9",
    x"3E8988B7",
    x"3E897787",
    x"3E896659",
    x"3E89552E",
    x"3E894404",
    x"3E8932DD",
    x"3E8921B7",
    x"3E891094",
    x"3E88FF73",
    x"3E88EE54",
    x"3E88DD38",
    x"3E88CC1D",
    x"3E88BB05",
    x"3E88A9EE",
    x"3E8898DA",
    x"3E8887C8",
    x"3E8876B8",
    x"3E8865AA",
    x"3E88549F",
    x"3E884395",
    x"3E88328E",
    x"3E882189",
    x"3E881086",
    x"3E87FF85",
    x"3E87EE86",
    x"3E87DD89",
    x"3E87CC8E",
    x"3E87BB96",
    x"3E87AA9F",
    x"3E8799AB",
    x"3E8788B9",
    x"3E8777C9",
    x"3E8766DB",
    x"3E8755EF",
    x"3E874506",
    x"3E87341E",
    x"3E872338",
    x"3E871255",
    x"3E870174",
    x"3E86F095",
    x"3E86DFB8",
    x"3E86CEDD",
    x"3E86BE04",
    x"3E86AD2D",
    x"3E869C59",
    x"3E868B86",
    x"3E867AB6",
    x"3E8669E8",
    x"3E86591B",
    x"3E864851",
    x"3E863789",
    x"3E8626C3",
    x"3E861600",
    x"3E86053E",
    x"3E85F47E",
    x"3E85E3C1",
    x"3E85D305",
    x"3E85C24C",
    x"3E85B195",
    x"3E85A0E0",
    x"3E85902D",
    x"3E857F7C",
    x"3E856ECD",
    x"3E855E20",
    x"3E854D75",
    x"3E853CCD",
    x"3E852C26",
    x"3E851B81",
    x"3E850ADF",
    x"3E84FA3F",
    x"3E84E9A1",
    x"3E84D904",
    x"3E84C86A",
    x"3E84B7D2",
    x"3E84A73C",
    x"3E8496A8",
    x"3E848617",
    x"3E847587",
    x"3E8464F9",
    x"3E84546E",
    x"3E8443E4",
    x"3E84335D",
    x"3E8422D7",
    x"3E841254",
    x"3E8401D3",
    x"3E83F154",
    x"3E83E0D6",
    x"3E83D05B",
    x"3E83BFE2",
    x"3E83AF6B",
    x"3E839EF6",
    x"3E838E84",
    x"3E837E13",
    x"3E836DA4",
    x"3E835D37",
    x"3E834CCD",
    x"3E833C64",
    x"3E832BFE",
    x"3E831B99",
    x"3E830B37",
    x"3E82FAD6",
    x"3E82EA78",
    x"3E82DA1C",
    x"3E82C9C2",
    x"3E82B969",
    x"3E82A913",
    x"3E8298BF",
    x"3E82886D",
    x"3E82781D",
    x"3E8267CF",
    x"3E825783",
    x"3E824739",
    x"3E8236F1",
    x"3E8226AB",
    x"3E821668",
    x"3E820626",
    x"3E81F5E6",
    x"3E81E5A8",
    x"3E81D56D",
    x"3E81C533",
    x"3E81B4FB",
    x"3E81A4C6",
    x"3E819492",
    x"3E818461",
    x"3E817431",
    x"3E816404",
    x"3E8153D8",
    x"3E8143AF",
    x"3E813387",
    x"3E812362",
    x"3E81133E",
    x"3E81031D",
    x"3E80F2FD",
    x"3E80E2E0",
    x"3E80D2C5",
    x"3E80C2AB",
    x"3E80B294",
    x"3E80A27F",
    x"3E80926B",
    x"3E80825A",
    x"3E80724B",
    x"3E80623E",
    x"3E805232",
    x"3E804229",
    x"3E803222",
    x"3E80221D",
    x"3E801219",
    x"3E800218",
    x"3E7FE431",
    x"3E7FC437",
    x"3E7FA440",
    x"3E7F844E",
    x"3E7F645F",
    x"3E7F4475",
    x"3E7F248E",
    x"3E7F04AC",
    x"3E7EE4CD",
    x"3E7EC4F2",
    x"3E7EA51C",
    x"3E7E8549",
    x"3E7E657A",
    x"3E7E45B0",
    x"3E7E25E9",
    x"3E7E0626",
    x"3E7DE668",
    x"3E7DC6AD",
    x"3E7DA6F6",
    x"3E7D8743",
    x"3E7D6794",
    x"3E7D47E9",
    x"3E7D2842",
    x"3E7D089F",
    x"3E7CE900",
    x"3E7CC965",
    x"3E7CA9CE",
    x"3E7C8A3A",
    x"3E7C6AAB",
    x"3E7C4B20",
    x"3E7C2B98",
    x"3E7C0C15",
    x"3E7BEC95",
    x"3E7BCD1A",
    x"3E7BADA2",
    x"3E7B8E2E",
    x"3E7B6EBE",
    x"3E7B4F52",
    x"3E7B2FEB",
    x"3E7B1087",
    x"3E7AF126",
    x"3E7AD1CA",
    x"3E7AB272",
    x"3E7A931E",
    x"3E7A73CD",
    x"3E7A5481",
    x"3E7A3538",
    x"3E7A15F3",
    x"3E79F6B3",
    x"3E79D776",
    x"3E79B83D",
    x"3E799908",
    x"3E7979D6",
    x"3E795AA9",
    x"3E793B80",
    x"3E791C5A",
    x"3E78FD39",
    x"3E78DE1B",
    x"3E78BF01",
    x"3E789FEB",
    x"3E7880D9",
    x"3E7861CB",
    x"3E7842C1",
    x"3E7823BA",
    x"3E7804B8",
    x"3E77E5B9",
    x"3E77C6BE",
    x"3E77A7C7",
    x"3E7788D4",
    x"3E7769E5",
    x"3E774AFA",
    x"3E772C12",
    x"3E770D2F",
    x"3E76EE4F",
    x"3E76CF73",
    x"3E76B09B",
    x"3E7691C7",
    x"3E7672F7",
    x"3E76542A",
    x"3E763562",
    x"3E76169D",
    x"3E75F7DC",
    x"3E75D91F",
    x"3E75BA66",
    x"3E759BB1",
    x"3E757CFF",
    x"3E755E51",
    x"3E753FA7",
    x"3E752101",
    x"3E75025F",
    x"3E74E3C1",
    x"3E74C526",
    x"3E74A68F",
    x"3E7487FD",
    x"3E74696D",
    x"3E744AE2",
    x"3E742C5B",
    x"3E740DD7",
    x"3E73EF57",
    x"3E73D0DB",
    x"3E73B263",
    x"3E7393EF",
    x"3E73757E",
    x"3E735711",
    x"3E7338A8",
    x"3E731A43",
    x"3E72FBE2",
    x"3E72DD84",
    x"3E72BF2A",
    x"3E72A0D4",
    x"3E728282",
    x"3E726434",
    x"3E7245E9",
    x"3E7227A2",
    x"3E72095F",
    x"3E71EB20",
    x"3E71CCE4",
    x"3E71AEAD",
    x"3E719079",
    x"3E717249",
    x"3E71541C",
    x"3E7135F4",
    x"3E7117CF",
    x"3E70F9AE",
    x"3E70DB90",
    x"3E70BD77",
    x"3E709F61",
    x"3E70814F",
    x"3E706341",
    x"3E704536",
    x"3E70272F",
    x"3E70092C",
    x"3E6FEB2D",
    x"3E6FCD31",
    x"3E6FAF3A",
    x"3E6F9146",
    x"3E6F7355",
    x"3E6F5569",
    x"3E6F3780",
    x"3E6F199B",
    x"3E6EFBBA",
    x"3E6EDDDC",
    x"3E6EC002",
    x"3E6EA22C",
    x"3E6E845A",
    x"3E6E668B",
    x"3E6E48C0",
    x"3E6E2AF9",
    x"3E6E0D35",
    x"3E6DEF75",
    x"3E6DD1B9",
    x"3E6DB401",
    x"3E6D964C",
    x"3E6D789B",
    x"3E6D5AEE",
    x"3E6D3D45",
    x"3E6D1F9F",
    x"3E6D01FD",
    x"3E6CE45E",
    x"3E6CC6C4",
    x"3E6CA92D",
    x"3E6C8B99",
    x"3E6C6E0A",
    x"3E6C507E",
    x"3E6C32F6",
    x"3E6C1571",
    x"3E6BF7F0",
    x"3E6BDA73",
    x"3E6BBCFA",
    x"3E6B9F84",
    x"3E6B8212",
    x"3E6B64A3",
    x"3E6B4739",
    x"3E6B29D2",
    x"3E6B0C6E",
    x"3E6AEF0F",
    x"3E6AD1B2",
    x"3E6AB45A",
    x"3E6A9705",
    x"3E6A79B4",
    x"3E6A5C67",
    x"3E6A3F1D",
    x"3E6A21D7",
    x"3E6A0495",
    x"3E69E756",
    x"3E69CA1B",
    x"3E69ACE3",
    x"3E698FB0",
    x"3E697280",
    x"3E695553",
    x"3E69382A",
    x"3E691B05",
    x"3E68FDE3",
    x"3E68E0C6",
    x"3E68C3AB",
    x"3E68A695",
    x"3E688982",
    x"3E686C72",
    x"3E684F67",
    x"3E68325E",
    x"3E68155A",
    x"3E67F859",
    x"3E67DB5C",
    x"3E67BE62",
    x"3E67A16C",
    x"3E67847A",
    x"3E67678B",
    x"3E674AA0",
    x"3E672DB8",
    x"3E6710D5",
    x"3E66F3F4",
    x"3E66D718",
    x"3E66BA3E",
    x"3E669D69",
    x"3E668097",
    x"3E6663C9",
    x"3E6646FE",
    x"3E662A37",
    x"3E660D74",
    x"3E65F0B4",
    x"3E65D3F7",
    x"3E65B73F",
    x"3E659A8A",
    x"3E657DD8",
    x"3E65612A",
    x"3E654480",
    x"3E6527D9",
    x"3E650B36",
    x"3E64EE96",
    x"3E64D1FA",
    x"3E64B562",
    x"3E6498CD",
    x"3E647C3C",
    x"3E645FAE",
    x"3E644324",
    x"3E64269D",
    x"3E640A1A",
    x"3E63ED9B",
    x"3E63D11F",
    x"3E63B4A6",
    x"3E639831",
    x"3E637BC0",
    x"3E635F52",
    x"3E6342E8",
    x"3E632682",
    x"3E630A1F",
    x"3E62EDBF",
    x"3E62D163",
    x"3E62B50B",
    x"3E6298B6",
    x"3E627C65",
    x"3E626017",
    x"3E6243CD",
    x"3E622786",
    x"3E620B43",
    x"3E61EF03",
    x"3E61D2C7",
    x"3E61B68E",
    x"3E619A59",
    x"3E617E28",
    x"3E6161FA",
    x"3E6145CF",
    x"3E6129A8",
    x"3E610D85",
    x"3E60F165",
    x"3E60D549",
    x"3E60B930",
    x"3E609D1A",
    x"3E608108",
    x"3E6064FA",
    x"3E6048EF",
    x"3E602CE8",
    x"3E6010E4",
    x"3E5FF4E4",
    x"3E5FD8E7",
    x"3E5FBCED",
    x"3E5FA0F8",
    x"3E5F8505",
    x"3E5F6916",
    x"3E5F4D2B",
    x"3E5F3143",
    x"3E5F155F",
    x"3E5EF97E",
    x"3E5EDDA0",
    x"3E5EC1C6",
    x"3E5EA5F0",
    x"3E5E8A1D",
    x"3E5E6E4D",
    x"3E5E5281",
    x"3E5E36B9",
    x"3E5E1AF3",
    x"3E5DFF32",
    x"3E5DE374",
    x"3E5DC7B9",
    x"3E5DAC02",
    x"3E5D904E",
    x"3E5D749E",
    x"3E5D58F1",
    x"3E5D3D47",
    x"3E5D21A2",
    x"3E5D05FF",
    x"3E5CEA60",
    x"3E5CCEC4",
    x"3E5CB32C",
    x"3E5C9798",
    x"3E5C7C06",
    x"3E5C6079",
    x"3E5C44EE",
    x"3E5C2967",
    x"3E5C0DE4",
    x"3E5BF264",
    x"3E5BD6E7",
    x"3E5BBB6E",
    x"3E5B9FF8",
    x"3E5B8486",
    x"3E5B6917",
    x"3E5B4DAC",
    x"3E5B3244",
    x"3E5B16DF",
    x"3E5AFB7E",
    x"3E5AE020",
    x"3E5AC4C6",
    x"3E5AA96F",
    x"3E5A8E1C",
    x"3E5A72CC",
    x"3E5A577F",
    x"3E5A3C36",
    x"3E5A20F0",
    x"3E5A05AE",
    x"3E59EA6F",
    x"3E59CF33",
    x"3E59B3FB",
    x"3E5998C6",
    x"3E597D95",
    x"3E596267",
    x"3E59473C",
    x"3E592C15",
    x"3E5910F1",
    x"3E58F5D1",
    x"3E58DAB4",
    x"3E58BF9A",
    x"3E58A484",
    x"3E588971",
    x"3E586E61",
    x"3E585355",
    x"3E58384C",
    x"3E581D47",
    x"3E580245",
    x"3E57E747",
    x"3E57CC4B",
    x"3E57B153",
    x"3E57965F",
    x"3E577B6E",
    x"3E576080",
    x"3E574596",
    x"3E572AAF",
    x"3E570FCB",
    x"3E56F4EB",
    x"3E56DA0E",
    x"3E56BF34",
    x"3E56A45E",
    x"3E56898B",
    x"3E566EBC",
    x"3E5653F0",
    x"3E563927",
    x"3E561E61",
    x"3E56039F",
    x"3E55E8E0",
    x"3E55CE25",
    x"3E55B36D",
    x"3E5598B8",
    x"3E557E07",
    x"3E556359",
    x"3E5548AE",
    x"3E552E06",
    x"3E551362",
    x"3E54F8C2",
    x"3E54DE24",
    x"3E54C38A",
    x"3E54A8F3",
    x"3E548E60",
    x"3E5473D0",
    x"3E545943",
    x"3E543EB9",
    x"3E542433",
    x"3E5409B0",
    x"3E53EF31",
    x"3E53D4B4",
    x"3E53BA3B",
    x"3E539FC6",
    x"3E538554",
    x"3E536AE5",
    x"3E535079",
    x"3E533610",
    x"3E531BAB",
    x"3E53014A",
    x"3E52E6EB",
    x"3E52CC90",
    x"3E52B238",
    x"3E5297E3",
    x"3E527D92",
    x"3E526344",
    x"3E5248F9",
    x"3E522EB2",
    x"3E52146D",
    x"3E51FA2C",
    x"3E51DFEF",
    x"3E51C5B4",
    x"3E51AB7D",
    x"3E51914A",
    x"3E517719",
    x"3E515CEC",
    x"3E5142C2",
    x"3E51289B",
    x"3E510E78",
    x"3E50F458",
    x"3E50DA3B",
    x"3E50C021",
    x"3E50A60B",
    x"3E508BF7",
    x"3E5071E8",
    x"3E5057DB",
    x"3E503DD2",
    x"3E5023CC",
    x"3E5009C9",
    x"3E4FEFC9",
    x"3E4FD5CD",
    x"3E4FBBD4",
    x"3E4FA1DE",
    x"3E4F87EB",
    x"3E4F6DFC",
    x"3E4F5410",
    x"3E4F3A27",
    x"3E4F2041",
    x"3E4F065F",
    x"3E4EEC80",
    x"3E4ED2A4",
    x"3E4EB8CB",
    x"3E4E9EF5",
    x"3E4E8523",
    x"3E4E6B54",
    x"3E4E5188",
    x"3E4E37C0",
    x"3E4E1DFA",
    x"3E4E0438",
    x"3E4DEA79",
    x"3E4DD0BE",
    x"3E4DB705",
    x"3E4D9D50",
    x"3E4D839E",
    x"3E4D69EF",
    x"3E4D5043",
    x"3E4D369B",
    x"3E4D1CF6",
    x"3E4D0354",
    x"3E4CE9B5",
    x"3E4CD019",
    x"3E4CB681",
    x"3E4C9CEC",
    x"3E4C835A",
    x"3E4C69CB",
    x"3E4C503F",
    x"3E4C36B7",
    x"3E4C1D31",
    x"3E4C03AF",
    x"3E4BEA31",
    x"3E4BD0B5",
    x"3E4BB73C",
    x"3E4B9DC7",
    x"3E4B8455",
    x"3E4B6AE6",
    x"3E4B517A",
    x"3E4B3812",
    x"3E4B1EAC",
    x"3E4B054A",
    x"3E4AEBEB",
    x"3E4AD28F",
    x"3E4AB936",
    x"3E4A9FE1",
    x"3E4A868E",
    x"3E4A6D3F",
    x"3E4A53F3",
    x"3E4A3AAA",
    x"3E4A2164",
    x"3E4A0822",
    x"3E49EEE2",
    x"3E49D5A6",
    x"3E49BC6D",
    x"3E49A337",
    x"3E498A04",
    x"3E4970D4",
    x"3E4957A8",
    x"3E493E7E",
    x"3E492558",
    x"3E490C35",
    x"3E48F315",
    x"3E48D9F8",
    x"3E48C0DF",
    x"3E48A7C8",
    x"3E488EB5",
    x"3E4875A4",
    x"3E485C97",
    x"3E48438D",
    x"3E482A86",
    x"3E481183",
    x"3E47F882",
    x"3E47DF85",
    x"3E47C68A",
    x"3E47AD93",
    x"3E47949F",
    x"3E477BAE",
    x"3E4762C0",
    x"3E4749D5",
    x"3E4730ED",
    x"3E471809",
    x"3E46FF27",
    x"3E46E649",
    x"3E46CD6E",
    x"3E46B496",
    x"3E469BC1",
    x"3E4682EF",
    x"3E466A20",
    x"3E465154",
    x"3E46388C",
    x"3E461FC6",
    x"3E460704",
    x"3E45EE44",
    x"3E45D588",
    x"3E45BCCF",
    x"3E45A419",
    x"3E458B66",
    x"3E4572B6",
    x"3E455A09",
    x"3E45415F",
    x"3E4528B9",
    x"3E451015",
    x"3E44F775",
    x"3E44DED7",
    x"3E44C63D",
    x"3E44ADA6",
    x"3E449512",
    x"3E447C81",
    x"3E4463F3",
    x"3E444B68",
    x"3E4432E0",
    x"3E441A5B",
    x"3E4401D9",
    x"3E43E95A",
    x"3E43D0DF",
    x"3E43B866",
    x"3E439FF1",
    x"3E43877E",
    x"3E436F0F",
    x"3E4356A2",
    x"3E433E39",
    x"3E4325D3",
    x"3E430D70",
    x"3E42F510",
    x"3E42DCB2",
    x"3E42C458",
    x"3E42AC01",
    x"3E4293AD",
    x"3E427B5C",
    x"3E42630F",
    x"3E424AC4",
    x"3E42327C",
    x"3E421A37",
    x"3E4201F5",
    x"3E41E9B7",
    x"3E41D17B",
    x"3E41B942",
    x"3E41A10D",
    x"3E4188DA",
    x"3E4170AA",
    x"3E41587E",
    x"3E414054",
    x"3E41282E",
    x"3E41100A",
    x"3E40F7EA",
    x"3E40DFCC",
    x"3E40C7B2",
    x"3E40AF9A",
    x"3E409786",
    x"3E407F74",
    x"3E406766",
    x"3E404F5B",
    x"3E403752",
    x"3E401F4D",
    x"3E40074A",
    x"3E3FEF4B",
    x"3E3FD74E",
    x"3E3FBF55",
    x"3E3FA75F",
    x"3E3F8F6B",
    x"3E3F777B",
    x"3E3F5F8D",
    x"3E3F47A3",
    x"3E3F2FBB",
    x"3E3F17D7",
    x"3E3EFFF5",
    x"3E3EE817",
    x"3E3ED03B",
    x"3E3EB863",
    x"3E3EA08D",
    x"3E3E88BB",
    x"3E3E70EB",
    x"3E3E591F",
    x"3E3E4155",
    x"3E3E298E",
    x"3E3E11CA",
    x"3E3DFA0A",
    x"3E3DE24C",
    x"3E3DCA91",
    x"3E3DB2D9",
    x"3E3D9B24",
    x"3E3D8373",
    x"3E3D6BC4",
    x"3E3D5418",
    x"3E3D3C6F",
    x"3E3D24C9",
    x"3E3D0D25",
    x"3E3CF585",
    x"3E3CDDE8",
    x"3E3CC64E",
    x"3E3CAEB6",
    x"3E3C9722",
    x"3E3C7F91",
    x"3E3C6802",
    x"3E3C5077",
    x"3E3C38EE",
    x"3E3C2168",
    x"3E3C09E6",
    x"3E3BF266",
    x"3E3BDAE9",
    x"3E3BC36F",
    x"3E3BABF8",
    x"3E3B9484",
    x"3E3B7D13",
    x"3E3B65A5",
    x"3E3B4E3A",
    x"3E3B36D1",
    x"3E3B1F6C",
    x"3E3B080A",
    x"3E3AF0AA",
    x"3E3AD94D",
    x"3E3AC1F4",
    x"3E3AAA9D",
    x"3E3A9349",
    x"3E3A7BF8",
    x"3E3A64AA",
    x"3E3A4D5F",
    x"3E3A3617",
    x"3E3A1ED1",
    x"3E3A078F",
    x"3E39F04F",
    x"3E39D913",
    x"3E39C1D9",
    x"3E39AAA2",
    x"3E39936F",
    x"3E397C3E",
    x"3E39650F",
    x"3E394DE4",
    x"3E3936BC",
    x"3E391F97",
    x"3E390874",
    x"3E38F155",
    x"3E38DA38",
    x"3E38C31E",
    x"3E38AC07",
    x"3E3894F3",
    x"3E387DE2",
    x"3E3866D3",
    x"3E384FC8",
    x"3E3838C0",
    x"3E3821BA",
    x"3E380AB7",
    x"3E37F3B7",
    x"3E37DCBA",
    x"3E37C5C0",
    x"3E37AEC9",
    x"3E3797D4",
    x"3E3780E3",
    x"3E3769F4",
    x"3E375308",
    x"3E373C1F",
    x"3E372539",
    x"3E370E56",
    x"3E36F776",
    x"3E36E098",
    x"3E36C9BE",
    x"3E36B2E6",
    x"3E369C11",
    x"3E36853F",
    x"3E366E6F",
    x"3E3657A3",
    x"3E3640DA",
    x"3E362A13",
    x"3E36134F",
    x"3E35FC8E",
    x"3E35E5D0",
    x"3E35CF15",
    x"3E35B85C",
    x"3E35A1A7",
    x"3E358AF4",
    x"3E357444",
    x"3E355D97",
    x"3E3546EC",
    x"3E353045",
    x"3E3519A0",
    x"3E3502FF",
    x"3E34EC60",
    x"3E34D5C3",
    x"3E34BF2A",
    x"3E34A894",
    x"3E349200",
    x"3E347B6F",
    x"3E3464E1",
    x"3E344E56",
    x"3E3437CE",
    x"3E342148",
    x"3E340AC5",
    x"3E33F445",
    x"3E33DDC8",
    x"3E33C74E",
    x"3E33B0D6",
    x"3E339A62",
    x"3E3383F0",
    x"3E336D81",
    x"3E335714",
    x"3E3340AB",
    x"3E332A44",
    x"3E3313E0",
    x"3E32FD7F",
    x"3E32E721",
    x"3E32D0C5",
    x"3E32BA6D",
    x"3E32A417",
    x"3E328DC4",
    x"3E327773",
    x"3E326126",
    x"3E324ADB",
    x"3E323493",
    x"3E321E4E",
    x"3E32080C",
    x"3E31F1CC",
    x"3E31DB8F",
    x"3E31C555",
    x"3E31AF1E",
    x"3E3198E9",
    x"3E3182B8",
    x"3E316C89",
    x"3E31565C",
    x"3E314033",
    x"3E312A0C",
    x"3E3113E8",
    x"3E30FDC7",
    x"3E30E7A9",
    x"3E30D18D",
    x"3E30BB75",
    x"3E30A55F",
    x"3E308F4B",
    x"3E30793B",
    x"3E30632D",
    x"3E304D22",
    x"3E30371A",
    x"3E302114",
    x"3E300B11",
    x"3E2FF511",
    x"3E2FDF14",
    x"3E2FC91A",
    x"3E2FB322",
    x"3E2F9D2D",
    x"3E2F873B",
    x"3E2F714B",
    x"3E2F5B5E",
    x"3E2F4574",
    x"3E2F2F8D",
    x"3E2F19A8",
    x"3E2F03C7",
    x"3E2EEDE7",
    x"3E2ED80B",
    x"3E2EC231",
    x"3E2EAC5A",
    x"3E2E9686",
    x"3E2E80B5",
    x"3E2E6AE6",
    x"3E2E551A",
    x"3E2E3F51",
    x"3E2E298A",
    x"3E2E13C6",
    x"3E2DFE05",
    x"3E2DE847",
    x"3E2DD28B",
    x"3E2DBCD2",
    x"3E2DA71C",
    x"3E2D9169",
    x"3E2D7BB8",
    x"3E2D660A",
    x"3E2D505E",
    x"3E2D3AB6",
    x"3E2D2510",
    x"3E2D0F6C",
    x"3E2CF9CC",
    x"3E2CE42E",
    x"3E2CCE93",
    x"3E2CB8FA",
    x"3E2CA364",
    x"3E2C8DD1",
    x"3E2C7841",
    x"3E2C62B3",
    x"3E2C4D28",
    x"3E2C37A0",
    x"3E2C221A",
    x"3E2C0C97",
    x"3E2BF717",
    x"3E2BE19A",
    x"3E2BCC1F",
    x"3E2BB6A7",
    x"3E2BA131",
    x"3E2B8BBE",
    x"3E2B764E",
    x"3E2B60E1",
    x"3E2B4B76",
    x"3E2B360E",
    x"3E2B20A8",
    x"3E2B0B46",
    x"3E2AF5E6",
    x"3E2AE088",
    x"3E2ACB2E",
    x"3E2AB5D5",
    x"3E2AA080",
    x"3E2A8B2D",
    x"3E2A75DD",
    x"3E2A6090",
    x"3E2A4B45",
    x"3E2A35FD",
    x"3E2A20B8",
    x"3E2A0B75",
    x"3E29F635",
    x"3E29E0F7",
    x"3E29CBBD",
    x"3E29B684",
    x"3E29A14F",
    x"3E298C1C",
    x"3E2976EC",
    x"3E2961BE",
    x"3E294C93",
    x"3E29376B",
    x"3E292246",
    x"3E290D23",
    x"3E28F802",
    x"3E28E2E5",
    x"3E28CDCA",
    x"3E28B8B1",
    x"3E28A39B",
    x"3E288E88",
    x"3E287978",
    x"3E28646A",
    x"3E284F5F",
    x"3E283A56",
    x"3E282550",
    x"3E28104D",
    x"3E27FB4C",
    x"3E27E64E",
    x"3E27D152",
    x"3E27BC5A",
    x"3E27A763",
    x"3E279270",
    x"3E277D7F",
    x"3E276890",
    x"3E2753A5",
    x"3E273EBB",
    x"3E2729D5",
    x"3E2714F1",
    x"3E270010",
    x"3E26EB31",
    x"3E26D655",
    x"3E26C17B",
    x"3E26ACA4",
    x"3E2697D0",
    x"3E2682FF",
    x"3E266E2F",
    x"3E265963",
    x"3E264499",
    x"3E262FD2",
    x"3E261B0D",
    x"3E26064B",
    x"3E25F18C",
    x"3E25DCCF",
    x"3E25C814",
    x"3E25B35D",
    x"3E259EA8",
    x"3E2589F5",
    x"3E257545",
    x"3E256098",
    x"3E254BED",
    x"3E253745",
    x"3E25229F",
    x"3E250DFC",
    x"3E24F95C",
    x"3E24E4BE",
    x"3E24D022",
    x"3E24BB8A",
    x"3E24A6F4",
    x"3E249260",
    x"3E247DCF",
    x"3E246940",
    x"3E2454B5",
    x"3E24402B",
    x"3E242BA5",
    x"3E241720",
    x"3E24029F",
    x"3E23EE20",
    x"3E23D9A3",
    x"3E23C529",
    x"3E23B0B2",
    x"3E239C3D",
    x"3E2387CB",
    x"3E23735B",
    x"3E235EEE",
    x"3E234A83",
    x"3E23361B",
    x"3E2321B6",
    x"3E230D53",
    x"3E22F8F3",
    x"3E22E495",
    x"3E22D039",
    x"3E22BBE1",
    x"3E22A78B",
    x"3E229337",
    x"3E227EE6",
    x"3E226A97",
    x"3E22564B",
    x"3E224202",
    x"3E222DBB",
    x"3E221976",
    x"3E220534",
    x"3E21F0F5",
    x"3E21DCB8",
    x"3E21C87E",
    x"3E21B446",
    x"3E21A011",
    x"3E218BDE",
    x"3E2177AE",
    x"3E216380",
    x"3E214F55",
    x"3E213B2C",
    x"3E212706",
    x"3E2112E2",
    x"3E20FEC1",
    x"3E20EAA3",
    x"3E20D687",
    x"3E20C26D",
    x"3E20AE56",
    x"3E209A41",
    x"3E20862F",
    x"3E207220",
    x"3E205E13",
    x"3E204A08",
    x"3E203600",
    x"3E2021FB",
    x"3E200DF8",
    x"3E1FF9F7",
    x"3E1FE5F9",
    x"3E1FD1FE",
    x"3E1FBE05",
    x"3E1FAA0E",
    x"3E1F961A",
    x"3E1F8229",
    x"3E1F6E3A",
    x"3E1F5A4D",
    x"3E1F4663",
    x"3E1F327C",
    x"3E1F1E97",
    x"3E1F0AB4",
    x"3E1EF6D4",
    x"3E1EE2F6",
    x"3E1ECF1B",
    x"3E1EBB43",
    x"3E1EA76C",
    x"3E1E9399",
    x"3E1E7FC7",
    x"3E1E6BF9",
    x"3E1E582C",
    x"3E1E4463",
    x"3E1E309B",
    x"3E1E1CD7",
    x"3E1E0914",
    x"3E1DF554",
    x"3E1DE197",
    x"3E1DCDDC",
    x"3E1DBA23",
    x"3E1DA66D",
    x"3E1D92BA",
    x"3E1D7F09",
    x"3E1D6B5A",
    x"3E1D57AE",
    x"3E1D4404",
    x"3E1D305D",
    x"3E1D1CB8",
    x"3E1D0916",
    x"3E1CF576",
    x"3E1CE1D8",
    x"3E1CCE3D",
    x"3E1CBAA5",
    x"3E1CA70F",
    x"3E1C937B",
    x"3E1C7FEA",
    x"3E1C6C5B",
    x"3E1C58CF",
    x"3E1C4545",
    x"3E1C31BD",
    x"3E1C1E38",
    x"3E1C0AB6",
    x"3E1BF736",
    x"3E1BE3B8",
    x"3E1BD03D",
    x"3E1BBCC4",
    x"3E1BA94E",
    x"3E1B95DA",
    x"3E1B8268",
    x"3E1B6EF9",
    x"3E1B5B8C",
    x"3E1B4822",
    x"3E1B34BA",
    x"3E1B2155",
    x"3E1B0DF2",
    x"3E1AFA91",
    x"3E1AE733",
    x"3E1AD3D8",
    x"3E1AC07E",
    x"3E1AAD27",
    x"3E1A99D3",
    x"3E1A8681",
    x"3E1A7331",
    x"3E1A5FE4",
    x"3E1A4C99",
    x"3E1A3951",
    x"3E1A260B",
    x"3E1A12C8",
    x"3E19FF86",
    x"3E19EC48",
    x"3E19D90B",
    x"3E19C5D1",
    x"3E19B29A",
    x"3E199F65",
    x"3E198C32",
    x"3E197902",
    x"3E1965D4",
    x"3E1952A8",
    x"3E193F7F",
    x"3E192C58",
    x"3E191934",
    x"3E190612",
    x"3E18F2F3",
    x"3E18DFD5",
    x"3E18CCBB",
    x"3E18B9A2",
    x"3E18A68C",
    x"3E189379",
    x"3E188067",
    x"3E186D58",
    x"3E185A4C",
    x"3E184742",
    x"3E18343A",
    x"3E182135",
    x"3E180E32",
    x"3E17FB31",
    x"3E17E833",
    x"3E17D537",
    x"3E17C23E",
    x"3E17AF47",
    x"3E179C52",
    x"3E178960",
    x"3E177670",
    x"3E176382",
    x"3E175097",
    x"3E173DAE",
    x"3E172AC7",
    x"3E1717E3",
    x"3E170501",
    x"3E16F222",
    x"3E16DF45",
    x"3E16CC6A",
    x"3E16B992",
    x"3E16A6BC",
    x"3E1693E8",
    x"3E168117",
    x"3E166E48",
    x"3E165B7B",
    x"3E1648B1",
    x"3E1635E9",
    x"3E162323",
    x"3E161060",
    x"3E15FD9F",
    x"3E15EAE1",
    x"3E15D825",
    x"3E15C56B",
    x"3E15B2B3",
    x"3E159FFE",
    x"3E158D4B",
    x"3E157A9B",
    x"3E1567ED",
    x"3E155541",
    x"3E154297",
    x"3E152FF0",
    x"3E151D4B",
    x"3E150AA9",
    x"3E14F809",
    x"3E14E56B",
    x"3E14D2CF",
    x"3E14C036",
    x"3E14AD9F",
    x"3E149B0B",
    x"3E148878",
    x"3E1475E9",
    x"3E14635B",
    x"3E1450D0",
    x"3E143E47",
    x"3E142BC0",
    x"3E14193C",
    x"3E1406BA",
    x"3E13F43A",
    x"3E13E1BD",
    x"3E13CF42",
    x"3E13BCC9",
    x"3E13AA52",
    x"3E1397DE",
    x"3E13856D",
    x"3E1372FD",
    x"3E136090",
    x"3E134E25",
    x"3E133BBC",
    x"3E132956",
    x"3E1316F2",
    x"3E130490",
    x"3E12F231",
    x"3E12DFD4",
    x"3E12CD79",
    x"3E12BB20",
    x"3E12A8CA",
    x"3E129676",
    x"3E128424",
    x"3E1271D5",
    x"3E125F88",
    x"3E124D3D",
    x"3E123AF5",
    x"3E1228AE",
    x"3E12166A",
    x"3E120429",
    x"3E11F1E9",
    x"3E11DFAC",
    x"3E11CD71",
    x"3E11BB39",
    x"3E11A903",
    x"3E1196CF",
    x"3E11849D",
    x"3E11726E",
    x"3E116040",
    x"3E114E15",
    x"3E113BED",
    x"3E1129C7",
    x"3E1117A2",
    x"3E110581",
    x"3E10F361",
    x"3E10E144",
    x"3E10CF29",
    x"3E10BD10",
    x"3E10AAF9",
    x"3E1098E5",
    x"3E1086D3",
    x"3E1074C4",
    x"3E1062B6",
    x"3E1050AB",
    x"3E103EA2",
    x"3E102C9B",
    x"3E101A97",
    x"3E100895",
    x"3E0FF695",
    x"3E0FE497",
    x"3E0FD29B",
    x"3E0FC0A2",
    x"3E0FAEAB",
    x"3E0F9CB7",
    x"3E0F8AC4",
    x"3E0F78D4",
    x"3E0F66E6",
    x"3E0F54FA",
    x"3E0F4311",
    x"3E0F3129",
    x"3E0F1F44",
    x"3E0F0D62",
    x"3E0EFB81",
    x"3E0EE9A3",
    x"3E0ED7C7",
    x"3E0EC5ED",
    x"3E0EB415",
    x"3E0EA240",
    x"3E0E906D",
    x"3E0E7E9C",
    x"3E0E6CCD",
    x"3E0E5B00",
    x"3E0E4936",
    x"3E0E376E",
    x"3E0E25A8",
    x"3E0E13E5",
    x"3E0E0223",
    x"3E0DF064",
    x"3E0DDEA7",
    x"3E0DCCEC",
    x"3E0DBB34",
    x"3E0DA97E",
    x"3E0D97CA",
    x"3E0D8618",
    x"3E0D7468",
    x"3E0D62BB",
    x"3E0D510F",
    x"3E0D3F66",
    x"3E0D2DC0",
    x"3E0D1C1B",
    x"3E0D0A79",
    x"3E0CF8D8",
    x"3E0CE73A",
    x"3E0CD59F",
    x"3E0CC405",
    x"3E0CB26E",
    x"3E0CA0D8",
    x"3E0C8F45",
    x"3E0C7DB4",
    x"3E0C6C26",
    x"3E0C5A99",
    x"3E0C490F",
    x"3E0C3787",
    x"3E0C2601",
    x"3E0C147E",
    x"3E0C02FC",
    x"3E0BF17D",
    x"3E0BE000",
    x"3E0BCE85",
    x"3E0BBD0C",
    x"3E0BAB96",
    x"3E0B9A21",
    x"3E0B88AF",
    x"3E0B773F",
    x"3E0B65D1",
    x"3E0B5466",
    x"3E0B42FC",
    x"3E0B3195",
    x"3E0B2030",
    x"3E0B0ECD",
    x"3E0AFD6C",
    x"3E0AEC0E",
    x"3E0ADAB1",
    x"3E0AC957",
    x"3E0AB7FF",
    x"3E0AA6A9",
    x"3E0A9555",
    x"3E0A8404",
    x"3E0A72B4",
    x"3E0A6167",
    x"3E0A501C",
    x"3E0A3ED3",
    x"3E0A2D8C",
    x"3E0A1C47",
    x"3E0A0B05",
    x"3E09F9C5",
    x"3E09E887",
    x"3E09D74B",
    x"3E09C611",
    x"3E09B4D9",
    x"3E09A3A4",
    x"3E099270",
    x"3E09813F",
    x"3E097010",
    x"3E095EE3",
    x"3E094DB8",
    x"3E093C8F",
    x"3E092B69",
    x"3E091A45",
    x"3E090922",
    x"3E08F802",
    x"3E08E6E4",
    x"3E08D5C9",
    x"3E08C4AF",
    x"3E08B397",
    x"3E08A282",
    x"3E08916F",
    x"3E08805E",
    x"3E086F4F",
    x"3E085E42",
    x"3E084D37",
    x"3E083C2F",
    x"3E082B28",
    x"3E081A24",
    x"3E080922",
    x"3E07F821",
    x"3E07E724",
    x"3E07D628",
    x"3E07C52E",
    x"3E07B436",
    x"3E07A341",
    x"3E07924E",
    x"3E07815C",
    x"3E07706D",
    x"3E075F80",
    x"3E074E95",
    x"3E073DAD",
    x"3E072CC6",
    x"3E071BE1",
    x"3E070AFF",
    x"3E06FA1F",
    x"3E06E940",
    x"3E06D864",
    x"3E06C78A",
    x"3E06B6B2",
    x"3E06A5DD",
    x"3E069509",
    x"3E068437",
    x"3E067368",
    x"3E06629B",
    x"3E0651CF",
    x"3E064106",
    x"3E06303F",
    x"3E061F7A",
    x"3E060EB7",
    x"3E05FDF6",
    x"3E05ED38",
    x"3E05DC7B",
    x"3E05CBC1",
    x"3E05BB08",
    x"3E05AA52",
    x"3E05999E",
    x"3E0588EB",
    x"3E05783B",
    x"3E05678D",
    x"3E0556E1",
    x"3E054638",
    x"3E053590",
    x"3E0524EA",
    x"3E051447",
    x"3E0503A5",
    x"3E04F306",
    x"3E04E268",
    x"3E04D1CD",
    x"3E04C134",
    x"3E04B09D",
    x"3E04A008",
    x"3E048F75",
    x"3E047EE4",
    x"3E046E55",
    x"3E045DC8",
    x"3E044D3E",
    x"3E043CB5",
    x"3E042C2E",
    x"3E041BAA",
    x"3E040B28",
    x"3E03FAA7",
    x"3E03EA29",
    x"3E03D9AD",
    x"3E03C932",
    x"3E03B8BA",
    x"3E03A844",
    x"3E0397D0",
    x"3E03875E",
    x"3E0376EE",
    x"3E036681",
    x"3E035615",
    x"3E0345AB",
    x"3E033543",
    x"3E0324DE",
    x"3E03147A",
    x"3E030419",
    x"3E02F3B9",
    x"3E02E35C",
    x"3E02D300",
    x"3E02C2A7",
    x"3E02B250",
    x"3E02A1FA",
    x"3E0291A7",
    x"3E028156",
    x"3E027107",
    x"3E0260BA",
    x"3E02506F",
    x"3E024026",
    x"3E022FDF",
    x"3E021F9A",
    x"3E020F57",
    x"3E01FF16",
    x"3E01EED7",
    x"3E01DE9A",
    x"3E01CE5F",
    x"3E01BE27",
    x"3E01ADF0",
    x"3E019DBB",
    x"3E018D88",
    x"3E017D58",
    x"3E016D29",
    x"3E015CFC",
    x"3E014CD2",
    x"3E013CA9",
    x"3E012C83",
    x"3E011C5E",
    x"3E010C3B",
    x"3E00FC1B",
    x"3E00EBFC",
    x"3E00DBE0",
    x"3E00CBC5",
    x"3E00BBAD",
    x"3E00AB97",
    x"3E009B82",
    x"3E008B70",
    x"3E007B5F",
    x"3E006B51",
    x"3E005B44",
    x"3E004B3A",
    x"3E003B32",
    x"3E002B2B",
    x"3E001B27",
    x"3E000B24",
    x"3DFFF648",
    x"3DFFD64B",
    x"3DFFB653",
    x"3DFF965E",
    x"3DFF766D",
    x"3DFF5680",
    x"3DFF3697",
    x"3DFF16B2",
    x"3DFEF6D2",
    x"3DFED6F5",
    x"3DFEB71C",
    x"3DFE9747",
    x"3DFE7776",
    x"3DFE57A9",
    x"3DFE37E0",
    x"3DFE181B",
    x"3DFDF85A",
    x"3DFDD89D",
    x"3DFDB8E4",
    x"3DFD992F",
    x"3DFD797E",
    x"3DFD59D0",
    x"3DFD3A27",
    x"3DFD1A82",
    x"3DFCFAE1",
    x"3DFCDB43",
    x"3DFCBBAA",
    x"3DFC9C14",
    x"3DFC7C83",
    x"3DFC5CF5",
    x"3DFC3D6C",
    x"3DFC1DE6",
    x"3DFBFE64",
    x"3DFBDEE6",
    x"3DFBBF6C",
    x"3DFB9FF6",
    x"3DFB8084",
    x"3DFB6116",
    x"3DFB41AC",
    x"3DFB2246",
    x"3DFB02E3",
    x"3DFAE385",
    x"3DFAC42B",
    x"3DFAA4D4",
    x"3DFA8581",
    x"3DFA6633",
    x"3DFA46E8",
    x"3DFA27A1",
    x"3DFA085E",
    x"3DF9E91F",
    x"3DF9C9E4",
    x"3DF9AAAC",
    x"3DF98B79",
    x"3DF96C49",
    x"3DF94D1E",
    x"3DF92DF6",
    x"3DF90ED2",
    x"3DF8EFB3",
    x"3DF8D096",
    x"3DF8B17E",
    x"3DF8926A",
    x"3DF8735A",
    x"3DF8544D",
    x"3DF83545",
    x"3DF81640",
    x"3DF7F73F",
    x"3DF7D842",
    x"3DF7B949",
    x"3DF79A54",
    x"3DF77B62",
    x"3DF75C75",
    x"3DF73D8B",
    x"3DF71EA6",
    x"3DF6FFC4",
    x"3DF6E0E6",
    x"3DF6C20B",
    x"3DF6A335",
    x"3DF68463",
    x"3DF66594",
    x"3DF646C9",
    x"3DF62802",
    x"3DF6093F",
    x"3DF5EA80",
    x"3DF5CBC5",
    x"3DF5AD0D",
    x"3DF58E59",
    x"3DF56FAA",
    x"3DF550FD",
    x"3DF53255",
    x"3DF513B1",
    x"3DF4F510",
    x"3DF4D674",
    x"3DF4B7DB",
    x"3DF49946",
    x"3DF47AB4",
    x"3DF45C27",
    x"3DF43D9D",
    x"3DF41F18",
    x"3DF40096",
    x"3DF3E217",
    x"3DF3C39D",
    x"3DF3A527",
    x"3DF386B4",
    x"3DF36845",
    x"3DF349DA",
    x"3DF32B72",
    x"3DF30D0F",
    x"3DF2EEAF",
    x"3DF2D053",
    x"3DF2B1FB",
    x"3DF293A7",
    x"3DF27556",
    x"3DF25709",
    x"3DF238C0",
    x"3DF21A7B",
    x"3DF1FC3A",
    x"3DF1DDFC",
    x"3DF1BFC2",
    x"3DF1A18C",
    x"3DF1835A",
    x"3DF1652B",
    x"3DF14701",
    x"3DF128DA",
    x"3DF10AB6",
    x"3DF0EC97",
    x"3DF0CE7B",
    x"3DF0B063",
    x"3DF0924F",
    x"3DF0743F",
    x"3DF05632",
    x"3DF03829",
    x"3DF01A24",
    x"3DEFFC23",
    x"3DEFDE25",
    x"3DEFC02B",
    x"3DEFA235",
    x"3DEF8443",
    x"3DEF6654",
    x"3DEF4869",
    x"3DEF2A82",
    x"3DEF0C9E",
    x"3DEEEEBF",
    x"3DEED0E3",
    x"3DEEB30A",
    x"3DEE9536",
    x"3DEE7765",
    x"3DEE5998",
    x"3DEE3BCF",
    x"3DEE1E09",
    x"3DEE0047",
    x"3DEDE289",
    x"3DEDC4CF",
    x"3DEDA718",
    x"3DED8965",
    x"3DED6BB5",
    x"3DED4E0A",
    x"3DED3062",
    x"3DED12BE",
    x"3DECF51D",
    x"3DECD780",
    x"3DECB9E7",
    x"3DEC9C52",
    x"3DEC7EC0",
    x"3DEC6132",
    x"3DEC43A8",
    x"3DEC2621",
    x"3DEC089E",
    x"3DEBEB1F",
    x"3DEBCDA4",
    x"3DEBB02C",
    x"3DEB92B8",
    x"3DEB7547",
    x"3DEB57DA",
    x"3DEB3A71",
    x"3DEB1D0C",
    x"3DEAFFAA",
    x"3DEAE24C",
    x"3DEAC4F1",
    x"3DEAA79B",
    x"3DEA8A47",
    x"3DEA6CF8",
    x"3DEA4FAC",
    x"3DEA3264",
    x"3DEA1520",
    x"3DE9F7DF",
    x"3DE9DAA2",
    x"3DE9BD68",
    x"3DE9A032",
    x"3DE98300",
    x"3DE965D2",
    x"3DE948A7",
    x"3DE92B7F",
    x"3DE90E5C",
    x"3DE8F13C",
    x"3DE8D41F",
    x"3DE8B707",
    x"3DE899F2",
    x"3DE87CE0",
    x"3DE85FD2",
    x"3DE842C8",
    x"3DE825C2",
    x"3DE808BF",
    x"3DE7EBC0",
    x"3DE7CEC4",
    x"3DE7B1CC",
    x"3DE794D7",
    x"3DE777E7",
    x"3DE75AF9",
    x"3DE73E10",
    x"3DE7212A",
    x"3DE70448",
    x"3DE6E769",
    x"3DE6CA8E",
    x"3DE6ADB6",
    x"3DE690E2",
    x"3DE67412",
    x"3DE65745",
    x"3DE63A7C",
    x"3DE61DB7",
    x"3DE600F5",
    x"3DE5E436",
    x"3DE5C77C",
    x"3DE5AAC5",
    x"3DE58E11",
    x"3DE57161",
    x"3DE554B5",
    x"3DE5380C",
    x"3DE51B67",
    x"3DE4FEC5",
    x"3DE4E227",
    x"3DE4C58D",
    x"3DE4A8F6",
    x"3DE48C62",
    x"3DE46FD3",
    x"3DE45346",
    x"3DE436BE",
    x"3DE41A39",
    x"3DE3FDB7",
    x"3DE3E139",
    x"3DE3C4BF",
    x"3DE3A848",
    x"3DE38BD5",
    x"3DE36F65",
    x"3DE352F9",
    x"3DE33690",
    x"3DE31A2B",
    x"3DE2FDCA",
    x"3DE2E16C",
    x"3DE2C511",
    x"3DE2A8BB",
    x"3DE28C67",
    x"3DE27017",
    x"3DE253CB",
    x"3DE23782",
    x"3DE21B3D",
    x"3DE1FEFC",
    x"3DE1E2BE",
    x"3DE1C683",
    x"3DE1AA4C",
    x"3DE18E18",
    x"3DE171E8",
    x"3DE155BC",
    x"3DE13993",
    x"3DE11D6E",
    x"3DE1014C",
    x"3DE0E52D",
    x"3DE0C912",
    x"3DE0ACFB",
    x"3DE090E7",
    x"3DE074D7",
    x"3DE058CA",
    x"3DE03CC1",
    x"3DE020BB",
    x"3DE004B8",
    x"3DDFE8BA",
    x"3DDFCCBE",
    x"3DDFB0C6",
    x"3DDF94D2",
    x"3DDF78E1",
    x"3DDF5CF4",
    x"3DDF410A",
    x"3DDF2523",
    x"3DDF0941",
    x"3DDEED61",
    x"3DDED185",
    x"3DDEB5AD",
    x"3DDE99D8",
    x"3DDE7E06",
    x"3DDE6238",
    x"3DDE466E",
    x"3DDE2AA7",
    x"3DDE0EE3",
    x"3DDDF323",
    x"3DDDD766",
    x"3DDDBBAD",
    x"3DDD9FF7",
    x"3DDD8445",
    x"3DDD6896",
    x"3DDD4CEB",
    x"3DDD3143",
    x"3DDD159F",
    x"3DDCF9FE",
    x"3DDCDE60",
    x"3DDCC2C6",
    x"3DDCA72F",
    x"3DDC8B9C",
    x"3DDC700D",
    x"3DDC5480",
    x"3DDC38F7",
    x"3DDC1D72",
    x"3DDC01F0",
    x"3DDBE672",
    x"3DDBCAF6",
    x"3DDBAF7F",
    x"3DDB940B",
    x"3DDB789A",
    x"3DDB5D2C",
    x"3DDB41C3",
    x"3DDB265C",
    x"3DDB0AF9",
    x"3DDAEF99",
    x"3DDAD43D",
    x"3DDAB8E4",
    x"3DDA9D8F",
    x"3DDA823D",
    x"3DDA66EE",
    x"3DDA4BA3",
    x"3DDA305B",
    x"3DDA1517",
    x"3DD9F9D6",
    x"3DD9DE99",
    x"3DD9C35E",
    x"3DD9A828",
    x"3DD98CF4",
    x"3DD971C4",
    x"3DD95698",
    x"3DD93B6F",
    x"3DD92049",
    x"3DD90527",
    x"3DD8EA08",
    x"3DD8CEEC",
    x"3DD8B3D4",
    x"3DD898BF",
    x"3DD87DAE",
    x"3DD862A0",
    x"3DD84795",
    x"3DD82C8E",
    x"3DD8118A",
    x"3DD7F68A",
    x"3DD7DB8C",
    x"3DD7C093",
    x"3DD7A59C",
    x"3DD78AA9",
    x"3DD76FBA",
    x"3DD754CD",
    x"3DD739E4",
    x"3DD71EFF",
    x"3DD7041D",
    x"3DD6E93E",
    x"3DD6CE62",
    x"3DD6B38A",
    x"3DD698B5",
    x"3DD67DE4",
    x"3DD66316",
    x"3DD6484B",
    x"3DD62D84",
    x"3DD612C0",
    x"3DD5F7FF",
    x"3DD5DD42",
    x"3DD5C288",
    x"3DD5A7D1",
    x"3DD58D1E",
    x"3DD5726E",
    x"3DD557C1",
    x"3DD53D18",
    x"3DD52272",
    x"3DD507CF",
    x"3DD4ED30",
    x"3DD4D294",
    x"3DD4B7FC",
    x"3DD49D66",
    x"3DD482D4",
    x"3DD46845",
    x"3DD44DBA",
    x"3DD43332",
    x"3DD418AD",
    x"3DD3FE2C",
    x"3DD3E3AE",
    x"3DD3C933",
    x"3DD3AEBB",
    x"3DD39447",
    x"3DD379D6",
    x"3DD35F69",
    x"3DD344FF",
    x"3DD32A98",
    x"3DD31034",
    x"3DD2F5D4",
    x"3DD2DB76",
    x"3DD2C11D",
    x"3DD2A6C6",
    x"3DD28C73",
    x"3DD27223",
    x"3DD257D6",
    x"3DD23D8D",
    x"3DD22347",
    x"3DD20904",
    x"3DD1EEC5",
    x"3DD1D489",
    x"3DD1BA50",
    x"3DD1A01A",
    x"3DD185E8",
    x"3DD16BB9",
    x"3DD1518D",
    x"3DD13764",
    x"3DD11D3F",
    x"3DD1031D",
    x"3DD0E8FE",
    x"3DD0CEE3",
    x"3DD0B4CA",
    x"3DD09AB5",
    x"3DD080A4",
    x"3DD06695",
    x"3DD04C8A",
    x"3DD03282",
    x"3DD0187D",
    x"3DCFFE7C",
    x"3DCFE47E",
    x"3DCFCA83",
    x"3DCFB08B",
    x"3DCF9697",
    x"3DCF7CA5",
    x"3DCF62B8",
    x"3DCF48CD",
    x"3DCF2EE5",
    x"3DCF1501",
    x"3DCEFB20",
    x"3DCEE142",
    x"3DCEC768",
    x"3DCEAD90",
    x"3DCE93BC",
    x"3DCE79EC",
    x"3DCE601E",
    x"3DCE4653",
    x"3DCE2C8C",
    x"3DCE12C8",
    x"3DCDF908",
    x"3DCDDF4A",
    x"3DCDC590",
    x"3DCDABD9",
    x"3DCD9225",
    x"3DCD7874",
    x"3DCD5EC7",
    x"3DCD451C",
    x"3DCD2B75",
    x"3DCD11D2",
    x"3DCCF831",
    x"3DCCDE94",
    x"3DCCC4F9",
    x"3DCCAB62",
    x"3DCC91CE",
    x"3DCC783E",
    x"3DCC5EB0",
    x"3DCC4526",
    x"3DCC2B9F",
    x"3DCC121B",
    x"3DCBF89B",
    x"3DCBDF1D",
    x"3DCBC5A3",
    x"3DCBAC2C",
    x"3DCB92B8",
    x"3DCB7947",
    x"3DCB5FD9",
    x"3DCB466F",
    x"3DCB2D08",
    x"3DCB13A4",
    x"3DCAFA43",
    x"3DCAE0E5",
    x"3DCAC78B",
    x"3DCAAE33",
    x"3DCA94DF",
    x"3DCA7B8E",
    x"3DCA6240",
    x"3DCA48F6",
    x"3DCA2FAE",
    x"3DCA166A",
    x"3DC9FD28",
    x"3DC9E3EA",
    x"3DC9CAAF",
    x"3DC9B178",
    x"3DC99843",
    x"3DC97F12",
    x"3DC965E3",
    x"3DC94CB8",
    x"3DC93390",
    x"3DC91A6B",
    x"3DC9014A",
    x"3DC8E82B",
    x"3DC8CF0F",
    x"3DC8B5F7",
    x"3DC89CE2",
    x"3DC883D0",
    x"3DC86AC1",
    x"3DC851B5",
    x"3DC838AD",
    x"3DC81FA7",
    x"3DC806A5",
    x"3DC7EDA5",
    x"3DC7D4A9",
    x"3DC7BBB0",
    x"3DC7A2BA",
    x"3DC789C8",
    x"3DC770D8",
    x"3DC757EB",
    x"3DC73F02",
    x"3DC7261C",
    x"3DC70D38",
    x"3DC6F458",
    x"3DC6DB7B",
    x"3DC6C2A1",
    x"3DC6A9CB",
    x"3DC690F7",
    x"3DC67826",
    x"3DC65F59",
    x"3DC6468F",
    x"3DC62DC7",
    x"3DC61503",
    x"3DC5FC42",
    x"3DC5E384",
    x"3DC5CAC9",
    x"3DC5B211",
    x"3DC5995D",
    x"3DC580AB",
    x"3DC567FC",
    x"3DC54F51",
    x"3DC536A9",
    x"3DC51E03",
    x"3DC50561",
    x"3DC4ECC2",
    x"3DC4D426",
    x"3DC4BB8D",
    x"3DC4A2F7",
    x"3DC48A64",
    x"3DC471D4",
    x"3DC45948",
    x"3DC440BE",
    x"3DC42838",
    x"3DC40FB4",
    x"3DC3F734",
    x"3DC3DEB6",
    x"3DC3C63C",
    x"3DC3ADC5",
    x"3DC39551",
    x"3DC37CDF",
    x"3DC36471",
    x"3DC34C06",
    x"3DC3339E",
    x"3DC31B39",
    x"3DC302D8",
    x"3DC2EA79",
    x"3DC2D21D",
    x"3DC2B9C4",
    x"3DC2A16E",
    x"3DC2891C",
    x"3DC270CC",
    x"3DC25880",
    x"3DC24036",
    x"3DC227F0",
    x"3DC20FAC",
    x"3DC1F76C",
    x"3DC1DF2E",
    x"3DC1C6F4",
    x"3DC1AEBC",
    x"3DC19688",
    x"3DC17E57",
    x"3DC16629",
    x"3DC14DFD",
    x"3DC135D5",
    x"3DC11DB0",
    x"3DC1058E",
    x"3DC0ED6E",
    x"3DC0D552",
    x"3DC0BD39",
    x"3DC0A523",
    x"3DC08D10",
    x"3DC07500",
    x"3DC05CF3",
    x"3DC044E8",
    x"3DC02CE1",
    x"3DC014DD",
    x"3DBFFCDC",
    x"3DBFE4DE",
    x"3DBFCCE3",
    x"3DBFB4EB",
    x"3DBF9CF6",
    x"3DBF8504",
    x"3DBF6D14",
    x"3DBF5528",
    x"3DBF3D3F",
    x"3DBF2559",
    x"3DBF0D76",
    x"3DBEF596",
    x"3DBEDDB8",
    x"3DBEC5DE",
    x"3DBEAE07",
    x"3DBE9633",
    x"3DBE7E61",
    x"3DBE6693",
    x"3DBE4EC8",
    x"3DBE36FF",
    x"3DBE1F3A",
    x"3DBE0778",
    x"3DBDEFB8",
    x"3DBDD7FC",
    x"3DBDC042",
    x"3DBDA88C",
    x"3DBD90D8",
    x"3DBD7927",
    x"3DBD617A",
    x"3DBD49CF",
    x"3DBD3227",
    x"3DBD1A82",
    x"3DBD02E1",
    x"3DBCEB42",
    x"3DBCD3A6",
    x"3DBCBC0D",
    x"3DBCA477",
    x"3DBC8CE4",
    x"3DBC7554",
    x"3DBC5DC6",
    x"3DBC463C",
    x"3DBC2EB5",
    x"3DBC1730",
    x"3DBBFFAF",
    x"3DBBE831",
    x"3DBBD0B5",
    x"3DBBB93C",
    x"3DBBA1C7",
    x"3DBB8A54",
    x"3DBB72E4",
    x"3DBB5B77",
    x"3DBB440D",
    x"3DBB2CA6",
    x"3DBB1542",
    x"3DBAFDE1",
    x"3DBAE683",
    x"3DBACF27",
    x"3DBAB7CF",
    x"3DBAA079",
    x"3DBA8927",
    x"3DBA71D7",
    x"3DBA5A8A",
    x"3DBA4340",
    x"3DBA2BF9",
    x"3DBA14B5",
    x"3DB9FD74",
    x"3DB9E636",
    x"3DB9CEFB",
    x"3DB9B7C2",
    x"3DB9A08D",
    x"3DB9895A",
    x"3DB9722A",
    x"3DB95AFE",
    x"3DB943D4",
    x"3DB92CAD",
    x"3DB91588",
    x"3DB8FE67",
    x"3DB8E749",
    x"3DB8D02D",
    x"3DB8B915",
    x"3DB8A1FF",
    x"3DB88AEC",
    x"3DB873DC",
    x"3DB85CCF",
    x"3DB845C5",
    x"3DB82EBE",
    x"3DB817BA",
    x"3DB800B8",
    x"3DB7E9B9",
    x"3DB7D2BE",
    x"3DB7BBC5",
    x"3DB7A4CF",
    x"3DB78DDB",
    x"3DB776EB",
    x"3DB75FFE",
    x"3DB74913",
    x"3DB7322B",
    x"3DB71B47",
    x"3DB70465",
    x"3DB6ED86",
    x"3DB6D6A9",
    x"3DB6BFD0",
    x"3DB6A8F9",
    x"3DB69226",
    x"3DB67B55",
    x"3DB66487",
    x"3DB64DBC",
    x"3DB636F3",
    x"3DB6202E",
    x"3DB6096B",
    x"3DB5F2AC",
    x"3DB5DBEF",
    x"3DB5C535",
    x"3DB5AE7D",
    x"3DB597C9",
    x"3DB58117",
    x"3DB56A69",
    x"3DB553BD",
    x"3DB53D14",
    x"3DB5266E",
    x"3DB50FCA",
    x"3DB4F92A",
    x"3DB4E28C",
    x"3DB4CBF1",
    x"3DB4B559",
    x"3DB49EC4",
    x"3DB48831",
    x"3DB471A2",
    x"3DB45B15",
    x"3DB4448B",
    x"3DB42E04",
    x"3DB4177F",
    x"3DB400FE",
    x"3DB3EA7F",
    x"3DB3D403",
    x"3DB3BD8A",
    x"3DB3A714",
    x"3DB390A0",
    x"3DB37A30",
    x"3DB363C2",
    x"3DB34D57",
    x"3DB336EE",
    x"3DB32089",
    x"3DB30A26",
    x"3DB2F3C6",
    x"3DB2DD69",
    x"3DB2C70F",
    x"3DB2B0B8",
    x"3DB29A63",
    x"3DB28411",
    x"3DB26DC2",
    x"3DB25775",
    x"3DB2412C",
    x"3DB22AE5",
    x"3DB214A1",
    x"3DB1FE60",
    x"3DB1E822",
    x"3DB1D1E6",
    x"3DB1BBAD",
    x"3DB1A577",
    x"3DB18F44",
    x"3DB17913",
    x"3DB162E6",
    x"3DB14CBB",
    x"3DB13692",
    x"3DB1206D",
    x"3DB10A4A",
    x"3DB0F42A",
    x"3DB0DE0D",
    x"3DB0C7F3",
    x"3DB0B1DB",
    x"3DB09BC6",
    x"3DB085B4",
    x"3DB06FA5",
    x"3DB05998",
    x"3DB0438F",
    x"3DB02D87",
    x"3DB01783",
    x"3DB00182",
    x"3DAFEB83",
    x"3DAFD587",
    x"3DAFBF8D",
    x"3DAFA997",
    x"3DAF93A3",
    x"3DAF7DB2",
    x"3DAF67C4",
    x"3DAF51D8",
    x"3DAF3BEF",
    x"3DAF2609",
    x"3DAF1026",
    x"3DAEFA45",
    x"3DAEE467",
    x"3DAECE8C",
    x"3DAEB8B3",
    x"3DAEA2DE",
    x"3DAE8D0B",
    x"3DAE773A",
    x"3DAE616D",
    x"3DAE4BA2",
    x"3DAE35DA",
    x"3DAE2015",
    x"3DAE0A52",
    x"3DADF492",
    x"3DADDED5",
    x"3DADC91A",
    x"3DADB363",
    x"3DAD9DAD",
    x"3DAD87FB",
    x"3DAD724B",
    x"3DAD5C9F",
    x"3DAD46F4",
    x"3DAD314D",
    x"3DAD1BA8",
    x"3DAD0606",
    x"3DACF066",
    x"3DACDACA",
    x"3DACC530",
    x"3DACAF98",
    x"3DAC9A04",
    x"3DAC8472",
    x"3DAC6EE3",
    x"3DAC5956",
    x"3DAC43CC",
    x"3DAC2E45",
    x"3DAC18C1",
    x"3DAC033F",
    x"3DABEDC0",
    x"3DABD844",
    x"3DABC2CA",
    x"3DABAD53",
    x"3DAB97DF",
    x"3DAB826D",
    x"3DAB6CFE",
    x"3DAB5792",
    x"3DAB4228",
    x"3DAB2CC1",
    x"3DAB175D",
    x"3DAB01FB",
    x"3DAAEC9C",
    x"3DAAD740",
    x"3DAAC1E7",
    x"3DAAAC90",
    x"3DAA973C",
    x"3DAA81EA",
    x"3DAA6C9B",
    x"3DAA574F",
    x"3DAA4205",
    x"3DAA2CBE",
    x"3DAA177A",
    x"3DAA0238",
    x"3DA9ECF9",
    x"3DA9D7BD",
    x"3DA9C284",
    x"3DA9AD4D",
    x"3DA99818",
    x"3DA982E7",
    x"3DA96DB7",
    x"3DA9588B",
    x"3DA94361",
    x"3DA92E3A",
    x"3DA91916",
    x"3DA903F4",
    x"3DA8EED5",
    x"3DA8D9B8",
    x"3DA8C49E",
    x"3DA8AF87",
    x"3DA89A72",
    x"3DA88560",
    x"3DA87051",
    x"3DA85B44",
    x"3DA8463A",
    x"3DA83133",
    x"3DA81C2E",
    x"3DA8072C",
    x"3DA7F22C",
    x"3DA7DD2F",
    x"3DA7C835",
    x"3DA7B33D",
    x"3DA79E48",
    x"3DA78956",
    x"3DA77466",
    x"3DA75F79",
    x"3DA74A8E",
    x"3DA735A6",
    x"3DA720C1",
    x"3DA70BDE",
    x"3DA6F6FE",
    x"3DA6E220",
    x"3DA6CD45",
    x"3DA6B86D",
    x"3DA6A397",
    x"3DA68EC4",
    x"3DA679F3",
    x"3DA66525",
    x"3DA6505A",
    x"3DA63B91",
    x"3DA626CB",
    x"3DA61207",
    x"3DA5FD47",
    x"3DA5E888",
    x"3DA5D3CC",
    x"3DA5BF13",
    x"3DA5AA5D",
    x"3DA595A9",
    x"3DA580F7",
    x"3DA56C48",
    x"3DA5579C",
    x"3DA542F2",
    x"3DA52E4B",
    x"3DA519A7",
    x"3DA50505",
    x"3DA4F066",
    x"3DA4DBC9",
    x"3DA4C72F",
    x"3DA4B297",
    x"3DA49E02",
    x"3DA48970",
    x"3DA474E0",
    x"3DA46052",
    x"3DA44BC8",
    x"3DA4373F",
    x"3DA422BA",
    x"3DA40E37",
    x"3DA3F9B6",
    x"3DA3E538",
    x"3DA3D0BD",
    x"3DA3BC44",
    x"3DA3A7CE",
    x"3DA3935A",
    x"3DA37EE9",
    x"3DA36A7A",
    x"3DA3560E",
    x"3DA341A5",
    x"3DA32D3E",
    x"3DA318DA",
    x"3DA30478",
    x"3DA2F019",
    x"3DA2DBBC",
    x"3DA2C762",
    x"3DA2B30A",
    x"3DA29EB5",
    x"3DA28A62",
    x"3DA27612",
    x"3DA261C5",
    x"3DA24D7A",
    x"3DA23931",
    x"3DA224EB",
    x"3DA210A8",
    x"3DA1FC67",
    x"3DA1E829",
    x"3DA1D3ED",
    x"3DA1BFB4",
    x"3DA1AB7D",
    x"3DA19749",
    x"3DA18318",
    x"3DA16EE8",
    x"3DA15ABC",
    x"3DA14692",
    x"3DA1326A",
    x"3DA11E45",
    x"3DA10A23",
    x"3DA0F603",
    x"3DA0E1E5",
    x"3DA0CDCA",
    x"3DA0B9B2",
    x"3DA0A59C",
    x"3DA09188",
    x"3DA07D77",
    x"3DA06969",
    x"3DA0555D",
    x"3DA04154",
    x"3DA02D4D",
    x"3DA01948",
    x"3DA00546",
    x"3D9FF147",
    x"3D9FDD4A",
    x"3D9FC950",
    x"3D9FB558",
    x"3D9FA162",
    x"3D9F8D6F",
    x"3D9F797F",
    x"3D9F6591",
    x"3D9F51A5",
    x"3D9F3DBD",
    x"3D9F29D6",
    x"3D9F15F2",
    x"3D9F0211",
    x"3D9EEE32",
    x"3D9EDA55",
    x"3D9EC67B",
    x"3D9EB2A3",
    x"3D9E9ECE",
    x"3D9E8AFC",
    x"3D9E772C",
    x"3D9E635E",
    x"3D9E4F93",
    x"3D9E3BCA",
    x"3D9E2804",
    x"3D9E1440",
    x"3D9E007F",
    x"3D9DECC0",
    x"3D9DD903",
    x"3D9DC54A",
    x"3D9DB192",
    x"3D9D9DDD",
    x"3D9D8A2B",
    x"3D9D767B",
    x"3D9D62CD",
    x"3D9D4F22",
    x"3D9D3B79",
    x"3D9D27D3",
    x"3D9D142F",
    x"3D9D008E",
    x"3D9CECEF",
    x"3D9CD953",
    x"3D9CC5B9",
    x"3D9CB221",
    x"3D9C9E8C",
    x"3D9C8AFA",
    x"3D9C776A",
    x"3D9C63DC",
    x"3D9C5051",
    x"3D9C3CC8",
    x"3D9C2941",
    x"3D9C15BE",
    x"3D9C023C",
    x"3D9BEEBD",
    x"3D9BDB40",
    x"3D9BC7C6",
    x"3D9BB44E",
    x"3D9BA0D9",
    x"3D9B8D66",
    x"3D9B79F6",
    x"3D9B6688",
    x"3D9B531C",
    x"3D9B3FB3",
    x"3D9B2C4C",
    x"3D9B18E8",
    x"3D9B0586",
    x"3D9AF226",
    x"3D9ADEC9",
    x"3D9ACB6F",
    x"3D9AB817",
    x"3D9AA4C1",
    x"3D9A916D",
    x"3D9A7E1C",
    x"3D9A6ACE",
    x"3D9A5782",
    x"3D9A4438",
    x"3D9A30F1",
    x"3D9A1DAC",
    x"3D9A0A69",
    x"3D99F729",
    x"3D99E3EB",
    x"3D99D0B0",
    x"3D99BD77",
    x"3D99AA41",
    x"3D99970D",
    x"3D9983DB",
    x"3D9970AC",
    x"3D995D7F",
    x"3D994A54",
    x"3D99372C",
    x"3D992407",
    x"3D9910E3",
    x"3D98FDC2",
    x"3D98EAA4",
    x"3D98D788",
    x"3D98C46E",
    x"3D98B157",
    x"3D989E42",
    x"3D988B2F",
    x"3D98781F",
    x"3D986511",
    x"3D985206",
    x"3D983EFC",
    x"3D982BF6",
    x"3D9818F1",
    x"3D9805F0",
    x"3D97F2F0",
    x"3D97DFF3",
    x"3D97CCF8",
    x"3D97BA00",
    x"3D97A709",
    x"3D979416",
    x"3D978124",
    x"3D976E35",
    x"3D975B49",
    x"3D97485F",
    x"3D973577",
    x"3D972291",
    x"3D970FAE",
    x"3D96FCCD",
    x"3D96E9EF",
    x"3D96D713",
    x"3D96C439",
    x"3D96B162",
    x"3D969E8D",
    x"3D968BBA",
    x"3D9678EA",
    x"3D96661C",
    x"3D965350",
    x"3D964087",
    x"3D962DC0",
    x"3D961AFC",
    x"3D96083A",
    x"3D95F57A",
    x"3D95E2BC",
    x"3D95D001",
    x"3D95BD48",
    x"3D95AA92",
    x"3D9597DD",
    x"3D95852C",
    x"3D95727C",
    x"3D955FCF",
    x"3D954D24",
    x"3D953A7C",
    x"3D9527D6",
    x"3D951532",
    x"3D950290",
    x"3D94EFF1",
    x"3D94DD54",
    x"3D94CABA",
    x"3D94B822",
    x"3D94A58C",
    x"3D9492F8",
    x"3D948067",
    x"3D946DD8",
    x"3D945B4C",
    x"3D9448C1",
    x"3D943639",
    x"3D9423B4",
    x"3D941130",
    x"3D93FEAF",
    x"3D93EC31",
    x"3D93D9B4",
    x"3D93C73A",
    x"3D93B4C3",
    x"3D93A24D",
    x"3D938FDA",
    x"3D937D69",
    x"3D936AFB",
    x"3D93588E",
    x"3D934625",
    x"3D9333BD",
    x"3D932158",
    x"3D930EF5",
    x"3D92FC94",
    x"3D92EA35",
    x"3D92D7D9",
    x"3D92C580",
    x"3D92B328",
    x"3D92A0D3",
    x"3D928E80",
    x"3D927C2F",
    x"3D9269E1",
    x"3D925795",
    x"3D92454B",
    x"3D923303",
    x"3D9220BE",
    x"3D920E7B",
    x"3D91FC3A",
    x"3D91E9FC",
    x"3D91D7C0",
    x"3D91C586",
    x"3D91B34F",
    x"3D91A119",
    x"3D918EE6",
    x"3D917CB6",
    x"3D916A87",
    x"3D91585B",
    x"3D914631",
    x"3D913409",
    x"3D9121E4",
    x"3D910FC1",
    x"3D90FDA0",
    x"3D90EB82",
    x"3D90D965",
    x"3D90C74B",
    x"3D90B533",
    x"3D90A31E",
    x"3D90910B",
    x"3D907EFA",
    x"3D906CEB",
    x"3D905ADE",
    x"3D9048D4",
    x"3D9036CC",
    x"3D9024C6",
    x"3D9012C3",
    x"3D9000C2",
    x"3D8FEEC3",
    x"3D8FDCC6",
    x"3D8FCACC",
    x"3D8FB8D3",
    x"3D8FA6DD",
    x"3D8F94EA",
    x"3D8F82F8",
    x"3D8F7109",
    x"3D8F5F1C",
    x"3D8F4D31",
    x"3D8F3B49",
    x"3D8F2962",
    x"3D8F177E",
    x"3D8F059C",
    x"3D8EF3BD",
    x"3D8EE1DF",
    x"3D8ED004",
    x"3D8EBE2B",
    x"3D8EAC55",
    x"3D8E9A80",
    x"3D8E88AE",
    x"3D8E76DE",
    x"3D8E6510",
    x"3D8E5345",
    x"3D8E417C",
    x"3D8E2FB5",
    x"3D8E1DF0",
    x"3D8E0C2D",
    x"3D8DFA6D",
    x"3D8DE8AF",
    x"3D8DD6F3",
    x"3D8DC539",
    x"3D8DB381",
    x"3D8DA1CC",
    x"3D8D9019",
    x"3D8D7E68",
    x"3D8D6CB9",
    x"3D8D5B0D",
    x"3D8D4962",
    x"3D8D37BA",
    x"3D8D2614",
    x"3D8D1471",
    x"3D8D02CF",
    x"3D8CF130",
    x"3D8CDF93",
    x"3D8CCDF8",
    x"3D8CBC60",
    x"3D8CAAC9",
    x"3D8C9935",
    x"3D8C87A3",
    x"3D8C7613",
    x"3D8C6485",
    x"3D8C52FA",
    x"3D8C4171",
    x"3D8C2FE9",
    x"3D8C1E65",
    x"3D8C0CE2",
    x"3D8BFB61",
    x"3D8BE9E3",
    x"3D8BD867",
    x"3D8BC6ED",
    x"3D8BB575",
    x"3D8BA400",
    x"3D8B928C",
    x"3D8B811B",
    x"3D8B6FAC",
    x"3D8B5E3F",
    x"3D8B4CD4",
    x"3D8B3B6C",
    x"3D8B2A05",
    x"3D8B18A1",
    x"3D8B073F",
    x"3D8AF5DF",
    x"3D8AE482",
    x"3D8AD326",
    x"3D8AC1CD",
    x"3D8AB076",
    x"3D8A9F21",
    x"3D8A8DCE",
    x"3D8A7C7D",
    x"3D8A6B2F",
    x"3D8A59E3",
    x"3D8A4899",
    x"3D8A3751",
    x"3D8A260B",
    x"3D8A14C7",
    x"3D8A0386",
    x"3D89F246",
    x"3D89E109",
    x"3D89CFCE",
    x"3D89BE95",
    x"3D89AD5E",
    x"3D899C2A",
    x"3D898AF7",
    x"3D8979C7",
    x"3D896899",
    x"3D89576D",
    x"3D894643",
    x"3D89351B",
    x"3D8923F6",
    x"3D8912D2",
    x"3D8901B1",
    x"3D88F092",
    x"3D88DF75",
    x"3D88CE5A",
    x"3D88BD41",
    x"3D88AC2B",
    x"3D889B16",
    x"3D888A04",
    x"3D8878F4",
    x"3D8867E6",
    x"3D8856DA",
    x"3D8845D0",
    x"3D8834C8",
    x"3D8823C3",
    x"3D8812BF",
    x"3D8801BE",
    x"3D87F0BF",
    x"3D87DFC2",
    x"3D87CEC7",
    x"3D87BDCE",
    x"3D87ACD7",
    x"3D879BE3",
    x"3D878AF0",
    x"3D877A00",
    x"3D876912",
    x"3D875826",
    x"3D87473C",
    x"3D873654",
    x"3D87256E",
    x"3D87148B",
    x"3D8703A9",
    x"3D86F2CA",
    x"3D86E1ED",
    x"3D86D111",
    x"3D86C038",
    x"3D86AF61",
    x"3D869E8C",
    x"3D868DBA",
    x"3D867CE9",
    x"3D866C1A",
    x"3D865B4E",
    x"3D864A84",
    x"3D8639BB",
    x"3D8628F5",
    x"3D861831",
    x"3D86076F",
    x"3D85F6AF",
    x"3D85E5F1",
    x"3D85D536",
    x"3D85C47C",
    x"3D85B3C5",
    x"3D85A30F",
    x"3D85925C",
    x"3D8581AB",
    x"3D8570FB",
    x"3D85604E",
    x"3D854FA3",
    x"3D853EFA",
    x"3D852E54",
    x"3D851DAF",
    x"3D850D0C",
    x"3D84FC6C",
    x"3D84EBCD",
    x"3D84DB31",
    x"3D84CA96",
    x"3D84B9FE",
    x"3D84A968",
    x"3D8498D4",
    x"3D848842",
    x"3D8477B2",
    x"3D846724",
    x"3D845698",
    x"3D84460E",
    x"3D843586",
    x"3D842501",
    x"3D84147D",
    x"3D8403FC",
    x"3D83F37C",
    x"3D83E2FF",
    x"3D83D283",
    x"3D83C20A",
    x"3D83B193",
    x"3D83A11E",
    x"3D8390AB",
    x"3D838039",
    x"3D836FCA",
    x"3D835F5D",
    x"3D834EF3",
    x"3D833E8A",
    x"3D832E23",
    x"3D831DBE",
    x"3D830D5C",
    x"3D82FCFB",
    x"3D82EC9C",
    x"3D82DC40",
    x"3D82CBE5",
    x"3D82BB8D",
    x"3D82AB36",
    x"3D829AE2",
    x"3D828A90",
    x"3D827A3F",
    x"3D8269F1",
    x"3D8259A5",
    x"3D82495B",
    x"3D823912",
    x"3D8228CC",
    x"3D821888",
    x"3D820846",
    x"3D81F806",
    x"3D81E7C8",
    x"3D81D78C",
    x"3D81C752",
    x"3D81B71A",
    x"3D81A6E5",
    x"3D8196B1",
    x"3D81867F",
    x"3D81764F",
    x"3D816621",
    x"3D8155F6",
    x"3D8145CC",
    x"3D8135A4",
    x"3D81257E",
    x"3D81155B",
    x"3D810539",
    x"3D80F519",
    x"3D80E4FC",
    x"3D80D4E0",
    x"3D80C4C7",
    x"3D80B4AF",
    x"3D80A499",
    x"3D809486",
    x"3D808474",
    x"3D807465",
    x"3D806457",
    x"3D80544C",
    x"3D804442",
    x"3D80343B",
    x"3D802435",
    x"3D801432",
    x"3D800430",
    x"3D7FE861",
    x"3D7FC866",
    x"3D7FA86F",
    x"3D7F887C",
    x"3D7F688D",
    x"3D7F48A2",
    x"3D7F28BB",
    x"3D7F08D7",
    x"3D7EE8F8",
    x"3D7EC91D",
    x"3D7EA946",
    x"3D7E8973",
    x"3D7E69A4",
    x"3D7E49D9",
    x"3D7E2A11",
    x"3D7E0A4E",
    x"3D7DEA8F",
    x"3D7DCAD3",
    x"3D7DAB1C",
    x"3D7D8B69",
    x"3D7D6BB9",
    x"3D7D4C0E",
    x"3D7D2C66",
    x"3D7D0CC3",
    x"3D7CED23",
    x"3D7CCD87",
    x"3D7CADF0",
    x"3D7C8E5C",
    x"3D7C6ECC",
    x"3D7C4F40",
    x"3D7C2FB8",
    x"3D7C1034",
    x"3D7BF0B4",
    x"3D7BD138",
    x"3D7BB1C0",
    x"3D7B924C",
    x"3D7B72DB",
    x"3D7B536F",
    x"3D7B3406",
    x"3D7B14A2",
    x"3D7AF541",
    x"3D7AD5E4",
    x"3D7AB68C",
    x"3D7A9737",
    x"3D7A77E6",
    x"3D7A5899",
    x"3D7A3950",
    x"3D7A1A0B",
    x"3D79FAC9",
    x"3D79DB8C",
    x"3D79BC52",
    x"3D799D1D",
    x"3D797DEB",
    x"3D795EBD",
    x"3D793F93",
    x"3D79206D",
    x"3D79014B",
    x"3D78E22D",
    x"3D78C313",
    x"3D78A3FC",
    x"3D7884EA",
    x"3D7865DB",
    x"3D7846D0",
    x"3D7827C9",
    x"3D7808C6",
    x"3D77E9C7",
    x"3D77CACC",
    x"3D77ABD4",
    x"3D778CE1",
    x"3D776DF1",
    x"3D774F05",
    x"3D77301E",
    x"3D771139",
    x"3D76F259",
    x"3D76D37D",
    x"3D76B4A4",
    x"3D7695D0",
    x"3D7676FF",
    x"3D765832",
    x"3D763969",
    x"3D761AA4",
    x"3D75FBE2",
    x"3D75DD25",
    x"3D75BE6B",
    x"3D759FB5",
    x"3D758103",
    x"3D756255",
    x"3D7543AA",
    x"3D752504",
    x"3D750661",
    x"3D74E7C2",
    x"3D74C927",
    x"3D74AA90",
    x"3D748BFD",
    x"3D746D6D",
    x"3D744EE1",
    x"3D743059",
    x"3D7411D5",
    x"3D73F355",
    x"3D73D4D8",
    x"3D73B660",
    x"3D7397EB",
    x"3D73797A",
    x"3D735B0C",
    x"3D733CA3",
    x"3D731E3D",
    x"3D72FFDB",
    x"3D72E17D",
    x"3D72C323",
    x"3D72A4CC",
    x"3D72867A",
    x"3D72682B",
    x"3D7249E0",
    x"3D722B98",
    x"3D720D55",
    x"3D71EF15",
    x"3D71D0D9",
    x"3D71B2A1",
    x"3D71946C",
    x"3D71763C",
    x"3D71580F",
    x"3D7139E6",
    x"3D711BC0",
    x"3D70FD9F",
    x"3D70DF81",
    x"3D70C167",
    x"3D70A351",
    x"3D70853E",
    x"3D70672F",
    x"3D704924",
    x"3D702B1D",
    x"3D700D19",
    x"3D6FEF1A",
    x"3D6FD11E",
    x"3D6FB325",
    x"3D6F9531",
    x"3D6F7740",
    x"3D6F5953",
    x"3D6F3B6A",
    x"3D6F1D84",
    x"3D6EFFA2",
    x"3D6EE1C4",
    x"3D6EC3EA",
    x"3D6EA613",
    x"3D6E8840",
    x"3D6E6A71",
    x"3D6E4CA6",
    x"3D6E2EDE",
    x"3D6E111A",
    x"3D6DF35A",
    x"3D6DD59D",
    x"3D6DB7E4",
    x"3D6D9A2F",
    x"3D6D7C7E",
    x"3D6D5ED0",
    x"3D6D4126",
    x"3D6D2380",
    x"3D6D05DD",
    x"3D6CE83E",
    x"3D6CCAA3",
    x"3D6CAD0C",
    x"3D6C8F78",
    x"3D6C71E8",
    x"3D6C545B",
    x"3D6C36D3",
    x"3D6C194E",
    x"3D6BFBCC",
    x"3D6BDE4F",
    x"3D6BC0D5",
    x"3D6BA35F",
    x"3D6B85EC",
    x"3D6B687D",
    x"3D6B4B12",
    x"3D6B2DAA",
    x"3D6B1046",
    x"3D6AF2E6",
    x"3D6AD58A",
    x"3D6AB831",
    x"3D6A9ADC",
    x"3D6A7D8A",
    x"3D6A603C",
    x"3D6A42F2",
    x"3D6A25AC",
    x"3D6A0869",
    x"3D69EB29",
    x"3D69CDEE",
    x"3D69B0B6",
    x"3D699382",
    x"3D697651",
    x"3D695924",
    x"3D693BFB",
    x"3D691ED5",
    x"3D6901B3",
    x"3D68E495",
    x"3D68C77A",
    x"3D68AA63",
    x"3D688D4F",
    x"3D687040",
    x"3D685333",
    x"3D68362B",
    x"3D681926",
    x"3D67FC24",
    x"3D67DF27",
    x"3D67C22D",
    x"3D67A536",
    x"3D678843",
    x"3D676B54",
    x"3D674E69",
    x"3D673181",
    x"3D67149C",
    x"3D66F7BB",
    x"3D66DADE",
    x"3D66BE05",
    x"3D66A12F",
    x"3D66845C",
    x"3D66678E",
    x"3D664AC2",
    x"3D662DFB",
    x"3D661137",
    x"3D65F477",
    x"3D65D7BA",
    x"3D65BB01",
    x"3D659E4B",
    x"3D658199",
    x"3D6564EB",
    x"3D654840",
    x"3D652B99",
    x"3D650EF5",
    x"3D64F255",
    x"3D64D5B8",
    x"3D64B91F",
    x"3D649C8A",
    x"3D647FF8",
    x"3D64636A",
    x"3D6446DF",
    x"3D642A58",
    x"3D640DD5",
    x"3D63F155",
    x"3D63D4D9",
    x"3D63B860",
    x"3D639BEA",
    x"3D637F79",
    x"3D63630B",
    x"3D6346A0",
    x"3D632A39",
    x"3D630DD5",
    x"3D62F175",
    x"3D62D519",
    x"3D62B8C0",
    x"3D629C6B",
    x"3D628019",
    x"3D6263CB",
    x"3D624780",
    x"3D622B39",
    x"3D620EF5",
    x"3D61F2B5",
    x"3D61D679",
    x"3D61BA40",
    x"3D619E0A",
    x"3D6181D8",
    x"3D6165AA",
    x"3D61497F",
    x"3D612D57",
    x"3D611133",
    x"3D60F513",
    x"3D60D8F6",
    x"3D60BCDD",
    x"3D60A0C7",
    x"3D6084B5",
    x"3D6068A6",
    x"3D604C9A",
    x"3D603093",
    x"3D60148E",
    x"3D5FF88D",
    x"3D5FDC90",
    x"3D5FC096",
    x"3D5FA4A0",
    x"3D5F88AD",
    x"3D5F6CBE",
    x"3D5F50D2",
    x"3D5F34EA",
    x"3D5F1905",
    x"3D5EFD23",
    x"3D5EE145",
    x"3D5EC56B",
    x"3D5EA994",
    x"3D5E8DC1",
    x"3D5E71F1",
    x"3D5E5624",
    x"3D5E3A5B",
    x"3D5E1E96",
    x"3D5E02D3",
    x"3D5DE715",
    x"3D5DCB5A",
    x"3D5DAFA2",
    x"3D5D93EE",
    x"3D5D783D",
    x"3D5D5C90",
    x"3D5D40E6",
    x"3D5D253F",
    x"3D5D099D",
    x"3D5CEDFD",
    x"3D5CD261",
    x"3D5CB6C8",
    x"3D5C9B33",
    x"3D5C7FA2",
    x"3D5C6413",
    x"3D5C4889",
    x"3D5C2D01",
    x"3D5C117D",
    x"3D5BF5FD",
    x"3D5BDA80",
    x"3D5BBF06",
    x"3D5BA390",
    x"3D5B881D",
    x"3D5B6CAE",
    x"3D5B5142",
    x"3D5B35DA",
    x"3D5B1A75",
    x"3D5AFF13",
    x"3D5AE3B5",
    x"3D5AC85A",
    x"3D5AAD03",
    x"3D5A91AF",
    x"3D5A765E",
    x"3D5A5B11",
    x"3D5A3FC8",
    x"3D5A2481",
    x"3D5A093F",
    x"3D59EDFF",
    x"3D59D2C3",
    x"3D59B78A",
    x"3D599C55",
    x"3D598123",
    x"3D5965F5",
    x"3D594ACA",
    x"3D592FA2",
    x"3D59147E",
    x"3D58F95D",
    x"3D58DE40",
    x"3D58C326",
    x"3D58A80F",
    x"3D588CFC",
    x"3D5871EC",
    x"3D5856DF",
    x"3D583BD6",
    x"3D5820D0",
    x"3D5805CE",
    x"3D57EACF",
    x"3D57CFD3",
    x"3D57B4DB",
    x"3D5799E6",
    x"3D577EF4",
    x"3D576406",
    x"3D57491B",
    x"3D572E34",
    x"3D571350",
    x"3D56F86F",
    x"3D56DD92",
    x"3D56C2B8",
    x"3D56A7E1",
    x"3D568D0E",
    x"3D56723E",
    x"3D565771",
    x"3D563CA8",
    x"3D5621E2",
    x"3D56071F",
    x"3D55EC60",
    x"3D55D1A4",
    x"3D55B6EC",
    x"3D559C36",
    x"3D558185",
    x"3D5566D6",
    x"3D554C2B",
    x"3D553183",
    x"3D5516DE",
    x"3D54FC3D",
    x"3D54E19F",
    x"3D54C705",
    x"3D54AC6E",
    x"3D5491DA",
    x"3D547749",
    x"3D545CBC",
    x"3D544232",
    x"3D5427AB",
    x"3D540D28",
    x"3D53F2A8",
    x"3D53D82B",
    x"3D53BDB2",
    x"3D53A33C",
    x"3D5388C9",
    x"3D536E5A",
    x"3D5353EE",
    x"3D533985",
    x"3D531F1F",
    x"3D5304BD",
    x"3D52EA5E",
    x"3D52D002",
    x"3D52B5AA",
    x"3D529B55",
    x"3D528103",
    x"3D5266B5",
    x"3D524C6A",
    x"3D523222",
    x"3D5217DD",
    x"3D51FD9C",
    x"3D51E35E",
    x"3D51C923",
    x"3D51AEEB",
    x"3D5194B7",
    x"3D517A86",
    x"3D516059",
    x"3D51462E",
    x"3D512C07",
    x"3D5111E3",
    x"3D50F7C3",
    x"3D50DDA5",
    x"3D50C38B",
    x"3D50A974",
    x"3D508F61",
    x"3D507550",
    x"3D505B43",
    x"3D50413A",
    x"3D502733",
    x"3D500D30",
    x"3D4FF330",
    x"3D4FD933",
    x"3D4FBF39",
    x"3D4FA543",
    x"3D4F8B50",
    x"3D4F7160",
    x"3D4F5774",
    x"3D4F3D8B",
    x"3D4F23A4",
    x"3D4F09C2",
    x"3D4EEFE2",
    x"3D4ED606",
    x"3D4EBC2D",
    x"3D4EA257",
    x"3D4E8884",
    x"3D4E6EB4",
    x"3D4E54E8",
    x"3D4E3B1F",
    x"3D4E2159",
    x"3D4E0797",
    x"3D4DEDD8",
    x"3D4DD41B",
    x"3D4DBA63",
    x"3D4DA0AD",
    x"3D4D86FA",
    x"3D4D6D4B",
    x"3D4D539F",
    x"3D4D39F6",
    x"3D4D2051",
    x"3D4D06AE",
    x"3D4CED0F",
    x"3D4CD373",
    x"3D4CB9DA",
    x"3D4CA044",
    x"3D4C86B2",
    x"3D4C6D23",
    x"3D4C5397",
    x"3D4C3A0E",
    x"3D4C2088",
    x"3D4C0706",
    x"3D4BED86",
    x"3D4BD40A",
    x"3D4BBA91",
    x"3D4BA11C",
    x"3D4B87A9",
    x"3D4B6E3A",
    x"3D4B54CE",
    x"3D4B3B65",
    x"3D4B21FF",
    x"3D4B089C",
    x"3D4AEF3D",
    x"3D4AD5E0",
    x"3D4ABC87",
    x"3D4AA331",
    x"3D4A89DE",
    x"3D4A708F",
    x"3D4A5742",
    x"3D4A3DF9",
    x"3D4A24B3",
    x"3D4A0B70",
    x"3D49F230",
    x"3D49D8F3",
    x"3D49BFBA",
    x"3D49A683",
    x"3D498D50",
    x"3D497420",
    x"3D495AF3",
    x"3D4941C9",
    x"3D4928A2",
    x"3D490F7F",
    x"3D48F65F",
    x"3D48DD41",
    x"3D48C427",
    x"3D48AB10",
    x"3D4891FC",
    x"3D4878EC",
    x"3D485FDE",
    x"3D4846D4",
    x"3D482DCD",
    x"3D4814C8",
    x"3D47FBC7",
    x"3D47E2C9",
    x"3D47C9CF",
    x"3D47B0D7",
    x"3D4797E2",
    x"3D477EF1",
    x"3D476603",
    x"3D474D18",
    x"3D47342F",
    x"3D471B4A",
    x"3D470269",
    x"3D46E98A",
    x"3D46D0AE",
    x"3D46B7D6",
    x"3D469F00",
    x"3D46862E",
    x"3D466D5F",
    x"3D465493",
    x"3D463BCA",
    x"3D462304",
    x"3D460A41",
    x"3D45F181",
    x"3D45D8C4",
    x"3D45C00B",
    x"3D45A754",
    x"3D458EA1",
    x"3D4575F1",
    x"3D455D44",
    x"3D454499",
    x"3D452BF2",
    x"3D45134E",
    x"3D44FAAE",
    x"3D44E210",
    x"3D44C975",
    x"3D44B0DD",
    x"3D449849",
    x"3D447FB7",
    x"3D446729",
    x"3D444E9E",
    x"3D443615",
    x"3D441D90",
    x"3D44050E",
    x"3D43EC8F",
    x"3D43D413",
    x"3D43BB9A",
    x"3D43A324",
    x"3D438AB1",
    x"3D437241",
    x"3D4359D4",
    x"3D43416B",
    x"3D432904",
    x"3D4310A0",
    x"3D42F840",
    x"3D42DFE2",
    x"3D42C788",
    x"3D42AF31",
    x"3D4296DC",
    x"3D427E8B",
    x"3D42663D",
    x"3D424DF1",
    x"3D4235A9",
    x"3D421D64",
    x"3D420522",
    x"3D41ECE3",
    x"3D41D4A6",
    x"3D41BC6D",
    x"3D41A437",
    x"3D418C04",
    x"3D4173D4",
    x"3D415BA7",
    x"3D41437D",
    x"3D412B57",
    x"3D411333",
    x"3D40FB12",
    x"3D40E2F4",
    x"3D40CAD9",
    x"3D40B2C1",
    x"3D409AAC",
    x"3D40829A",
    x"3D406A8C",
    x"3D405280",
    x"3D403A77",
    x"3D402271",
    x"3D400A6E",
    x"3D3FF26F",
    x"3D3FDA72",
    x"3D3FC278",
    x"3D3FAA81",
    x"3D3F928D",
    x"3D3F7A9D",
    x"3D3F62AF",
    x"3D3F4AC4",
    x"3D3F32DC",
    x"3D3F1AF7",
    x"3D3F0315",
    x"3D3EEB36",
    x"3D3ED35A",
    x"3D3EBB82",
    x"3D3EA3AC",
    x"3D3E8BD9",
    x"3D3E7409",
    x"3D3E5C3C",
    x"3D3E4472",
    x"3D3E2CAA",
    x"3D3E14E6",
    x"3D3DFD25",
    x"3D3DE567",
    x"3D3DCDAC",
    x"3D3DB5F4",
    x"3D3D9E3E",
    x"3D3D868C",
    x"3D3D6EDD",
    x"3D3D5730",
    x"3D3D3F87",
    x"3D3D27E1",
    x"3D3D103D",
    x"3D3CF89C",
    x"3D3CE0FF",
    x"3D3CC964",
    x"3D3CB1CD",
    x"3D3C9A38",
    x"3D3C82A6",
    x"3D3C6B17",
    x"3D3C538B",
    x"3D3C3C02",
    x"3D3C247C",
    x"3D3C0CF9",
    x"3D3BF579",
    x"3D3BDDFC",
    x"3D3BC681",
    x"3D3BAF0A",
    x"3D3B9796",
    x"3D3B8024",
    x"3D3B68B6",
    x"3D3B514A",
    x"3D3B39E1",
    x"3D3B227C",
    x"3D3B0B19",
    x"3D3AF3B9",
    x"3D3ADC5C",
    x"3D3AC502",
    x"3D3AADAB",
    x"3D3A9656",
    x"3D3A7F05",
    x"3D3A67B7",
    x"3D3A506B",
    x"3D3A3922",
    x"3D3A21DD",
    x"3D3A0A9A",
    x"3D39F35A",
    x"3D39DC1D",
    x"3D39C4E3",
    x"3D39ADAC",
    x"3D399678",
    x"3D397F46",
    x"3D396818",
    x"3D3950EC",
    x"3D3939C4",
    x"3D39229E",
    x"3D390B7B",
    x"3D38F45B",
    x"3D38DD3E",
    x"3D38C624",
    x"3D38AF0C",
    x"3D3897F8",
    x"3D3880E6",
    x"3D3869D8",
    x"3D3852CC",
    x"3D383BC3",
    x"3D3824BD",
    x"3D380DBA",
    x"3D37F6B9",
    x"3D37DFBC",
    x"3D37C8C2",
    x"3D37B1CA",
    x"3D379AD5",
    x"3D3783E3",
    x"3D376CF4",
    x"3D375608",
    x"3D373F1F",
    x"3D372838",
    x"3D371155",
    x"3D36FA74",
    x"3D36E396",
    x"3D36CCBB",
    x"3D36B5E3",
    x"3D369F0D",
    x"3D36883B",
    x"3D36716B",
    x"3D365A9F",
    x"3D3643D5",
    x"3D362D0E",
    x"3D361649",
    x"3D35FF88",
    x"3D35E8CA",
    x"3D35D20E",
    x"3D35BB55",
    x"3D35A49F",
    x"3D358DEC",
    x"3D35773C",
    x"3D35608E",
    x"3D3549E3",
    x"3D35333C",
    x"3D351C97",
    x"3D3505F4",
    x"3D34EF55",
    x"3D34D8B9",
    x"3D34C21F",
    x"3D34AB88",
    x"3D3494F4",
    x"3D347E63",
    x"3D3467D4",
    x"3D345149",
    x"3D343AC0",
    x"3D34243A",
    x"3D340DB7",
    x"3D33F737",
    x"3D33E0B9",
    x"3D33CA3F",
    x"3D33B3C7",
    x"3D339D52",
    x"3D3386DF",
    x"3D337070",
    x"3D335A03",
    x"3D334399",
    x"3D332D32",
    x"3D3316CE",
    x"3D33006D",
    x"3D32EA0E",
    x"3D32D3B2",
    x"3D32BD59",
    x"3D32A703",
    x"3D3290AF",
    x"3D327A5F",
    x"3D326411",
    x"3D324DC6",
    x"3D32377D",
    x"3D322138",
    x"3D320AF5",
    x"3D31F4B5",
    x"3D31DE78",
    x"3D31C83D",
    x"3D31B206",
    x"3D319BD1",
    x"3D31859F",
    x"3D316F70",
    x"3D315943",
    x"3D314319",
    x"3D312CF2",
    x"3D3116CE",
    x"3D3100AD",
    x"3D30EA8E",
    x"3D30D472",
    x"3D30BE59",
    x"3D30A842",
    x"3D30922F",
    x"3D307C1E",
    x"3D306610",
    x"3D305004",
    x"3D3039FC",
    x"3D3023F6",
    x"3D300DF3",
    x"3D2FF7F2",
    x"3D2FE1F5",
    x"3D2FCBFA",
    x"3D2FB602",
    x"3D2FA00C",
    x"3D2F8A1A",
    x"3D2F742A",
    x"3D2F5E3D",
    x"3D2F4852",
    x"3D2F326A",
    x"3D2F1C86",
    x"3D2F06A3",
    x"3D2EF0C4",
    x"3D2EDAE7",
    x"3D2EC50D",
    x"3D2EAF36",
    x"3D2E9961",
    x"3D2E8390",
    x"3D2E6DC0",
    x"3D2E57F4",
    x"3D2E422A",
    x"3D2E2C64",
    x"3D2E169F",
    x"3D2E00DE",
    x"3D2DEB1F",
    x"3D2DD563",
    x"3D2DBFAA",
    x"3D2DA9F3",
    x"3D2D943F",
    x"3D2D7E8E",
    x"3D2D68E0",
    x"3D2D5334",
    x"3D2D3D8B",
    x"3D2D27E5",
    x"3D2D1241",
    x"3D2CFCA0",
    x"3D2CE702",
    x"3D2CD166",
    x"3D2CBBCD",
    x"3D2CA637",
    x"3D2C90A4",
    x"3D2C7B13",
    x"3D2C6585",
    x"3D2C4FFA",
    x"3D2C3A71",
    x"3D2C24EB",
    x"3D2C0F68",
    x"3D2BF9E7",
    x"3D2BE469",
    x"3D2BCEEE",
    x"3D2BB976",
    x"3D2BA400",
    x"3D2B8E8D",
    x"3D2B791C",
    x"3D2B63AE",
    x"3D2B4E43",
    x"3D2B38DB",
    x"3D2B2375",
    x"3D2B0E12",
    x"3D2AF8B2",
    x"3D2AE354",
    x"3D2ACDF9",
    x"3D2AB8A0",
    x"3D2AA34B",
    x"3D2A8DF7",
    x"3D2A78A7",
    x"3D2A6359",
    x"3D2A4E0E",
    x"3D2A38C6",
    x"3D2A2380",
    x"3D2A0E3D",
    x"3D29F8FC",
    x"3D29E3BF",
    x"3D29CE84",
    x"3D29B94B",
    x"3D29A415",
    x"3D298EE2",
    x"3D2979B1",
    x"3D296484",
    x"3D294F58",
    x"3D293A30",
    x"3D29250A",
    x"3D290FE6",
    x"3D28FAC6",
    x"3D28E5A8",
    x"3D28D08C",
    x"3D28BB74",
    x"3D28A65E",
    x"3D28914A",
    x"3D287C39",
    x"3D28672B",
    x"3D28521F",
    x"3D283D16",
    x"3D282810",
    x"3D28130C",
    x"3D27FE0B",
    x"3D27E90D",
    x"3D27D411",
    x"3D27BF18",
    x"3D27AA21",
    x"3D27952D",
    x"3D27803C",
    x"3D276B4D",
    x"3D275661",
    x"3D274178",
    x"3D272C91",
    x"3D2717AD",
    x"3D2702CB",
    x"3D26EDEC",
    x"3D26D90F",
    x"3D26C436",
    x"3D26AF5E",
    x"3D269A8A",
    x"3D2685B8",
    x"3D2670E8",
    x"3D265C1C",
    x"3D264751",
    x"3D26328A",
    x"3D261DC5",
    x"3D260902",
    x"3D25F442",
    x"3D25DF85",
    x"3D25CACB",
    x"3D25B613",
    x"3D25A15D",
    x"3D258CAA",
    x"3D2577FA",
    x"3D25634C",
    x"3D254EA1",
    x"3D2539F9",
    x"3D252553",
    x"3D2510AF",
    x"3D24FC0E",
    x"3D24E770",
    x"3D24D2D5",
    x"3D24BE3B",
    x"3D24A9A5",
    x"3D249511",
    x"3D248080",
    x"3D246BF1",
    x"3D245765",
    x"3D2442DB",
    x"3D242E54",
    x"3D2419D0",
    x"3D24054E",
    x"3D23F0CE",
    x"3D23DC51",
    x"3D23C7D7",
    x"3D23B35F",
    x"3D239EEA",
    x"3D238A78",
    x"3D237608",
    x"3D23619A",
    x"3D234D2F",
    x"3D2338C7",
    x"3D232461",
    x"3D230FFE",
    x"3D22FB9D",
    x"3D22E73F",
    x"3D22D2E3",
    x"3D22BE8A",
    x"3D22AA34",
    x"3D2295E0",
    x"3D22818E",
    x"3D226D3F",
    x"3D2258F3",
    x"3D2244A9",
    x"3D223062",
    x"3D221C1D",
    x"3D2207DB",
    x"3D21F39B",
    x"3D21DF5E",
    x"3D21CB23",
    x"3D21B6EB",
    x"3D21A2B5",
    x"3D218E82",
    x"3D217A52",
    x"3D216624",
    x"3D2151F8",
    x"3D213DCF",
    x"3D2129A9",
    x"3D211585",
    x"3D210163",
    x"3D20ED44",
    x"3D20D928",
    x"3D20C50E",
    x"3D20B0F7",
    x"3D209CE2",
    x"3D2088D0",
    x"3D2074C0",
    x"3D2060B2",
    x"3D204CA8",
    x"3D20389F",
    x"3D202499",
    x"3D201096",
    x"3D1FFC95",
    x"3D1FE897",
    x"3D1FD49B",
    x"3D1FC0A2",
    x"3D1FACAB",
    x"3D1F98B7",
    x"3D1F84C5",
    x"3D1F70D5",
    x"3D1F5CE9",
    x"3D1F48FE",
    x"3D1F3516",
    x"3D1F2131",
    x"3D1F0D4E",
    x"3D1EF96E",
    x"3D1EE590",
    x"3D1ED1B4",
    x"3D1EBDDB",
    x"3D1EAA05",
    x"3D1E9631",
    x"3D1E825F",
    x"3D1E6E90",
    x"3D1E5AC4",
    x"3D1E46F9",
    x"3D1E3332",
    x"3D1E1F6D",
    x"3D1E0BAA",
    x"3D1DF7EA",
    x"3D1DE42C",
    x"3D1DD071",
    x"3D1DBCB8",
    x"3D1DA901",
    x"3D1D954E",
    x"3D1D819C",
    x"3D1D6DED",
    x"3D1D5A41",
    x"3D1D4697",
    x"3D1D32EF",
    x"3D1D1F4A",
    x"3D1D0BA7",
    x"3D1CF807",
    x"3D1CE469",
    x"3D1CD0CE",
    x"3D1CBD35",
    x"3D1CA99F",
    x"3D1C960B",
    x"3D1C8279",
    x"3D1C6EEA",
    x"3D1C5B5D",
    x"3D1C47D3",
    x"3D1C344B",
    x"3D1C20C6",
    x"3D1C0D43",
    x"3D1BF9C3",
    x"3D1BE645",
    x"3D1BD2C9",
    x"3D1BBF50",
    x"3D1BABD9",
    x"3D1B9865",
    x"3D1B84F3",
    x"3D1B7184",
    x"3D1B5E17",
    x"3D1B4AAC",
    x"3D1B3744",
    x"3D1B23DE",
    x"3D1B107B",
    x"3D1AFD1A",
    x"3D1AE9BC",
    x"3D1AD660",
    x"3D1AC306",
    x"3D1AAFAF",
    x"3D1A9C5A",
    x"3D1A8908",
    x"3D1A75B8",
    x"3D1A626B",
    x"3D1A4F20",
    x"3D1A3BD7",
    x"3D1A2891",
    x"3D1A154D",
    x"3D1A020B",
    x"3D19EECC",
    x"3D19DB90",
    x"3D19C855",
    x"3D19B51D",
    x"3D19A1E8",
    x"3D198EB5",
    x"3D197B84",
    x"3D196856",
    x"3D19552A",
    x"3D194201",
    x"3D192EDA",
    x"3D191BB5",
    x"3D190893",
    x"3D18F573",
    x"3D18E255",
    x"3D18CF3A",
    x"3D18BC22",
    x"3D18A90B",
    x"3D1895F7",
    x"3D1882E6",
    x"3D186FD7",
    x"3D185CCA",
    x"3D1849C0",
    x"3D1836B7",
    x"3D1823B2",
    x"3D1810AF",
    x"3D17FDAE",
    x"3D17EAAF",
    x"3D17D7B3",
    x"3D17C4B9",
    x"3D17B1C2",
    x"3D179ECD",
    x"3D178BDA",
    x"3D1778EA",
    x"3D1765FC",
    x"3D175310",
    x"3D174027",
    x"3D172D40",
    x"3D171A5C",
    x"3D17077A",
    x"3D16F49A",
    x"3D16E1BD",
    x"3D16CEE1",
    x"3D16BC09",
    x"3D16A932",
    x"3D16965F",
    x"3D16838D",
    x"3D1670BE",
    x"3D165DF1",
    x"3D164B26",
    x"3D16385E",
    x"3D162598",
    x"3D1612D5",
    x"3D160013",
    x"3D15ED54",
    x"3D15DA98",
    x"3D15C7DE",
    x"3D15B526",
    x"3D15A271",
    x"3D158FBD",
    x"3D157D0D",
    x"3D156A5E",
    x"3D1557B2",
    x"3D154508",
    x"3D153261",
    x"3D151FBC",
    x"3D150D19",
    x"3D14FA78",
    x"3D14E7DA",
    x"3D14D53E",
    x"3D14C2A5",
    x"3D14B00E",
    x"3D149D79",
    x"3D148AE6",
    x"3D147856",
    x"3D1465C8",
    x"3D14533D",
    x"3D1440B3",
    x"3D142E2D",
    x"3D141BA8",
    x"3D140926",
    x"3D13F6A6",
    x"3D13E428",
    x"3D13D1AD",
    x"3D13BF34",
    x"3D13ACBD",
    x"3D139A48",
    x"3D1387D6",
    x"3D137566",
    x"3D1362F9",
    x"3D13508E",
    x"3D133E25",
    x"3D132BBE",
    x"3D13195A",
    x"3D1306F8",
    x"3D12F498",
    x"3D12E23B",
    x"3D12CFE0",
    x"3D12BD87",
    x"3D12AB30",
    x"3D1298DC",
    x"3D12868A",
    x"3D12743A",
    x"3D1261ED",
    x"3D124FA2",
    x"3D123D59",
    x"3D122B12",
    x"3D1218CE",
    x"3D12068C",
    x"3D11F44D",
    x"3D11E20F",
    x"3D11CFD4",
    x"3D11BD9B",
    x"3D11AB65",
    x"3D119930",
    x"3D1186FE",
    x"3D1174CF",
    x"3D1162A1",
    x"3D115076",
    x"3D113E4D",
    x"3D112C26",
    x"3D111A02",
    x"3D1107E0",
    x"3D10F5C0",
    x"3D10E3A2",
    x"3D10D187",
    x"3D10BF6E",
    x"3D10AD57",
    x"3D109B43",
    x"3D108930",
    x"3D107720",
    x"3D106513",
    x"3D105307",
    x"3D1040FE",
    x"3D102EF7",
    x"3D101CF2",
    x"3D100AF0",
    x"3D0FF8EF",
    x"3D0FE6F1",
    x"3D0FD4F6",
    x"3D0FC2FC",
    x"3D0FB105",
    x"3D0F9F10",
    x"3D0F8D1D",
    x"3D0F7B2D",
    x"3D0F693E",
    x"3D0F5752",
    x"3D0F4569",
    x"3D0F3381",
    x"3D0F219C",
    x"3D0F0FB9",
    x"3D0EFDD8",
    x"3D0EEBF9",
    x"3D0EDA1D",
    x"3D0EC843",
    x"3D0EB66B",
    x"3D0EA495",
    x"3D0E92C2",
    x"3D0E80F0",
    x"3D0E6F21",
    x"3D0E5D55",
    x"3D0E4B8A",
    x"3D0E39C2",
    x"3D0E27FC",
    x"3D0E1638",
    x"3D0E0476",
    x"3D0DF2B7",
    x"3D0DE0F9",
    x"3D0DCF3E",
    x"3D0DBD85",
    x"3D0DABCF",
    x"3D0D9A1B",
    x"3D0D8868",
    x"3D0D76B8",
    x"3D0D650B",
    x"3D0D535F",
    x"3D0D41B6",
    x"3D0D300F",
    x"3D0D1E6A",
    x"3D0D0CC7",
    x"3D0CFB27",
    x"3D0CE988",
    x"3D0CD7EC",
    x"3D0CC652",
    x"3D0CB4BB",
    x"3D0CA325",
    x"3D0C9192",
    x"3D0C8001",
    x"3D0C6E72",
    x"3D0C5CE5",
    x"3D0C4B5B",
    x"3D0C39D2",
    x"3D0C284C",
    x"3D0C16C8",
    x"3D0C0546",
    x"3D0BF3C7",
    x"3D0BE24A",
    x"3D0BD0CE",
    x"3D0BBF55",
    x"3D0BADDF",
    x"3D0B9C6A",
    x"3D0B8AF7",
    x"3D0B7987",
    x"3D0B6819",
    x"3D0B56AD",
    x"3D0B4543",
    x"3D0B33DC",
    x"3D0B2276",
    x"3D0B1113",
    x"3D0AFFB2",
    x"3D0AEE53",
    x"3D0ADCF7",
    x"3D0ACB9C",
    x"3D0ABA44",
    x"3D0AA8ED",
    x"3D0A9799",
    x"3D0A8648",
    x"3D0A74F8",
    x"3D0A63AA",
    x"3D0A525F",
    x"3D0A4116",
    x"3D0A2FCF",
    x"3D0A1E8A",
    x"3D0A0D47",
    x"3D09FC06",
    x"3D09EAC8",
    x"3D09D98C",
    x"3D09C852",
    x"3D09B71A",
    x"3D09A5E4",
    x"3D0994B0",
    x"3D09837F",
    x"3D09724F",
    x"3D096122",
    x"3D094FF7",
    x"3D093ECE",
    x"3D092DA7",
    x"3D091C83",
    x"3D090B60",
    x"3D08FA40",
    x"3D08E922",
    x"3D08D806",
    x"3D08C6EC",
    x"3D08B5D4",
    x"3D08A4BE",
    x"3D0893AB",
    x"3D088299",
    x"3D08718A",
    x"3D08607D",
    x"3D084F72",
    x"3D083E69",
    x"3D082D62",
    x"3D081C5E",
    x"3D080B5B",
    x"3D07FA5B",
    x"3D07E95D",
    x"3D07D860",
    x"3D07C767",
    x"3D07B66F",
    x"3D07A579",
    x"3D079485",
    x"3D078394",
    x"3D0772A4",
    x"3D0761B7",
    x"3D0750CC",
    x"3D073FE3",
    x"3D072EFC",
    x"3D071E17",
    x"3D070D34",
    x"3D06FC54",
    x"3D06EB75",
    x"3D06DA99",
    x"3D06C9BF",
    x"3D06B8E7",
    x"3D06A810",
    x"3D06973D",
    x"3D06866B",
    x"3D06759B",
    x"3D0664CD",
    x"3D065402",
    x"3D064338",
    x"3D063271",
    x"3D0621AC",
    x"3D0610E9",
    x"3D060027",
    x"3D05EF68",
    x"3D05DEAC",
    x"3D05CDF1",
    x"3D05BD38",
    x"3D05AC82",
    x"3D059BCD",
    x"3D058B1B",
    x"3D057A6A",
    x"3D0569BC",
    x"3D055910",
    x"3D054866",
    x"3D0537BE",
    x"3D052718",
    x"3D051674",
    x"3D0505D2",
    x"3D04F532",
    x"3D04E495",
    x"3D04D3F9",
    x"3D04C360",
    x"3D04B2C8",
    x"3D04A233",
    x"3D0491A0",
    x"3D04810F",
    x"3D047080",
    x"3D045FF3",
    x"3D044F68",
    x"3D043EDF",
    x"3D042E58",
    x"3D041DD3",
    x"3D040D50",
    x"3D03FCD0",
    x"3D03EC51",
    x"3D03DBD5",
    x"3D03CB5A",
    x"3D03BAE2",
    x"3D03AA6C",
    x"3D0399F7",
    x"3D038985",
    x"3D037915",
    x"3D0368A7",
    x"3D03583B",
    x"3D0347D1",
    x"3D033769",
    x"3D032703",
    x"3D03169F",
    x"3D03063D",
    x"3D02F5DE",
    x"3D02E580",
    x"3D02D524",
    x"3D02C4CB",
    x"3D02B473",
    x"3D02A41D",
    x"3D0293CA",
    x"3D028378",
    x"3D027329",
    x"3D0262DC",
    x"3D025290",
    x"3D024247",
    x"3D023200",
    x"3D0221BB",
    x"3D021177",
    x"3D020136",
    x"3D01F0F7",
    x"3D01E0BA",
    x"3D01D07F",
    x"3D01C046",
    x"3D01B00F",
    x"3D019FDA",
    x"3D018FA7",
    x"3D017F76",
    x"3D016F47",
    x"3D015F1A",
    x"3D014EEF",
    x"3D013EC6",
    x"3D012E9F",
    x"3D011E7B",
    x"3D010E58",
    x"3D00FE37",
    x"3D00EE18",
    x"3D00DDFC",
    x"3D00CDE1",
    x"3D00BDC8",
    x"3D00ADB1",
    x"3D009D9D",
    x"3D008D8A",
    x"3D007D79",
    x"3D006D6B",
    x"3D005D5E",
    x"3D004D53",
    x"3D003D4B",
    x"3D002D44",
    x"3D001D3F",
    x"3D000D3D",
    x"3CFFFA78",
    x"3CFFDA7B",
    x"3CFFBA81",
    x"3CFF9A8C",
    x"3CFF7A9B",
    x"3CFF5AAD",
    x"3CFF3AC4",
    x"3CFF1ADF",
    x"3CFEFAFD",
    x"3CFEDB20",
    x"3CFEBB46",
    x"3CFE9B71",
    x"3CFE7BA0",
    x"3CFE5BD2",
    x"3CFE3C09",
    x"3CFE1C43",
    x"3CFDFC82",
    x"3CFDDCC4",
    x"3CFDBD0A",
    x"3CFD9D55",
    x"3CFD7DA3",
    x"3CFD5DF5",
    x"3CFD3E4C",
    x"3CFD1EA6",
    x"3CFCFF04",
    x"3CFCDF66",
    x"3CFCBFCC",
    x"3CFCA036",
    x"3CFC80A4",
    x"3CFC6116",
    x"3CFC418C",
    x"3CFC2206",
    x"3CFC0283",
    x"3CFBE305",
    x"3CFBC38A",
    x"3CFBA414",
    x"3CFB84A1",
    x"3CFB6533",
    x"3CFB45C8",
    x"3CFB2661",
    x"3CFB06FF",
    x"3CFAE7A0",
    x"3CFAC845",
    x"3CFAA8EE",
    x"3CFA899A",
    x"3CFA6A4B",
    x"3CFA4B00",
    x"3CFA2BB8",
    x"3CFA0C75",
    x"3CF9ED35",
    x"3CF9CDFA",
    x"3CF9AEC2",
    x"3CF98F8E",
    x"3CF9705E",
    x"3CF95132",
    x"3CF9320A",
    x"3CF912E5",
    x"3CF8F3C5",
    x"3CF8D4A8",
    x"3CF8B590",
    x"3CF8967B",
    x"3CF8776A",
    x"3CF8585D",
    x"3CF83954",
    x"3CF81A4F",
    x"3CF7FB4D",
    x"3CF7DC50",
    x"3CF7BD56",
    x"3CF79E61",
    x"3CF77F6F",
    x"3CF76081",
    x"3CF74197",
    x"3CF722B0",
    x"3CF703CE",
    x"3CF6E4EF",
    x"3CF6C615",
    x"3CF6A73E",
    x"3CF6886B",
    x"3CF6699C",
    x"3CF64AD1",
    x"3CF62C09",
    x"3CF60D46",
    x"3CF5EE86",
    x"3CF5CFCA",
    x"3CF5B112",
    x"3CF5925E",
    x"3CF573AD",
    x"3CF55501",
    x"3CF53658",
    x"3CF517B3",
    x"3CF4F912",
    x"3CF4DA75",
    x"3CF4BBDB",
    x"3CF49D46",
    x"3CF47EB4",
    x"3CF46026",
    x"3CF4419C",
    x"3CF42316",
    x"3CF40493",
    x"3CF3E615",
    x"3CF3C79A",
    x"3CF3A923",
    x"3CF38AB0",
    x"3CF36C40",
    x"3CF34DD4",
    x"3CF32F6D",
    x"3CF31109",
    x"3CF2F2A8",
    x"3CF2D44C",
    x"3CF2B5F3",
    x"3CF2979E",
    x"3CF2794D",
    x"3CF25B00",
    x"3CF23CB7",
    x"3CF21E71",
    x"3CF2002F",
    x"3CF1E1F1",
    x"3CF1C3B7",
    x"3CF1A580",
    x"3CF1874D",
    x"3CF1691E",
    x"3CF14AF3",
    x"3CF12CCB",
    x"3CF10EA8",
    x"3CF0F088",
    x"3CF0D26C",
    x"3CF0B453",
    x"3CF0963E",
    x"3CF0782E",
    x"3CF05A20",
    x"3CF03C17",
    x"3CF01E11",
    x"3CF00010",
    x"3CEFE211",
    x"3CEFC417",
    x"3CEFA620",
    x"3CEF882D",
    x"3CEF6A3E",
    x"3CEF4C53",
    x"3CEF2E6B",
    x"3CEF1087",
    x"3CEEF2A7",
    x"3CEED4CB",
    x"3CEEB6F2",
    x"3CEE991D",
    x"3CEE7B4C",
    x"3CEE5D7E",
    x"3CEE3FB4",
    x"3CEE21EE",
    x"3CEE042C",
    x"3CEDE66D",
    x"3CEDC8B2",
    x"3CEDAAFB",
    x"3CED8D47",
    x"3CED6F98",
    x"3CED51EC",
    x"3CED3443",
    x"3CED169E",
    x"3CECF8FD",
    x"3CECDB60",
    x"3CECBDC7",
    x"3CECA031",
    x"3CEC829F",
    x"3CEC6510",
    x"3CEC4785",
    x"3CEC29FE",
    x"3CEC0C7B",
    x"3CEBEEFB",
    x"3CEBD17F",
    x"3CEBB407",
    x"3CEB9692",
    x"3CEB7921",
    x"3CEB5BB4",
    x"3CEB3E4A",
    x"3CEB20E4",
    x"3CEB0382",
    x"3CEAE623",
    x"3CEAC8C8",
    x"3CEAAB71",
    x"3CEA8E1E",
    x"3CEA70CE",
    x"3CEA5381",
    x"3CEA3639",
    x"3CEA18F4",
    x"3CE9FBB2",
    x"3CE9DE75",
    x"3CE9C13B",
    x"3CE9A405",
    x"3CE986D2",
    x"3CE969A3",
    x"3CE94C77",
    x"3CE92F50",
    x"3CE9122C",
    x"3CE8F50B",
    x"3CE8D7EE",
    x"3CE8BAD5",
    x"3CE89DC0",
    x"3CE880AE",
    x"3CE8639F",
    x"3CE84695",
    x"3CE8298E",
    x"3CE80C8A",
    x"3CE7EF8B",
    x"3CE7D28F",
    x"3CE7B596",
    x"3CE798A1",
    x"3CE77BB0",
    x"3CE75EC2",
    x"3CE741D8",
    x"3CE724F2",
    x"3CE7080F",
    x"3CE6EB30",
    x"3CE6CE54",
    x"3CE6B17C",
    x"3CE694A8",
    x"3CE677D7",
    x"3CE65B0A",
    x"3CE63E40",
    x"3CE6217A",
    x"3CE604B8",
    x"3CE5E7F9",
    x"3CE5CB3E",
    x"3CE5AE86",
    x"3CE591D2",
    x"3CE57522",
    x"3CE55875",
    x"3CE53BCC",
    x"3CE51F26",
    x"3CE50284",
    x"3CE4E5E5",
    x"3CE4C94A",
    x"3CE4ACB3",
    x"3CE4901F",
    x"3CE4738F",
    x"3CE45702",
    x"3CE43A79",
    x"3CE41DF4",
    x"3CE40172",
    x"3CE3E4F3",
    x"3CE3C879",
    x"3CE3AC01",
    x"3CE38F8E",
    x"3CE3731D",
    x"3CE356B1",
    x"3CE33A48",
    x"3CE31DE2",
    x"3CE30180",
    x"3CE2E522",
    x"3CE2C8C7",
    x"3CE2AC70",
    x"3CE2901C",
    x"3CE273CC",
    x"3CE2577F",
    x"3CE23B36",
    x"3CE21EF0",
    x"3CE202AE",
    x"3CE1E66F",
    x"3CE1CA34",
    x"3CE1ADFD",
    x"3CE191C9",
    x"3CE17598",
    x"3CE1596C",
    x"3CE13D42",
    x"3CE1211C",
    x"3CE104FA",
    x"3CE0E8DB",
    x"3CE0CCC0",
    x"3CE0B0A8",
    x"3CE09493",
    x"3CE07883",
    x"3CE05C75",
    x"3CE0406C",
    x"3CE02465",
    x"3CE00862",
    x"3CDFEC63",
    x"3CDFD067",
    x"3CDFB46F",
    x"3CDF987A",
    x"3CDF7C89",
    x"3CDF609B",
    x"3CDF44B1",
    x"3CDF28CA",
    x"3CDF0CE7",
    x"3CDEF107",
    x"3CDED52A",
    x"3CDEB951",
    x"3CDE9D7C",
    x"3CDE81AA",
    x"3CDE65DC",
    x"3CDE4A11",
    x"3CDE2E49",
    x"3CDE1285",
    x"3CDDF6C4",
    x"3CDDDB07",
    x"3CDDBF4E",
    x"3CDDA397",
    x"3CDD87E5",
    x"3CDD6C35",
    x"3CDD508A",
    x"3CDD34E1",
    x"3CDD193C",
    x"3CDCFD9B",
    x"3CDCE1FD",
    x"3CDCC663",
    x"3CDCAACB",
    x"3CDC8F38",
    x"3CDC73A8",
    x"3CDC581B",
    x"3CDC3C92",
    x"3CDC210C",
    x"3CDC0589",
    x"3CDBEA0A",
    x"3CDBCE8F",
    x"3CDBB317",
    x"3CDB97A2",
    x"3CDB7C31",
    x"3CDB60C3",
    x"3CDB4559",
    x"3CDB29F2",
    x"3CDB0E8E",
    x"3CDAF32E",
    x"3CDAD7D1",
    x"3CDABC78",
    x"3CDAA122",
    x"3CDA85D0",
    x"3CDA6A81",
    x"3CDA4F35",
    x"3CDA33ED",
    x"3CDA18A8",
    x"3CD9FD67",
    x"3CD9E229",
    x"3CD9C6EE",
    x"3CD9ABB7",
    x"3CD99083",
    x"3CD97553",
    x"3CD95A26",
    x"3CD93EFC",
    x"3CD923D6",
    x"3CD908B3",
    x"3CD8ED94",
    x"3CD8D278",
    x"3CD8B75F",
    x"3CD89C4A",
    x"3CD88138",
    x"3CD8662A",
    x"3CD84B1F",
    x"3CD83017",
    x"3CD81513",
    x"3CD7FA12",
    x"3CD7DF14",
    x"3CD7C41A",
    x"3CD7A923",
    x"3CD78E30",
    x"3CD77340",
    x"3CD75853",
    x"3CD73D6A",
    x"3CD72284",
    x"3CD707A1",
    x"3CD6ECC2",
    x"3CD6D1E6",
    x"3CD6B70D",
    x"3CD69C38",
    x"3CD68166",
    x"3CD66698",
    x"3CD64BCD",
    x"3CD63105",
    x"3CD61640",
    x"3CD5FB7F",
    x"3CD5E0C1",
    x"3CD5C607",
    x"3CD5AB50",
    x"3CD5909C",
    x"3CD575EC",
    x"3CD55B3F",
    x"3CD54095",
    x"3CD525EF",
    x"3CD50B4C",
    x"3CD4F0AC",
    x"3CD4D60F",
    x"3CD4BB76",
    x"3CD4A0E0",
    x"3CD4864E",
    x"3CD46BBF",
    x"3CD45133",
    x"3CD436AB",
    x"3CD41C25",
    x"3CD401A4",
    x"3CD3E725",
    x"3CD3CCAA",
    x"3CD3B232",
    x"3CD397BD",
    x"3CD37D4C",
    x"3CD362DE",
    x"3CD34873",
    x"3CD32E0C",
    x"3CD313A8",
    x"3CD2F947",
    x"3CD2DEE9",
    x"3CD2C48F",
    x"3CD2AA38",
    x"3CD28FE5",
    x"3CD27594",
    x"3CD25B47",
    x"3CD240FD",
    x"3CD226B7",
    x"3CD20C74",
    x"3CD1F234",
    x"3CD1D7F7",
    x"3CD1BDBE",
    x"3CD1A388",
    x"3CD18955",
    x"3CD16F25",
    x"3CD154F9",
    x"3CD13AD0",
    x"3CD120AA",
    x"3CD10688",
    x"3CD0EC69",
    x"3CD0D24D",
    x"3CD0B834",
    x"3CD09E1F",
    x"3CD0840D",
    x"3CD069FE",
    x"3CD04FF2",
    x"3CD035EA",
    x"3CD01BE5",
    x"3CD001E3",
    x"3CCFE7E4",
    x"3CCFCDE9",
    x"3CCFB3F1",
    x"3CCF99FC",
    x"3CCF800A",
    x"3CCF661C",
    x"3CCF4C31",
    x"3CCF3249",
    x"3CCF1864",
    x"3CCEFE83",
    x"3CCEE4A5",
    x"3CCECACA",
    x"3CCEB0F2",
    x"3CCE971D",
    x"3CCE7D4C",
    x"3CCE637E",
    x"3CCE49B3",
    x"3CCE2FEC",
    x"3CCE1627",
    x"3CCDFC66",
    x"3CCDE2A8",
    x"3CCDC8ED",
    x"3CCDAF36",
    x"3CCD9582",
    x"3CCD7BD1",
    x"3CCD6223",
    x"3CCD4878",
    x"3CCD2ED1",
    x"3CCD152C",
    x"3CCCFB8B",
    x"3CCCE1ED",
    x"3CCCC853",
    x"3CCCAEBB",
    x"3CCC9527",
    x"3CCC7B96",
    x"3CCC6208",
    x"3CCC487E",
    x"3CCC2EF6",
    x"3CCC1572",
    x"3CCBFBF1",
    x"3CCBE273",
    x"3CCBC8F8",
    x"3CCBAF81",
    x"3CCB960C",
    x"3CCB7C9B",
    x"3CCB632D",
    x"3CCB49C2",
    x"3CCB305B",
    x"3CCB16F6",
    x"3CCAFD95",
    x"3CCAE437",
    x"3CCACADC",
    x"3CCAB184",
    x"3CCA982F",
    x"3CCA7EDE",
    x"3CCA6590",
    x"3CCA4C45",
    x"3CCA32FD",
    x"3CCA19B8",
    x"3CCA0076",
    x"3CC9E738",
    x"3CC9CDFC",
    x"3CC9B4C4",
    x"3CC99B8F",
    x"3CC9825D",
    x"3CC9692F",
    x"3CC95003",
    x"3CC936DB",
    x"3CC91DB5",
    x"3CC90493",
    x"3CC8EB74",
    x"3CC8D258",
    x"3CC8B940",
    x"3CC8A02A",
    x"3CC88718",
    x"3CC86E08",
    x"3CC854FC",
    x"3CC83BF3",
    x"3CC822ED",
    x"3CC809EA",
    x"3CC7F0EB",
    x"3CC7D7EE",
    x"3CC7BEF5",
    x"3CC7A5FE",
    x"3CC78D0B",
    x"3CC7741B",
    x"3CC75B2E",
    x"3CC74244",
    x"3CC7295E",
    x"3CC7107A",
    x"3CC6F799",
    x"3CC6DEBC",
    x"3CC6C5E2",
    x"3CC6AD0B",
    x"3CC69436",
    x"3CC67B65",
    x"3CC66298",
    x"3CC649CD",
    x"3CC63105",
    x"3CC61841",
    x"3CC5FF7F",
    x"3CC5E6C1",
    x"3CC5CE05",
    x"3CC5B54D",
    x"3CC59C98",
    x"3CC583E6",
    x"3CC56B37",
    x"3CC5528B",
    x"3CC539E2",
    x"3CC5213D",
    x"3CC5089A",
    x"3CC4EFFB",
    x"3CC4D75E",
    x"3CC4BEC5",
    x"3CC4A62E",
    x"3CC48D9B",
    x"3CC4750B",
    x"3CC45C7E",
    x"3CC443F4",
    x"3CC42B6D",
    x"3CC412E9",
    x"3CC3FA68",
    x"3CC3E1EA",
    x"3CC3C970",
    x"3CC3B0F8",
    x"3CC39884",
    x"3CC38012",
    x"3CC367A4",
    x"3CC34F38",
    x"3CC336D0",
    x"3CC31E6A",
    x"3CC30608",
    x"3CC2EDA9",
    x"3CC2D54D",
    x"3CC2BCF4",
    x"3CC2A49D",
    x"3CC28C4A",
    x"3CC273FA",
    x"3CC25BAD",
    x"3CC24363",
    x"3CC22B1D",
    x"3CC212D9",
    x"3CC1FA98",
    x"3CC1E25A",
    x"3CC1CA1F",
    x"3CC1B1E8",
    x"3CC199B3",
    x"3CC18181",
    x"3CC16952",
    x"3CC15127",
    x"3CC138FE",
    x"3CC120D9",
    x"3CC108B6",
    x"3CC0F096",
    x"3CC0D87A",
    x"3CC0C060",
    x"3CC0A84A",
    x"3CC09036",
    x"3CC07826",
    x"3CC06018",
    x"3CC0480E",
    x"3CC03006",
    x"3CC01802",
    x"3CC00000",
    x"3CBFE802",
    x"3CBFD006",
    x"3CBFB80E",
    x"3CBFA018",
    x"3CBF8826",
    x"3CBF7036",
    x"3CBF5849",
    x"3CBF4060",
    x"3CBF2879",
    x"3CBF1096",
    x"3CBEF8B5",
    x"3CBEE0D8",
    x"3CBEC8FD",
    x"3CBEB125",
    x"3CBE9951",
    x"3CBE817F",
    x"3CBE69B0",
    x"3CBE51E5",
    x"3CBE3A1C",
    x"3CBE2256",
    x"3CBE0A93",
    x"3CBDF2D3",
    x"3CBDDB17",
    x"3CBDC35D",
    x"3CBDABA6",
    x"3CBD93F2",
    x"3CBD7C41",
    x"3CBD6493",
    x"3CBD4CE8",
    x"3CBD3540",
    x"3CBD1D9A",
    x"3CBD05F8",
    x"3CBCEE59",
    x"3CBCD6BD",
    x"3CBCBF23",
    x"3CBCA78D",
    x"3CBC8FF9",
    x"3CBC7869",
    x"3CBC60DB",
    x"3CBC4951",
    x"3CBC31C9",
    x"3CBC1A44",
    x"3CBC02C2",
    x"3CBBEB43",
    x"3CBBD3C7",
    x"3CBBBC4E",
    x"3CBBA4D8",
    x"3CBB8D65",
    x"3CBB75F5",
    x"3CBB5E88",
    x"3CBB471D",
    x"3CBB2FB6",
    x"3CBB1851",
    x"3CBB00F0",
    x"3CBAE991",
    x"3CBAD235",
    x"3CBABADD",
    x"3CBAA387",
    x"3CBA8C34",
    x"3CBA74E4",
    x"3CBA5D97",
    x"3CBA464C",
    x"3CBA2F05",
    x"3CBA17C1",
    x"3CBA007F",
    x"3CB9E940",
    x"3CB9D205",
    x"3CB9BACC",
    x"3CB9A396",
    x"3CB98C63",
    x"3CB97533",
    x"3CB95E06",
    x"3CB946DB",
    x"3CB92FB4",
    x"3CB91890",
    x"3CB9016E",
    x"3CB8EA4F",
    x"3CB8D333",
    x"3CB8BC1A",
    x"3CB8A504",
    x"3CB88DF1",
    x"3CB876E1",
    x"3CB85FD3",
    x"3CB848C9",
    x"3CB831C1",
    x"3CB81ABC",
    x"3CB803BB",
    x"3CB7ECBB",
    x"3CB7D5BF",
    x"3CB7BEC6",
    x"3CB7A7D0",
    x"3CB790DC",
    x"3CB779EB",
    x"3CB762FE",
    x"3CB74C13",
    x"3CB7352B",
    x"3CB71E45",
    x"3CB70763",
    x"3CB6F084",
    x"3CB6D9A7",
    x"3CB6C2CD",
    x"3CB6ABF6",
    x"3CB69522",
    x"3CB67E51",
    x"3CB66783",
    x"3CB650B7",
    x"3CB639EE",
    x"3CB62329",
    x"3CB60C66",
    x"3CB5F5A5",
    x"3CB5DEE8",
    x"3CB5C82E",
    x"3CB5B176",
    x"3CB59AC1",
    x"3CB5840F",
    x"3CB56D60",
    x"3CB556B4",
    x"3CB5400B",
    x"3CB52964",
    x"3CB512C0",
    x"3CB4FC1F",
    x"3CB4E581",
    x"3CB4CEE6",
    x"3CB4B84E",
    x"3CB4A1B8",
    x"3CB48B25",
    x"3CB47495",
    x"3CB45E08",
    x"3CB4477E",
    x"3CB430F6",
    x"3CB41A71",
    x"3CB403EF",
    x"3CB3ED70",
    x"3CB3D6F4",
    x"3CB3C07B",
    x"3CB3AA04",
    x"3CB39390",
    x"3CB37D1F",
    x"3CB366B1",
    x"3CB35045",
    x"3CB339DD",
    x"3CB32377",
    x"3CB30D14",
    x"3CB2F6B4",
    x"3CB2E056",
    x"3CB2C9FC",
    x"3CB2B3A4",
    x"3CB29D4F",
    x"3CB286FC",
    x"3CB270AD",
    x"3CB25A60",
    x"3CB24416",
    x"3CB22DCF",
    x"3CB2178B",
    x"3CB20149",
    x"3CB1EB0B",
    x"3CB1D4CF",
    x"3CB1BE95",
    x"3CB1A85F",
    x"3CB1922B",
    x"3CB17BFA",
    x"3CB165CC",
    x"3CB14FA1",
    x"3CB13978",
    x"3CB12353",
    x"3CB10D30",
    x"3CB0F70F",
    x"3CB0E0F2",
    x"3CB0CAD7",
    x"3CB0B4BF",
    x"3CB09EAA",
    x"3CB08897",
    x"3CB07288",
    x"3CB05C7B",
    x"3CB04671",
    x"3CB03069",
    x"3CB01A65",
    x"3CB00463",
    x"3CAFEE63",
    x"3CAFD867",
    x"3CAFC26D",
    x"3CAFAC76",
    x"3CAF9682",
    x"3CAF8091",
    x"3CAF6AA2",
    x"3CAF54B6",
    x"3CAF3ECD",
    x"3CAF28E6",
    x"3CAF1303",
    x"3CAEFD22",
    x"3CAEE743",
    x"3CAED168",
    x"3CAEBB8F",
    x"3CAEA5B9",
    x"3CAE8FE6",
    x"3CAE7A15",
    x"3CAE6447",
    x"3CAE4E7C",
    x"3CAE38B3",
    x"3CAE22EE",
    x"3CAE0D2B",
    x"3CADF76A",
    x"3CADE1AD",
    x"3CADCBF2",
    x"3CADB63A",
    x"3CADA084",
    x"3CAD8AD2",
    x"3CAD7522",
    x"3CAD5F74",
    x"3CAD49CA",
    x"3CAD3422",
    x"3CAD1E7D",
    x"3CAD08DA",
    x"3CACF33B",
    x"3CACDD9E",
    x"3CACC803",
    x"3CACB26C",
    x"3CAC9CD7",
    x"3CAC8744",
    x"3CAC71B5",
    x"3CAC5C28",
    x"3CAC469E",
    x"3CAC3116",
    x"3CAC1B91",
    x"3CAC060F",
    x"3CABF090",
    x"3CABDB13",
    x"3CABC599",
    x"3CABB022",
    x"3CAB9AAD",
    x"3CAB853B",
    x"3CAB6FCC",
    x"3CAB5A5F",
    x"3CAB44F5",
    x"3CAB2F8E",
    x"3CAB1A29",
    x"3CAB04C7",
    x"3CAAEF68",
    x"3CAADA0C",
    x"3CAAC4B2",
    x"3CAAAF5A",
    x"3CAA9A06",
    x"3CAA84B4",
    x"3CAA6F65",
    x"3CAA5A18",
    x"3CAA44CE",
    x"3CAA2F87",
    x"3CAA1A42",
    x"3CAA0500",
    x"3CA9EFC1",
    x"3CA9DA84",
    x"3CA9C54A",
    x"3CA9B013",
    x"3CA99ADE",
    x"3CA985AC",
    x"3CA9707D",
    x"3CA95B50",
    x"3CA94626",
    x"3CA930FF",
    x"3CA91BDA",
    x"3CA906B8",
    x"3CA8F198",
    x"3CA8DC7B",
    x"3CA8C761",
    x"3CA8B249",
    x"3CA89D34",
    x"3CA88822",
    x"3CA87312",
    x"3CA85E05",
    x"3CA848FB",
    x"3CA833F3",
    x"3CA81EEE",
    x"3CA809EB",
    x"3CA7F4EB",
    x"3CA7DFEE",
    x"3CA7CAF3",
    x"3CA7B5FB",
    x"3CA7A106",
    x"3CA78C13",
    x"3CA77723",
    x"3CA76235",
    x"3CA74D4A",
    x"3CA73862",
    x"3CA7237C",
    x"3CA70E99",
    x"3CA6F9B9",
    x"3CA6E4DB",
    x"3CA6CFFF",
    x"3CA6BB27",
    x"3CA6A651",
    x"3CA6917D",
    x"3CA67CAC",
    x"3CA667DE",
    x"3CA65312",
    x"3CA63E49",
    x"3CA62983",
    x"3CA614BF",
    x"3CA5FFFE",
    x"3CA5EB3F",
    x"3CA5D683",
    x"3CA5C1C9",
    x"3CA5AD12",
    x"3CA5985E",
    x"3CA583AC",
    x"3CA56EFD",
    x"3CA55A50",
    x"3CA545A6",
    x"3CA530FF",
    x"3CA51C5A",
    x"3CA507B8",
    x"3CA4F318",
    x"3CA4DE7B",
    x"3CA4C9E1",
    x"3CA4B549",
    x"3CA4A0B3",
    x"3CA48C21",
    x"3CA47790",
    x"3CA46303",
    x"3CA44E78",
    x"3CA439EF",
    x"3CA42569",
    x"3CA410E6",
    x"3CA3FC65",
    x"3CA3E7E7",
    x"3CA3D36B",
    x"3CA3BEF2",
    x"3CA3AA7B",
    x"3CA39607",
    x"3CA38196",
    x"3CA36D27",
    x"3CA358BA",
    x"3CA34451",
    x"3CA32FE9",
    x"3CA31B85",
    x"3CA30722",
    x"3CA2F2C3",
    x"3CA2DE66",
    x"3CA2CA0B",
    x"3CA2B5B3",
    x"3CA2A15E",
    x"3CA28D0B",
    x"3CA278BA",
    x"3CA2646D",
    x"3CA25021",
    x"3CA23BD9",
    x"3CA22792",
    x"3CA2134F",
    x"3CA1FF0E",
    x"3CA1EACF",
    x"3CA1D693",
    x"3CA1C259",
    x"3CA1AE22",
    x"3CA199EE",
    x"3CA185BC",
    x"3CA1718C",
    x"3CA15D5F",
    x"3CA14935",
    x"3CA1350D",
    x"3CA120E8",
    x"3CA10CC5",
    x"3CA0F8A5",
    x"3CA0E487",
    x"3CA0D06B",
    x"3CA0BC53",
    x"3CA0A83C",
    x"3CA09429",
    x"3CA08017",
    x"3CA06C09",
    x"3CA057FC",
    x"3CA043F3",
    x"3CA02FEB",
    x"3CA01BE7",
    x"3CA007E4",
    x"3C9FF3E5",
    x"3C9FDFE7",
    x"3C9FCBED",
    x"3C9FB7F4",
    x"3C9FA3FF",
    x"3C9F900B",
    x"3C9F7C1B",
    x"3C9F682C",
    x"3C9F5441",
    x"3C9F4057",
    x"3C9F2C71",
    x"3C9F188C",
    x"3C9F04AA",
    x"3C9EF0CB",
    x"3C9EDCEE",
    x"3C9EC914",
    x"3C9EB53C",
    x"3C9EA166",
    x"3C9E8D94",
    x"3C9E79C3",
    x"3C9E65F5",
    x"3C9E522A",
    x"3C9E3E61",
    x"3C9E2A9A",
    x"3C9E16D6",
    x"3C9E0314",
    x"3C9DEF55",
    x"3C9DDB98",
    x"3C9DC7DE",
    x"3C9DB426",
    x"3C9DA071",
    x"3C9D8CBE",
    x"3C9D790E",
    x"3C9D6560",
    x"3C9D51B5",
    x"3C9D3E0C",
    x"3C9D2A65",
    x"3C9D16C1",
    x"3C9D031F",
    x"3C9CEF80",
    x"3C9CDBE4",
    x"3C9CC849",
    x"3C9CB4B2",
    x"3C9CA11C",
    x"3C9C8D89",
    x"3C9C79F9",
    x"3C9C666B",
    x"3C9C52DF",
    x"3C9C3F56",
    x"3C9C2BCF",
    x"3C9C184B",
    x"3C9C04C9",
    x"3C9BF14A",
    x"3C9BDDCD",
    x"3C9BCA52",
    x"3C9BB6DA",
    x"3C9BA365",
    x"3C9B8FF2",
    x"3C9B7C81",
    x"3C9B6912",
    x"3C9B55A6",
    x"3C9B423D",
    x"3C9B2ED6",
    x"3C9B1B71",
    x"3C9B080F",
    x"3C9AF4AF",
    x"3C9AE152",
    x"3C9ACDF7",
    x"3C9ABA9E",
    x"3C9AA748",
    x"3C9A93F5",
    x"3C9A80A3",
    x"3C9A6D54",
    x"3C9A5A08",
    x"3C9A46BE",
    x"3C9A3376",
    x"3C9A2031",
    x"3C9A0CEE",
    x"3C99F9AE",
    x"3C99E670",
    x"3C99D334",
    x"3C99BFFB",
    x"3C99ACC4",
    x"3C999990",
    x"3C99865E",
    x"3C99732E",
    x"3C996001",
    x"3C994CD6",
    x"3C9939AE",
    x"3C992688",
    x"3C991364",
    x"3C990043",
    x"3C98ED24",
    x"3C98DA08",
    x"3C98C6EE",
    x"3C98B3D6",
    x"3C98A0C1",
    x"3C988DAE",
    x"3C987A9D",
    x"3C98678F",
    x"3C985483",
    x"3C98417A",
    x"3C982E73",
    x"3C981B6E",
    x"3C98086C",
    x"3C97F56C",
    x"3C97E26F",
    x"3C97CF74",
    x"3C97BC7B",
    x"3C97A985",
    x"3C979690",
    x"3C97839F",
    x"3C9770B0",
    x"3C975DC3",
    x"3C974AD8",
    x"3C9737F0",
    x"3C97250A",
    x"3C971227",
    x"3C96FF46",
    x"3C96EC67",
    x"3C96D98B",
    x"3C96C6B1",
    x"3C96B3D9",
    x"3C96A104",
    x"3C968E31",
    x"3C967B60",
    x"3C966892",
    x"3C9655C6",
    x"3C9642FC",
    x"3C963035",
    x"3C961D70",
    x"3C960AAE",
    x"3C95F7EE",
    x"3C95E530",
    x"3C95D274",
    x"3C95BFBB",
    x"3C95AD04",
    x"3C959A50",
    x"3C95879E",
    x"3C9574EE",
    x"3C956241",
    x"3C954F95",
    x"3C953CED",
    x"3C952A46",
    x"3C9517A2",
    x"3C950500",
    x"3C94F261",
    x"3C94DFC4",
    x"3C94CD29",
    x"3C94BA90",
    x"3C94A7FA",
    x"3C949566",
    x"3C9482D5",
    x"3C947046",
    x"3C945DB9",
    x"3C944B2E",
    x"3C9438A6",
    x"3C942620",
    x"3C94139D",
    x"3C94011B",
    x"3C93EE9C",
    x"3C93DC20",
    x"3C93C9A5",
    x"3C93B72D",
    x"3C93A4B7",
    x"3C939244",
    x"3C937FD3",
    x"3C936D64",
    x"3C935AF7",
    x"3C93488D",
    x"3C933625",
    x"3C9323C0",
    x"3C93115C",
    x"3C92FEFB",
    x"3C92EC9D",
    x"3C92DA40",
    x"3C92C7E6",
    x"3C92B58E",
    x"3C92A339",
    x"3C9290E5",
    x"3C927E94",
    x"3C926C46",
    x"3C9259F9",
    x"3C9247AF",
    x"3C923567",
    x"3C922322",
    x"3C9210DF",
    x"3C91FE9E",
    x"3C91EC5F",
    x"3C91DA23",
    x"3C91C7E9",
    x"3C91B5B1",
    x"3C91A37B",
    x"3C919148",
    x"3C917F17",
    x"3C916CE8",
    x"3C915ABC",
    x"3C914891",
    x"3C913669",
    x"3C912444",
    x"3C911220",
    x"3C90FFFF",
    x"3C90EDE0",
    x"3C90DBC4",
    x"3C90C9A9",
    x"3C90B791",
    x"3C90A57C",
    x"3C909368",
    x"3C908157",
    x"3C906F48",
    x"3C905D3B",
    x"3C904B30",
    x"3C903928",
    x"3C902722",
    x"3C90151E",
    x"3C90031D",
    x"3C8FF11D",
    x"3C8FDF20",
    x"3C8FCD26",
    x"3C8FBB2D",
    x"3C8FA937",
    x"3C8F9743",
    x"3C8F8551",
    x"3C8F7362",
    x"3C8F6174",
    x"3C8F4F89",
    x"3C8F3DA0",
    x"3C8F2BBA",
    x"3C8F19D5",
    x"3C8F07F3",
    x"3C8EF613",
    x"3C8EE436",
    x"3C8ED25A",
    x"3C8EC081",
    x"3C8EAEAA",
    x"3C8E9CD6",
    x"3C8E8B03",
    x"3C8E7933",
    x"3C8E6765",
    x"3C8E5599",
    x"3C8E43CF",
    x"3C8E3208",
    x"3C8E2043",
    x"3C8E0E80",
    x"3C8DFCBF",
    x"3C8DEB01",
    x"3C8DD944",
    x"3C8DC78A",
    x"3C8DB5D3",
    x"3C8DA41D",
    x"3C8D926A",
    x"3C8D80B8",
    x"3C8D6F09",
    x"3C8D5D5D",
    x"3C8D4BB2",
    x"3C8D3A0A",
    x"3C8D2864",
    x"3C8D16C0",
    x"3C8D051E",
    x"3C8CF37E",
    x"3C8CE1E1",
    x"3C8CD046",
    x"3C8CBEAD",
    x"3C8CAD16",
    x"3C8C9B82",
    x"3C8C89EF",
    x"3C8C785F",
    x"3C8C66D1",
    x"3C8C5545",
    x"3C8C43BC",
    x"3C8C3234",
    x"3C8C20AF",
    x"3C8C0F2C",
    x"3C8BFDAC",
    x"3C8BEC2D",
    x"3C8BDAB0",
    x"3C8BC936",
    x"3C8BB7BE",
    x"3C8BA648",
    x"3C8B94D5",
    x"3C8B8363",
    x"3C8B71F4",
    x"3C8B6087",
    x"3C8B4F1C",
    x"3C8B3DB3",
    x"3C8B2C4C",
    x"3C8B1AE8",
    x"3C8B0985",
    x"3C8AF825",
    x"3C8AE6C7",
    x"3C8AD56C",
    x"3C8AC412",
    x"3C8AB2BB",
    x"3C8AA165",
    x"3C8A9012",
    x"3C8A7EC1",
    x"3C8A6D73",
    x"3C8A5C26",
    x"3C8A4ADC",
    x"3C8A3993",
    x"3C8A284D",
    x"3C8A1709",
    x"3C8A05C7",
    x"3C89F488",
    x"3C89E34A",
    x"3C89D20F",
    x"3C89C0D6",
    x"3C89AF9F",
    x"3C899E6A",
    x"3C898D37",
    x"3C897C07",
    x"3C896AD8",
    x"3C8959AC",
    x"3C894882",
    x"3C89375A",
    x"3C892634",
    x"3C891510",
    x"3C8903EF",
    x"3C88F2CF",
    x"3C88E1B2",
    x"3C88D097",
    x"3C88BF7E",
    x"3C88AE67",
    x"3C889D52",
    x"3C888C40",
    x"3C887B2F",
    x"3C886A21",
    x"3C885915",
    x"3C88480B",
    x"3C883703",
    x"3C8825FD",
    x"3C8814F9",
    x"3C8803F8",
    x"3C87F2F8",
    x"3C87E1FB",
    x"3C87D100",
    x"3C87C007",
    x"3C87AF10",
    x"3C879E1B",
    x"3C878D28",
    x"3C877C37",
    x"3C876B49",
    x"3C875A5D",
    x"3C874972",
    x"3C87388A",
    x"3C8727A4",
    x"3C8716C0",
    x"3C8705DF",
    x"3C86F4FF",
    x"3C86E421",
    x"3C86D346",
    x"3C86C26D",
    x"3C86B195",
    x"3C86A0C0",
    x"3C868FED",
    x"3C867F1C",
    x"3C866E4D",
    x"3C865D81",
    x"3C864CB6",
    x"3C863BED",
    x"3C862B27",
    x"3C861A63",
    x"3C8609A0",
    x"3C85F8E0",
    x"3C85E822",
    x"3C85D766",
    x"3C85C6AC",
    x"3C85B5F4",
    x"3C85A53F",
    x"3C85948B",
    x"3C8583DA",
    x"3C85732A",
    x"3C85627D",
    x"3C8551D2",
    x"3C854128",
    x"3C853081",
    x"3C851FDC",
    x"3C850F39",
    x"3C84FE98",
    x"3C84EDFA",
    x"3C84DD5D",
    x"3C84CCC2",
    x"3C84BC2A",
    x"3C84AB93",
    x"3C849AFF",
    x"3C848A6D",
    x"3C8479DC",
    x"3C84694E",
    x"3C8458C2",
    x"3C844838",
    x"3C8437B0",
    x"3C84272A",
    x"3C8416A6",
    x"3C840624",
    x"3C83F5A5",
    x"3C83E527",
    x"3C83D4AB",
    x"3C83C432",
    x"3C83B3BA",
    x"3C83A345",
    x"3C8392D1",
    x"3C838260",
    x"3C8371F1",
    x"3C836184",
    x"3C835118",
    x"3C8340AF",
    x"3C833048",
    x"3C831FE3",
    x"3C830F80",
    x"3C82FF1F",
    x"3C82EEC1",
    x"3C82DE64",
    x"3C82CE09",
    x"3C82BDB0",
    x"3C82AD59",
    x"3C829D05",
    x"3C828CB2",
    x"3C827C62",
    x"3C826C13",
    x"3C825BC7",
    x"3C824B7C",
    x"3C823B34",
    x"3C822AED",
    x"3C821AA9",
    x"3C820A67",
    x"3C81FA26",
    x"3C81E9E8",
    x"3C81D9AC",
    x"3C81C972",
    x"3C81B93A",
    x"3C81A903",
    x"3C8198CF",
    x"3C81889D",
    x"3C81786D",
    x"3C81683F",
    x"3C815813",
    x"3C8147E9",
    x"3C8137C1",
    x"3C81279B",
    x"3C811777",
    x"3C810755",
    x"3C80F735",
    x"3C80E718",
    x"3C80D6FC",
    x"3C80C6E2",
    x"3C80B6CA",
    x"3C80A6B4",
    x"3C8096A0",
    x"3C80868E",
    x"3C80767F",
    x"3C806671",
    x"3C805665",
    x"3C80465B",
    x"3C803653",
    x"3C80264E",
    x"3C80164A",
    x"3C800648",
    x"3C7FEC91",
    x"3C7FCC95",
    x"3C7FAC9D",
    x"3C7F8CAA",
    x"3C7F6CBA",
    x"3C7F4CCF",
    x"3C7F2CE7",
    x"3C7F0D03",
    x"3C7EED24",
    x"3C7ECD48",
    x"3C7EAD70",
    x"3C7E8D9D",
    x"3C7E6DCD",
    x"3C7E4E01",
    x"3C7E2E3A",
    x"3C7E0E76",
    x"3C7DEEB6",
    x"3C7DCEFA",
    x"3C7DAF42",
    x"3C7D8F8E",
    x"3C7D6FDE",
    x"3C7D5032",
    x"3C7D308A",
    x"3C7D10E6",
    x"3C7CF146",
    x"3C7CD1AA",
    x"3C7CB212",
    x"3C7C927D",
    x"3C7C72ED",
    x"3C7C5361",
    x"3C7C33D8",
    x"3C7C1454",
    x"3C7BF4D3",
    x"3C7BD556",
    x"3C7BB5DE",
    x"3C7B9669",
    x"3C7B76F8",
    x"3C7B578B",
    x"3C7B3822",
    x"3C7B18BD",
    x"3C7AF95C",
    x"3C7AD9FF",
    x"3C7ABAA6",
    x"3C7A9B50",
    x"3C7A7BFF",
    x"3C7A5CB1",
    x"3C7A3D68",
    x"3C7A1E22",
    x"3C79FEE0",
    x"3C79DFA2",
    x"3C79C068",
    x"3C79A132",
    x"3C798200",
    x"3C7962D2",
    x"3C7943A7",
    x"3C792481",
    x"3C79055E",
    x"3C78E63F",
    x"3C78C724",
    x"3C78A80D",
    x"3C7888FA",
    x"3C7869EB",
    x"3C784AE0",
    x"3C782BD8",
    x"3C780CD5",
    x"3C77EDD5",
    x"3C77CED9",
    x"3C77AFE2",
    x"3C7790EE",
    x"3C7771FD",
    x"3C775311",
    x"3C773429",
    x"3C771544",
    x"3C76F663",
    x"3C76D786",
    x"3C76B8AD",
    x"3C7699D8",
    x"3C767B07",
    x"3C765C39",
    x"3C763D70",
    x"3C761EAA",
    x"3C75FFE8",
    x"3C75E12A",
    x"3C75C270",
    x"3C75A3BA",
    x"3C758507",
    x"3C756658",
    x"3C7547AD",
    x"3C752906",
    x"3C750A63",
    x"3C74EBC4",
    x"3C74CD28",
    x"3C74AE90",
    x"3C748FFD",
    x"3C74716C",
    x"3C7452E0",
    x"3C743458",
    x"3C7415D3",
    x"3C73F752",
    x"3C73D8D5",
    x"3C73BA5C",
    x"3C739BE7",
    x"3C737D75",
    x"3C735F07",
    x"3C73409D",
    x"3C732237",
    x"3C7303D5",
    x"3C72E576",
    x"3C72C71B",
    x"3C72A8C4",
    x"3C728A71",
    x"3C726C22",
    x"3C724DD6",
    x"3C722F8E",
    x"3C72114A",
    x"3C71F30A",
    x"3C71D4CE",
    x"3C71B695",
    x"3C719860",
    x"3C717A2F",
    x"3C715C01",
    x"3C713DD8",
    x"3C711FB2",
    x"3C710190",
    x"3C70E371",
    x"3C70C557",
    x"3C70A740",
    x"3C70892D",
    x"3C706B1E",
    x"3C704D12",
    x"3C702F0B",
    x"3C701107",
    x"3C6FF306",
    x"3C6FD50A",
    x"3C6FB711",
    x"3C6F991C",
    x"3C6F7B2B",
    x"3C6F5D3D",
    x"3C6F3F53",
    x"3C6F216D",
    x"3C6F038B",
    x"3C6EE5AD",
    x"3C6EC7D2",
    x"3C6EA9FB",
    x"3C6E8C27",
    x"3C6E6E58",
    x"3C6E508C",
    x"3C6E32C3",
    x"3C6E14FF",
    x"3C6DF73E",
    x"3C6DD981",
    x"3C6DBBC8",
    x"3C6D9E12",
    x"3C6D8060",
    x"3C6D62B2",
    x"3C6D4508",
    x"3C6D2761",
    x"3C6D09BE",
    x"3C6CEC1E",
    x"3C6CCE83",
    x"3C6CB0EB",
    x"3C6C9356",
    x"3C6C75C6",
    x"3C6C5839",
    x"3C6C3AB0",
    x"3C6C1D2A",
    x"3C6BFFA9",
    x"3C6BE22A",
    x"3C6BC4B0",
    x"3C6BA739",
    x"3C6B89C6",
    x"3C6B6C57",
    x"3C6B4EEB",
    x"3C6B3183",
    x"3C6B141F",
    x"3C6AF6BE",
    x"3C6AD961",
    x"3C6ABC08",
    x"3C6A9EB2",
    x"3C6A8160",
    x"3C6A6412",
    x"3C6A46C7",
    x"3C6A2980",
    x"3C6A0C3D",
    x"3C69EEFD",
    x"3C69D1C1",
    x"3C69B489",
    x"3C699754",
    x"3C697A23",
    x"3C695CF5",
    x"3C693FCB",
    x"3C6922A5",
    x"3C690583",
    x"3C68E864",
    x"3C68CB49",
    x"3C68AE31",
    x"3C68911D",
    x"3C68740D",
    x"3C685700",
    x"3C6839F7",
    x"3C681CF2",
    x"3C67FFF0",
    x"3C67E2F2",
    x"3C67C5F7",
    x"3C67A900",
    x"3C678C0D",
    x"3C676F1D",
    x"3C675231",
    x"3C673549",
    x"3C671864",
    x"3C66FB83",
    x"3C66DEA5",
    x"3C66C1CB",
    x"3C66A4F4",
    x"3C668822",
    x"3C666B52",
    x"3C664E87",
    x"3C6631BF",
    x"3C6614FA",
    x"3C65F83A",
    x"3C65DB7C",
    x"3C65BEC3",
    x"3C65A20D",
    x"3C65855A",
    x"3C6568AB",
    x"3C654C00",
    x"3C652F58",
    x"3C6512B4",
    x"3C64F614",
    x"3C64D977",
    x"3C64BCDD",
    x"3C64A047",
    x"3C6483B5",
    x"3C646726",
    x"3C644A9B",
    x"3C642E14",
    x"3C641190",
    x"3C63F50F",
    x"3C63D893",
    x"3C63BC19",
    x"3C639FA4",
    x"3C638331",
    x"3C6366C3",
    x"3C634A58",
    x"3C632DF0",
    x"3C63118C",
    x"3C62F52C",
    x"3C62D8CF",
    x"3C62BC76",
    x"3C62A020",
    x"3C6283CE",
    x"3C62677F",
    x"3C624B34",
    x"3C622EEC",
    x"3C6212A8",
    x"3C61F667",
    x"3C61DA2A",
    x"3C61BDF1",
    x"3C61A1BB",
    x"3C618588",
    x"3C616959",
    x"3C614D2E",
    x"3C613106",
    x"3C6114E2",
    x"3C60F8C1",
    x"3C60DCA4",
    x"3C60C08A",
    x"3C60A473",
    x"3C608861",
    x"3C606C51",
    x"3C605046",
    x"3C60343D",
    x"3C601839",
    x"3C5FFC37",
    x"3C5FE039",
    x"3C5FC43F",
    x"3C5FA848",
    x"3C5F8C55",
    x"3C5F7065",
    x"3C5F5479",
    x"3C5F3890",
    x"3C5F1CAB",
    x"3C5F00C9",
    x"3C5EE4EB",
    x"3C5EC910",
    x"3C5EAD38",
    x"3C5E9165",
    x"3C5E7594",
    x"3C5E59C7",
    x"3C5E3DFE",
    x"3C5E2238",
    x"3C5E0675",
    x"3C5DEAB6",
    x"3C5DCEFA",
    x"3C5DB342",
    x"3C5D978E",
    x"3C5D7BDC",
    x"3C5D602F",
    x"3C5D4484",
    x"3C5D28DD",
    x"3C5D0D3A",
    x"3C5CF19A",
    x"3C5CD5FE",
    x"3C5CBA65",
    x"3C5C9ECF",
    x"3C5C833D",
    x"3C5C67AE",
    x"3C5C4C23",
    x"3C5C309B",
    x"3C5C1517",
    x"3C5BF996",
    x"3C5BDE19",
    x"3C5BC29E",
    x"3C5BA728",
    x"3C5B8BB5",
    x"3C5B7045",
    x"3C5B54D9",
    x"3C5B3970",
    x"3C5B1E0A",
    x"3C5B02A8",
    x"3C5AE74A",
    x"3C5ACBEE",
    x"3C5AB097",
    x"3C5A9542",
    x"3C5A79F1",
    x"3C5A5EA4",
    x"3C5A435A",
    x"3C5A2813",
    x"3C5A0CD0",
    x"3C59F190",
    x"3C59D653",
    x"3C59BB1A",
    x"3C599FE4",
    x"3C5984B2",
    x"3C596983",
    x"3C594E58",
    x"3C593330",
    x"3C59180B",
    x"3C58FCEA",
    x"3C58E1CC",
    x"3C58C6B1",
    x"3C58AB9A",
    x"3C589086",
    x"3C587576",
    x"3C585A69",
    x"3C583F5F",
    x"3C582459",
    x"3C580956",
    x"3C57EE57",
    x"3C57D35B",
    x"3C57B862",
    x"3C579D6D",
    x"3C57827B",
    x"3C57678C",
    x"3C574CA1",
    x"3C5731B9",
    x"3C5716D4",
    x"3C56FBF3",
    x"3C56E115",
    x"3C56C63B",
    x"3C56AB64",
    x"3C569090",
    x"3C5675C0",
    x"3C565AF3",
    x"3C564029",
    x"3C562562",
    x"3C560A9F",
    x"3C55EFE0",
    x"3C55D524",
    x"3C55BA6B",
    x"3C559FB5",
    x"3C558503",
    x"3C556A54",
    x"3C554FA8",
    x"3C553500",
    x"3C551A5B",
    x"3C54FFB9",
    x"3C54E51B",
    x"3C54CA80",
    x"3C54AFE8",
    x"3C549554",
    x"3C547AC3",
    x"3C546035",
    x"3C5445AB",
    x"3C542B24",
    x"3C5410A0",
    x"3C53F620",
    x"3C53DBA3",
    x"3C53C129",
    x"3C53A6B2",
    x"3C538C3F",
    x"3C5371CF",
    x"3C535763",
    x"3C533CF9",
    x"3C532293",
    x"3C530831",
    x"3C52EDD1",
    x"3C52D375",
    x"3C52B91C",
    x"3C529EC7",
    x"3C528475",
    x"3C526A26",
    x"3C524FDA",
    x"3C523592",
    x"3C521B4D",
    x"3C52010B",
    x"3C51E6CD",
    x"3C51CC91",
    x"3C51B259",
    x"3C519825",
    x"3C517DF3",
    x"3C5163C5",
    x"3C51499A",
    x"3C512F73",
    x"3C51154F",
    x"3C50FB2E",
    x"3C50E110",
    x"3C50C6F5",
    x"3C50ACDE",
    x"3C5092CA",
    x"3C5078B9",
    x"3C505EAC",
    x"3C5044A2",
    x"3C502A9B",
    x"3C501097",
    x"3C4FF697",
    x"3C4FDC99",
    x"3C4FC29F",
    x"3C4FA8A9",
    x"3C4F8EB5",
    x"3C4F74C5",
    x"3C4F5AD8",
    x"3C4F40EE",
    x"3C4F2708",
    x"3C4F0D25",
    x"3C4EF345",
    x"3C4ED968",
    x"3C4EBF8E",
    x"3C4EA5B8",
    x"3C4E8BE5",
    x"3C4E7215",
    x"3C4E5848",
    x"3C4E3E7F",
    x"3C4E24B9",
    x"3C4E0AF6",
    x"3C4DF136",
    x"3C4DD779",
    x"3C4DBDC0",
    x"3C4DA40A",
    x"3C4D8A57",
    x"3C4D70A7",
    x"3C4D56FB",
    x"3C4D3D52",
    x"3C4D23AB",
    x"3C4D0A09",
    x"3C4CF069",
    x"3C4CD6CD",
    x"3C4CBD33",
    x"3C4CA39D",
    x"3C4C8A0A",
    x"3C4C707B",
    x"3C4C56EE",
    x"3C4C3D65",
    x"3C4C23DF",
    x"3C4C0A5C",
    x"3C4BF0DC",
    x"3C4BD760",
    x"3C4BBDE6",
    x"3C4BA470",
    x"3C4B8AFD",
    x"3C4B718E",
    x"3C4B5821",
    x"3C4B3EB8",
    x"3C4B2551",
    x"3C4B0BEE",
    x"3C4AF28E",
    x"3C4AD932",
    x"3C4ABFD8",
    x"3C4AA682",
    x"3C4A8D2E",
    x"3C4A73DE",
    x"3C4A5A91",
    x"3C4A4148",
    x"3C4A2801",
    x"3C4A0EBE",
    x"3C49F57D",
    x"3C49DC40",
    x"3C49C306",
    x"3C49A9D0",
    x"3C49909C",
    x"3C49776B",
    x"3C495E3E",
    x"3C494514",
    x"3C492BED",
    x"3C4912C9",
    x"3C48F9A8",
    x"3C48E08A",
    x"3C48C770",
    x"3C48AE59",
    x"3C489544",
    x"3C487C33",
    x"3C486325",
    x"3C484A1A",
    x"3C483113",
    x"3C48180E",
    x"3C47FF0D",
    x"3C47E60E",
    x"3C47CD13",
    x"3C47B41B",
    x"3C479B26",
    x"3C478234",
    x"3C476946",
    x"3C47505A",
    x"3C473772",
    x"3C471E8C",
    x"3C4705AA",
    x"3C46ECCB",
    x"3C46D3EF",
    x"3C46BB16",
    x"3C46A240",
    x"3C46896D",
    x"3C46709E",
    x"3C4657D1",
    x"3C463F08",
    x"3C462641",
    x"3C460D7E",
    x"3C45F4BE",
    x"3C45DC01",
    x"3C45C347",
    x"3C45AA90",
    x"3C4591DC",
    x"3C45792C",
    x"3C45607E",
    x"3C4547D4",
    x"3C452F2C",
    x"3C451688",
    x"3C44FDE6",
    x"3C44E548",
    x"3C44CCAD",
    x"3C44B415",
    x"3C449B80",
    x"3C4482EE",
    x"3C446A5F",
    x"3C4451D4",
    x"3C44394B",
    x"3C4420C5",
    x"3C440843",
    x"3C43EFC3",
    x"3C43D747",
    x"3C43BECD",
    x"3C43A657",
    x"3C438DE4",
    x"3C437574",
    x"3C435D06",
    x"3C43449C",
    x"3C432C35",
    x"3C4313D1",
    x"3C42FB70",
    x"3C42E312",
    x"3C42CAB8",
    x"3C42B260",
    x"3C429A0B",
    x"3C4281B9",
    x"3C42696B",
    x"3C42511F",
    x"3C4238D6",
    x"3C422091",
    x"3C42084E",
    x"3C41F00F",
    x"3C41D7D2",
    x"3C41BF99",
    x"3C41A762",
    x"3C418F2F",
    x"3C4176FE",
    x"3C415ED1",
    x"3C4146A7",
    x"3C412E7F",
    x"3C41165B",
    x"3C40FE3A",
    x"3C40E61C",
    x"3C40CE00",
    x"3C40B5E8",
    x"3C409DD3",
    x"3C4085C1",
    x"3C406DB1",
    x"3C4055A5",
    x"3C403D9C",
    x"3C402596",
    x"3C400D93",
    x"3C3FF592",
    x"3C3FDD95",
    x"3C3FC59B",
    x"3C3FADA4",
    x"3C3F95B0",
    x"3C3F7DBE",
    x"3C3F65D0",
    x"3C3F4DE5",
    x"3C3F35FD",
    x"3C3F1E17",
    x"3C3F0635",
    x"3C3EEE56",
    x"3C3ED67A",
    x"3C3EBEA0",
    x"3C3EA6CA",
    x"3C3E8EF7",
    x"3C3E7726",
    x"3C3E5F59",
    x"3C3E478E",
    x"3C3E2FC7",
    x"3C3E1802",
    x"3C3E0041",
    x"3C3DE882",
    x"3C3DD0C7",
    x"3C3DB90E",
    x"3C3DA158",
    x"3C3D89A6",
    x"3C3D71F6",
    x"3C3D5A49",
    x"3C3D429F",
    x"3C3D2AF9",
    x"3C3D1355",
    x"3C3CFBB4",
    x"3C3CE416",
    x"3C3CCC7B",
    x"3C3CB4E3",
    x"3C3C9D4E",
    x"3C3C85BB",
    x"3C3C6E2C",
    x"3C3C56A0",
    x"3C3C3F16",
    x"3C3C2790",
    x"3C3C100D",
    x"3C3BF88C",
    x"3C3BE10E",
    x"3C3BC994",
    x"3C3BB21C",
    x"3C3B9AA7",
    x"3C3B8335",
    x"3C3B6BC6",
    x"3C3B545A",
    x"3C3B3CF1",
    x"3C3B258B",
    x"3C3B0E28",
    x"3C3AF6C8",
    x"3C3ADF6A",
    x"3C3AC810",
    x"3C3AB0B8",
    x"3C3A9964",
    x"3C3A8212",
    x"3C3A6AC3",
    x"3C3A5377",
    x"3C3A3C2E",
    x"3C3A24E8",
    x"3C3A0DA5",
    x"3C39F665",
    x"3C39DF27",
    x"3C39C7ED",
    x"3C39B0B5",
    x"3C399981",
    x"3C39824F",
    x"3C396B20",
    x"3C3953F4",
    x"3C393CCB",
    x"3C3925A5",
    x"3C390E82",
    x"3C38F761",
    x"3C38E044",
    x"3C38C929",
    x"3C38B212",
    x"3C389AFD",
    x"3C3883EB",
    x"3C386CDC",
    x"3C3855D0",
    x"3C383EC6",
    x"3C3827C0",
    x"3C3810BC",
    x"3C37F9BC",
    x"3C37E2BE",
    x"3C37CBC3",
    x"3C37B4CB",
    x"3C379DD6",
    x"3C3786E4",
    x"3C376FF4",
    x"3C375908",
    x"3C37421E",
    x"3C372B37",
    x"3C371453",
    x"3C36FD72",
    x"3C36E694",
    x"3C36CFB8",
    x"3C36B8E0",
    x"3C36A20A",
    x"3C368B37",
    x"3C367467",
    x"3C365D9A",
    x"3C3646D0",
    x"3C363009",
    x"3C361944",
    x"3C360282",
    x"3C35EBC3",
    x"3C35D507",
    x"3C35BE4E",
    x"3C35A798",
    x"3C3590E4",
    x"3C357A33",
    x"3C356386",
    x"3C354CDB",
    x"3C353632",
    x"3C351F8D",
    x"3C3508EB",
    x"3C34F24B",
    x"3C34DBAE",
    x"3C34C514",
    x"3C34AE7D",
    x"3C3497E8",
    x"3C348157",
    x"3C346AC8",
    x"3C34543C",
    x"3C343DB3",
    x"3C34272D",
    x"3C3410A9",
    x"3C33FA28",
    x"3C33E3AB",
    x"3C33CD2F",
    x"3C33B6B7",
    x"3C33A042",
    x"3C3389CF",
    x"3C33735F",
    x"3C335CF2",
    x"3C334688",
    x"3C333021",
    x"3C3319BC",
    x"3C33035A",
    x"3C32ECFB",
    x"3C32D69F",
    x"3C32C046",
    x"3C32A9EF",
    x"3C32939B",
    x"3C327D4A",
    x"3C3266FC",
    x"3C3250B0",
    x"3C323A68",
    x"3C322422",
    x"3C320DDF",
    x"3C31F79E",
    x"3C31E161",
    x"3C31CB26",
    x"3C31B4EE",
    x"3C319EB9",
    x"3C318886",
    x"3C317257",
    x"3C315C2A",
    x"3C3145FF",
    x"3C312FD8",
    x"3C3119B4",
    x"3C310392",
    x"3C30ED73",
    x"3C30D756",
    x"3C30C13D",
    x"3C30AB26",
    x"3C309512",
    x"3C307F01",
    x"3C3068F2",
    x"3C3052E7",
    x"3C303CDE",
    x"3C3026D7",
    x"3C3010D4",
    x"3C2FFAD3",
    x"3C2FE4D5",
    x"3C2FCEDA",
    x"3C2FB8E1",
    x"3C2FA2EC",
    x"3C2F8CF9",
    x"3C2F7708",
    x"3C2F611B",
    x"3C2F4B30",
    x"3C2F3548",
    x"3C2F1F63",
    x"3C2F0980",
    x"3C2EF3A0",
    x"3C2EDDC3",
    x"3C2EC7E9",
    x"3C2EB211",
    x"3C2E9C3C",
    x"3C2E866A",
    x"3C2E709B",
    x"3C2E5ACE",
    x"3C2E4504",
    x"3C2E2F3D",
    x"3C2E1978",
    x"3C2E03B7",
    x"3C2DEDF7",
    x"3C2DD83B",
    x"3C2DC281",
    x"3C2DACCA",
    x"3C2D9716",
    x"3C2D8165",
    x"3C2D6BB6",
    x"3C2D560A",
    x"3C2D4060",
    x"3C2D2ABA",
    x"3C2D1516",
    x"3C2CFF74",
    x"3C2CE9D6",
    x"3C2CD43A",
    x"3C2CBEA1",
    x"3C2CA90A",
    x"3C2C9376",
    x"3C2C7DE5",
    x"3C2C6857",
    x"3C2C52CB",
    x"3C2C3D42",
    x"3C2C27BC",
    x"3C2C1238",
    x"3C2BFCB7",
    x"3C2BE739",
    x"3C2BD1BE",
    x"3C2BBC45",
    x"3C2BA6CF",
    x"3C2B915B",
    x"3C2B7BEA",
    x"3C2B667C",
    x"3C2B5111",
    x"3C2B3BA8",
    x"3C2B2642",
    x"3C2B10DE",
    x"3C2AFB7D",
    x"3C2AE61F",
    x"3C2AD0C4",
    x"3C2ABB6B",
    x"3C2AA615",
    x"3C2A90C2",
    x"3C2A7B71",
    x"3C2A6623",
    x"3C2A50D7",
    x"3C2A3B8F",
    x"3C2A2648",
    x"3C2A1105",
    x"3C29FBC4",
    x"3C29E686",
    x"3C29D14B",
    x"3C29BC12",
    x"3C29A6DC",
    x"3C2991A8",
    x"3C297C77",
    x"3C296749",
    x"3C29521D",
    x"3C293CF4",
    x"3C2927CE",
    x"3C2912AA",
    x"3C28FD89",
    x"3C28E86B",
    x"3C28D34F",
    x"3C28BE36",
    x"3C28A920",
    x"3C28940C",
    x"3C287EFB",
    x"3C2869EC",
    x"3C2854E0",
    x"3C283FD7",
    x"3C282AD0",
    x"3C2815CC",
    x"3C2800CB",
    x"3C27EBCC",
    x"3C27D6D0",
    x"3C27C1D6",
    x"3C27ACDF",
    x"3C2797EB",
    x"3C2782F9",
    x"3C276E0A",
    x"3C27591E",
    x"3C274434",
    x"3C272F4D",
    x"3C271A68",
    x"3C270586",
    x"3C26F0A7",
    x"3C26DBCA",
    x"3C26C6F0",
    x"3C26B218",
    x"3C269D43",
    x"3C268871",
    x"3C2673A1",
    x"3C265ED4",
    x"3C264A0A",
    x"3C263542",
    x"3C26207C",
    x"3C260BBA",
    x"3C25F6F9",
    x"3C25E23C",
    x"3C25CD81",
    x"3C25B8C8",
    x"3C25A413",
    x"3C258F5F",
    x"3C257AAF",
    x"3C256601",
    x"3C255155",
    x"3C253CAC",
    x"3C252806",
    x"3C251362",
    x"3C24FEC1",
    x"3C24EA23",
    x"3C24D587",
    x"3C24C0ED",
    x"3C24AC56",
    x"3C2497C2",
    x"3C248331",
    x"3C246EA1",
    x"3C245A15",
    x"3C24458B",
    x"3C243104",
    x"3C241C7F",
    x"3C2407FC",
    x"3C23F37D",
    x"3C23DF00",
    x"3C23CA85",
    x"3C23B60D",
    x"3C23A197",
    x"3C238D24",
    x"3C2378B4",
    x"3C236446",
    x"3C234FDB",
    x"3C233B72",
    x"3C23270C",
    x"3C2312A9",
    x"3C22FE48",
    x"3C22E9E9",
    x"3C22D58D",
    x"3C22C134",
    x"3C22ACDD",
    x"3C229888",
    x"3C228437",
    x"3C226FE7",
    x"3C225B9B",
    x"3C224750",
    x"3C223309",
    x"3C221EC4",
    x"3C220A81",
    x"3C21F641",
    x"3C21E204",
    x"3C21CDC9",
    x"3C21B990",
    x"3C21A55A",
    x"3C219127",
    x"3C217CF6",
    x"3C2168C8",
    x"3C21549C",
    x"3C214072",
    x"3C212C4C",
    x"3C211827",
    x"3C210406",
    x"3C20EFE6",
    x"3C20DBCA",
    x"3C20C7AF",
    x"3C20B398",
    x"3C209F82",
    x"3C208B70",
    x"3C207760",
    x"3C206352",
    x"3C204F47",
    x"3C203B3E",
    x"3C202738",
    x"3C201334",
    x"3C1FFF33",
    x"3C1FEB34",
    x"3C1FD738",
    x"3C1FC33F",
    x"3C1FAF48",
    x"3C1F9B53",
    x"3C1F8761",
    x"3C1F7371",
    x"3C1F5F84",
    x"3C1F4B99",
    x"3C1F37B1",
    x"3C1F23CB",
    x"3C1F0FE8",
    x"3C1EFC07",
    x"3C1EE829",
    x"3C1ED44D",
    x"3C1EC074",
    x"3C1EAC9D",
    x"3C1E98C9",
    x"3C1E84F7",
    x"3C1E7128",
    x"3C1E5D5B",
    x"3C1E4990",
    x"3C1E35C8",
    x"3C1E2203",
    x"3C1E0E40",
    x"3C1DFA7F",
    x"3C1DE6C1",
    x"3C1DD305",
    x"3C1DBF4C",
    x"3C1DAB96",
    x"3C1D97E1",
    x"3C1D8430",
    x"3C1D7080",
    x"3C1D5CD4",
    x"3C1D4929",
    x"3C1D3581",
    x"3C1D21DC",
    x"3C1D0E39",
    x"3C1CFA98",
    x"3C1CE6FA",
    x"3C1CD35E",
    x"3C1CBFC5",
    x"3C1CAC2F",
    x"3C1C989A",
    x"3C1C8508",
    x"3C1C7179",
    x"3C1C5DEC",
    x"3C1C4A62",
    x"3C1C36D9",
    x"3C1C2354",
    x"3C1C0FD1",
    x"3C1BFC50",
    x"3C1BE8D2",
    x"3C1BD556",
    x"3C1BC1DC",
    x"3C1BAE65",
    x"3C1B9AF1",
    x"3C1B877E",
    x"3C1B740F",
    x"3C1B60A1",
    x"3C1B4D37",
    x"3C1B39CE",
    x"3C1B2668",
    x"3C1B1305",
    x"3C1AFFA3",
    x"3C1AEC45",
    x"3C1AD8E8",
    x"3C1AC58E",
    x"3C1AB237",
    x"3C1A9EE2",
    x"3C1A8B8F",
    x"3C1A783F",
    x"3C1A64F1",
    x"3C1A51A6",
    x"3C1A3E5D",
    x"3C1A2B16",
    x"3C1A17D2",
    x"3C1A0490",
    x"3C19F151",
    x"3C19DE14",
    x"3C19CAD9",
    x"3C19B7A1",
    x"3C19A46B",
    x"3C199138",
    x"3C197E07",
    x"3C196AD9",
    x"3C1957AC",
    x"3C194483",
    x"3C19315B",
    x"3C191E36",
    x"3C190B14",
    x"3C18F7F3",
    x"3C18E4D6",
    x"3C18D1BA",
    x"3C18BEA1",
    x"3C18AB8B",
    x"3C189876",
    x"3C188564",
    x"3C187255",
    x"3C185F48",
    x"3C184C3D",
    x"3C183935",
    x"3C18262F",
    x"3C18132B",
    x"3C18002A",
    x"3C17ED2B",
    x"3C17DA2F",
    x"3C17C735",
    x"3C17B43D",
    x"3C17A148",
    x"3C178E55",
    x"3C177B64",
    x"3C176876",
    x"3C17558A",
    x"3C1742A0",
    x"3C172FB9",
    x"3C171CD5",
    x"3C1709F2",
    x"3C16F712",
    x"3C16E434",
    x"3C16D159",
    x"3C16BE80",
    x"3C16ABA9",
    x"3C1698D5",
    x"3C168603",
    x"3C167334",
    x"3C166066",
    x"3C164D9B",
    x"3C163AD3",
    x"3C16280D",
    x"3C161549",
    x"3C160287",
    x"3C15EFC8",
    x"3C15DD0B",
    x"3C15CA51",
    x"3C15B799",
    x"3C15A4E3",
    x"3C159230",
    x"3C157F7F",
    x"3C156CD0",
    x"3C155A23",
    x"3C154779",
    x"3C1534D2",
    x"3C15222C",
    x"3C150F89",
    x"3C14FCE8",
    x"3C14EA4A",
    x"3C14D7AE",
    x"3C14C514",
    x"3C14B27C",
    x"3C149FE7",
    x"3C148D54",
    x"3C147AC4",
    x"3C146836",
    x"3C1455AA",
    x"3C144320",
    x"3C143099",
    x"3C141E14",
    x"3C140B92",
    x"3C13F911",
    x"3C13E693",
    x"3C13D418",
    x"3C13C19E",
    x"3C13AF27",
    x"3C139CB2",
    x"3C138A40",
    x"3C1377D0",
    x"3C136562",
    x"3C1352F7",
    x"3C13408D",
    x"3C132E26",
    x"3C131BC2",
    x"3C13095F",
    x"3C12F6FF",
    x"3C12E4A2",
    x"3C12D246",
    x"3C12BFED",
    x"3C12AD96",
    x"3C129B42",
    x"3C1288EF",
    x"3C12769F",
    x"3C126452",
    x"3C125206",
    x"3C123FBD",
    x"3C122D76",
    x"3C121B32",
    x"3C1208F0",
    x"3C11F6B0",
    x"3C11E472",
    x"3C11D237",
    x"3C11BFFD",
    x"3C11ADC7",
    x"3C119B92",
    x"3C118960",
    x"3C117730",
    x"3C116502",
    x"3C1152D6",
    x"3C1140AD",
    x"3C112E86",
    x"3C111C62",
    x"3C110A3F",
    x"3C10F81F",
    x"3C10E601",
    x"3C10D3E6",
    x"3C10C1CC",
    x"3C10AFB5",
    x"3C109DA0",
    x"3C108B8E",
    x"3C10797D",
    x"3C10676F",
    x"3C105563",
    x"3C10435A",
    x"3C103153",
    x"3C101F4E",
    x"3C100D4B",
    x"3C0FFB4A",
    x"3C0FE94C",
    x"3C0FD750",
    x"3C0FC556",
    x"3C0FB35F",
    x"3C0FA169",
    x"3C0F8F76",
    x"3C0F7D85",
    x"3C0F6B97",
    x"3C0F59AB",
    x"3C0F47C0",
    x"3C0F35D9",
    x"3C0F23F3",
    x"3C0F1210",
    x"3C0F002E",
    x"3C0EEE50",
    x"3C0EDC73",
    x"3C0ECA98",
    x"3C0EB8C0",
    x"3C0EA6EA",
    x"3C0E9517",
    x"3C0E8345",
    x"3C0E7176",
    x"3C0E5FA9",
    x"3C0E4DDE",
    x"3C0E3C15",
    x"3C0E2A4F",
    x"3C0E188B",
    x"3C0E06C9",
    x"3C0DF509",
    x"3C0DE34B",
    x"3C0DD190",
    x"3C0DBFD7",
    x"3C0DAE20",
    x"3C0D9C6B",
    x"3C0D8AB9",
    x"3C0D7909",
    x"3C0D675B",
    x"3C0D55AF",
    x"3C0D4405",
    x"3C0D325E",
    x"3C0D20B9",
    x"3C0D0F16",
    x"3C0CFD75",
    x"3C0CEBD6",
    x"3C0CDA3A",
    x"3C0CC8A0",
    x"3C0CB708",
    x"3C0CA572",
    x"3C0C93DE",
    x"3C0C824D",
    x"3C0C70BE",
    x"3C0C5F31",
    x"3C0C4DA6",
    x"3C0C3C1E",
    x"3C0C2A97",
    x"3C0C1913",
    x"3C0C0791",
    x"3C0BF611",
    x"3C0BE493",
    x"3C0BD318",
    x"3C0BC19F",
    x"3C0BB027",
    x"3C0B9EB2",
    x"3C0B8D40",
    x"3C0B7BCF",
    x"3C0B6A61",
    x"3C0B58F5",
    x"3C0B478B",
    x"3C0B3623",
    x"3C0B24BD",
    x"3C0B135A",
    x"3C0B01F8",
    x"3C0AF099",
    x"3C0ADF3C",
    x"3C0ACDE1",
    x"3C0ABC89",
    x"3C0AAB32",
    x"3C0A99DE",
    x"3C0A888C",
    x"3C0A773C",
    x"3C0A65EE",
    x"3C0A54A2",
    x"3C0A4359",
    x"3C0A3211",
    x"3C0A20CC",
    x"3C0A0F89",
    x"3C09FE48",
    x"3C09ED0A",
    x"3C09DBCD",
    x"3C09CA93",
    x"3C09B95A",
    x"3C09A824",
    x"3C0996F0",
    x"3C0985BF",
    x"3C09748F",
    x"3C096361",
    x"3C095236",
    x"3C09410D",
    x"3C092FE6",
    x"3C091EC1",
    x"3C090D9E",
    x"3C08FC7D",
    x"3C08EB5F",
    x"3C08DA43",
    x"3C08C928",
    x"3C08B810",
    x"3C08A6FA",
    x"3C0895E7",
    x"3C0884D5",
    x"3C0873C5",
    x"3C0862B8",
    x"3C0851AD",
    x"3C0840A4",
    x"3C082F9D",
    x"3C081E98",
    x"3C080D95",
    x"3C07FC94",
    x"3C07EB96",
    x"3C07DA99",
    x"3C07C99F",
    x"3C07B8A7",
    x"3C07A7B1",
    x"3C0796BD",
    x"3C0785CB",
    x"3C0774DC",
    x"3C0763EE",
    x"3C075303",
    x"3C074219",
    x"3C073132",
    x"3C07204D",
    x"3C070F6A",
    x"3C06FE89",
    x"3C06EDAA",
    x"3C06DCCE",
    x"3C06CBF3",
    x"3C06BB1B",
    x"3C06AA44",
    x"3C069970",
    x"3C06889E",
    x"3C0677CE",
    x"3C066700",
    x"3C065634",
    x"3C06456A",
    x"3C0634A3",
    x"3C0623DD",
    x"3C06131A",
    x"3C060259",
    x"3C05F199",
    x"3C05E0DC",
    x"3C05D021",
    x"3C05BF68",
    x"3C05AEB1",
    x"3C059DFC",
    x"3C058D4A",
    x"3C057C99",
    x"3C056BEB",
    x"3C055B3E",
    x"3C054A94",
    x"3C0539EC",
    x"3C052945",
    x"3C0518A1",
    x"3C0507FF",
    x"3C04F75F",
    x"3C04E6C1",
    x"3C04D625",
    x"3C04C58C",
    x"3C04B4F4",
    x"3C04A45F",
    x"3C0493CB",
    x"3C04833A",
    x"3C0472AA",
    x"3C04621D",
    x"3C045192",
    x"3C044109",
    x"3C043081",
    x"3C041FFC",
    x"3C040F79",
    x"3C03FEF9",
    x"3C03EE7A",
    x"3C03DDFD",
    x"3C03CD82",
    x"3C03BD0A",
    x"3C03AC93",
    x"3C039C1E",
    x"3C038BAC",
    x"3C037B3B",
    x"3C036ACD",
    x"3C035A61",
    x"3C0349F6",
    x"3C03398E",
    x"3C032928",
    x"3C0318C4",
    x"3C030862",
    x"3C02F802",
    x"3C02E7A4",
    x"3C02D748",
    x"3C02C6EE",
    x"3C02B696",
    x"3C02A640",
    x"3C0295ED",
    x"3C02859B",
    x"3C02754B",
    x"3C0264FE",
    x"3C0254B2",
    x"3C024468",
    x"3C023421",
    x"3C0223DB",
    x"3C021398",
    x"3C020357",
    x"3C01F317",
    x"3C01E2DA",
    x"3C01D29E",
    x"3C01C265",
    x"3C01B22E",
    x"3C01A1F9",
    x"3C0191C5",
    x"3C018194",
    x"3C017165",
    x"3C016138",
    x"3C01510D",
    x"3C0140E4",
    x"3C0130BC",
    x"3C012097",
    x"3C011074",
    x"3C010053",
    x"3C00F034",
    x"3C00E017",
    x"3C00CFFC",
    x"3C00BFE3",
    x"3C00AFCC",
    x"3C009FB7",
    x"3C008FA4",
    x"3C007F93",
    x"3C006F84",
    x"3C005F77",
    x"3C004F6C",
    x"3C003F64",
    x"3C002F5D",
    x"3C001F58",
    x"3C000F55",
    x"3BFFFEA8",
    x"3BFFDEAA",
    x"3BFFBEB0",
    x"3BFF9EBA",
    x"3BFF7EC8",
    x"3BFF5EDB",
    x"3BFF3EF1",
    x"3BFF1F0B",
    x"3BFEFF29",
    x"3BFEDF4B",
    x"3BFEBF71",
    x"3BFE9F9B",
    x"3BFE7FC9",
    x"3BFE5FFB",
    x"3BFE4031",
    x"3BFE206B",
    x"3BFE00A9",
    x"3BFDE0EB",
    x"3BFDC131",
    x"3BFDA17B",
    x"3BFD81C9",
    x"3BFD621A",
    x"3BFD4270",
    x"3BFD22CA",
    x"3BFD0327",
    x"3BFCE389",
    x"3BFCC3EE",
    x"3BFCA458",
    x"3BFC84C5",
    x"3BFC6537",
    x"3BFC45AC",
    x"3BFC2625",
    x"3BFC06A2",
    x"3BFBE724",
    x"3BFBC7A9",
    x"3BFBA832",
    x"3BFB88BF",
    x"3BFB6950",
    x"3BFB49E4",
    x"3BFB2A7D",
    x"3BFB0B1A",
    x"3BFAEBBA",
    x"3BFACC5F",
    x"3BFAAD07",
    x"3BFA8DB4",
    x"3BFA6E64",
    x"3BFA4F18",
    x"3BFA2FD0",
    x"3BFA108C",
    x"3BF9F14C",
    x"3BF9D210",
    x"3BF9B2D7",
    x"3BF993A3",
    x"3BF97472",
    x"3BF95546",
    x"3BF9361D",
    x"3BF916F8",
    x"3BF8F7D7",
    x"3BF8D8BA",
    x"3BF8B9A1",
    x"3BF89A8C",
    x"3BF87B7B",
    x"3BF85C6D",
    x"3BF83D63",
    x"3BF81E5E",
    x"3BF7FF5C",
    x"3BF7E05E",
    x"3BF7C164",
    x"3BF7A26E",
    x"3BF7837B",
    x"3BF7648D",
    x"3BF745A2",
    x"3BF726BB",
    x"3BF707D8",
    x"3BF6E8F9",
    x"3BF6CA1E",
    x"3BF6AB47",
    x"3BF68C73",
    x"3BF66DA4",
    x"3BF64ED8",
    x"3BF63010",
    x"3BF6114C",
    x"3BF5F28C",
    x"3BF5D3CF",
    x"3BF5B517",
    x"3BF59662",
    x"3BF577B1",
    x"3BF55904",
    x"3BF53A5B",
    x"3BF51BB5",
    x"3BF4FD14",
    x"3BF4DE76",
    x"3BF4BFDC",
    x"3BF4A146",
    x"3BF482B4",
    x"3BF46425",
    x"3BF4459B",
    x"3BF42714",
    x"3BF40891",
    x"3BF3EA12",
    x"3BF3CB97",
    x"3BF3AD1F",
    x"3BF38EAB",
    x"3BF3703B",
    x"3BF351CF",
    x"3BF33367",
    x"3BF31502",
    x"3BF2F6A2",
    x"3BF2D845",
    x"3BF2B9EC",
    x"3BF29B96",
    x"3BF27D45",
    x"3BF25EF7",
    x"3BF240AD",
    x"3BF22267",
    x"3BF20424",
    x"3BF1E5E6",
    x"3BF1C7AB",
    x"3BF1A974",
    x"3BF18B41",
    x"3BF16D11",
    x"3BF14EE5",
    x"3BF130BD",
    x"3BF11299",
    x"3BF0F479",
    x"3BF0D65C",
    x"3BF0B843",
    x"3BF09A2E",
    x"3BF07C1D",
    x"3BF05E0F",
    x"3BF04005",
    x"3BF021FF",
    x"3BF003FC",
    x"3BEFE5FE",
    x"3BEFC803",
    x"3BEFAA0C",
    x"3BEF8C18",
    x"3BEF6E29",
    x"3BEF503D",
    x"3BEF3255",
    x"3BEF1470",
    x"3BEEF690",
    x"3BEED8B3",
    x"3BEEBAD9",
    x"3BEE9D04",
    x"3BEE7F32",
    x"3BEE6164",
    x"3BEE439A",
    x"3BEE25D3",
    x"3BEE0810",
    x"3BEDEA51",
    x"3BEDCC96",
    x"3BEDAEDE",
    x"3BED912A",
    x"3BED737A",
    x"3BED55CD",
    x"3BED3824",
    x"3BED1A7F",
    x"3BECFCDE",
    x"3BECDF40",
    x"3BECC1A6",
    x"3BECA410",
    x"3BEC867D",
    x"3BEC68EE",
    x"3BEC4B63",
    x"3BEC2DDB",
    x"3BEC1057",
    x"3BEBF2D7",
    x"3BEBD55B",
    x"3BEBB7E2",
    x"3BEB9A6D",
    x"3BEB7CFB",
    x"3BEB5F8D",
    x"3BEB4223",
    x"3BEB24BD",
    x"3BEB075A",
    x"3BEAE9FB",
    x"3BEACCA0",
    x"3BEAAF48",
    x"3BEA91F4",
    x"3BEA74A3",
    x"3BEA5757",
    x"3BEA3A0D",
    x"3BEA1CC8",
    x"3BE9FF86",
    x"3BE9E248",
    x"3BE9C50E",
    x"3BE9A7D7",
    x"3BE98AA4",
    x"3BE96D74",
    x"3BE95048",
    x"3BE93320",
    x"3BE915FC",
    x"3BE8F8DB",
    x"3BE8DBBD",
    x"3BE8BEA4",
    x"3BE8A18E",
    x"3BE8847B",
    x"3BE8676D",
    x"3BE84A61",
    x"3BE82D5A",
    x"3BE81056",
    x"3BE7F356",
    x"3BE7D659",
    x"3BE7B960",
    x"3BE79C6B",
    x"3BE77F79",
    x"3BE7628B",
    x"3BE745A1",
    x"3BE728BA",
    x"3BE70BD6",
    x"3BE6EEF7",
    x"3BE6D21B",
    x"3BE6B542",
    x"3BE6986D",
    x"3BE67B9C",
    x"3BE65ECE",
    x"3BE64204",
    x"3BE6253E",
    x"3BE6087B",
    x"3BE5EBBC",
    x"3BE5CF00",
    x"3BE5B248",
    x"3BE59594",
    x"3BE578E3",
    x"3BE55C35",
    x"3BE53F8C",
    x"3BE522E5",
    x"3BE50643",
    x"3BE4E9A4",
    x"3BE4CD08",
    x"3BE4B071",
    x"3BE493DC",
    x"3BE4774C",
    x"3BE45ABF",
    x"3BE43E35",
    x"3BE421AF",
    x"3BE4052D",
    x"3BE3E8AE",
    x"3BE3CC32",
    x"3BE3AFBB",
    x"3BE39346",
    x"3BE376D6",
    x"3BE35A69",
    x"3BE33DFF",
    x"3BE32199",
    x"3BE30537",
    x"3BE2E8D8",
    x"3BE2CC7D",
    x"3BE2B025",
    x"3BE293D1",
    x"3BE27780",
    x"3BE25B33",
    x"3BE23EE9",
    x"3BE222A3",
    x"3BE20660",
    x"3BE1EA21",
    x"3BE1CDE6",
    x"3BE1B1AE",
    x"3BE19579",
    x"3BE17949",
    x"3BE15D1B",
    x"3BE140F1",
    x"3BE124CB",
    x"3BE108A8",
    x"3BE0EC89",
    x"3BE0D06D",
    x"3BE0B455",
    x"3BE09840",
    x"3BE07C2F",
    x"3BE06021",
    x"3BE04417",
    x"3BE02810",
    x"3BE00C0D",
    x"3BDFF00D",
    x"3BDFD411",
    x"3BDFB818",
    x"3BDF9C22",
    x"3BDF8031",
    x"3BDF6442",
    x"3BDF4858",
    x"3BDF2C70",
    x"3BDF108D",
    x"3BDEF4AC",
    x"3BDED8CF",
    x"3BDEBCF6",
    x"3BDEA120",
    x"3BDE854E",
    x"3BDE697F",
    x"3BDE4DB3",
    x"3BDE31EB",
    x"3BDE1627",
    x"3BDDFA66",
    x"3BDDDEA8",
    x"3BDDC2EE",
    x"3BDDA738",
    x"3BDD8B84",
    x"3BDD6FD5",
    x"3BDD5428",
    x"3BDD3880",
    x"3BDD1CDA",
    x"3BDD0138",
    x"3BDCE59A",
    x"3BDCC9FF",
    x"3BDCAE67",
    x"3BDC92D3",
    x"3BDC7743",
    x"3BDC5BB6",
    x"3BDC402C",
    x"3BDC24A6",
    x"3BDC0923",
    x"3BDBEDA3",
    x"3BDBD227",
    x"3BDBB6AF",
    x"3BDB9B3A",
    x"3BDB7FC8",
    x"3BDB645A",
    x"3BDB48EF",
    x"3BDB2D87",
    x"3BDB1223",
    x"3BDAF6C3",
    x"3BDADB66",
    x"3BDAC00C",
    x"3BDAA4B6",
    x"3BDA8963",
    x"3BDA6E13",
    x"3BDA52C7",
    x"3BDA377F",
    x"3BDA1C39",
    x"3BDA00F8",
    x"3BD9E5B9",
    x"3BD9CA7E",
    x"3BD9AF47",
    x"3BD99412",
    x"3BD978E2",
    x"3BD95DB4",
    x"3BD9428A",
    x"3BD92764",
    x"3BD90C40",
    x"3BD8F120",
    x"3BD8D604",
    x"3BD8BAEB",
    x"3BD89FD5",
    x"3BD884C3",
    x"3BD869B4",
    x"3BD84EA9",
    x"3BD833A0",
    x"3BD8189C",
    x"3BD7FD9A",
    x"3BD7E29C",
    x"3BD7C7A2",
    x"3BD7ACAA",
    x"3BD791B6",
    x"3BD776C6",
    x"3BD75BD9",
    x"3BD740EF",
    x"3BD72609",
    x"3BD70B25",
    x"3BD6F046",
    x"3BD6D569",
    x"3BD6BA90",
    x"3BD69FBB",
    x"3BD684E8",
    x"3BD66A1A",
    x"3BD64F4E",
    x"3BD63486",
    x"3BD619C1",
    x"3BD5FEFF",
    x"3BD5E441",
    x"3BD5C986",
    x"3BD5AECF",
    x"3BD5941A",
    x"3BD5796A",
    x"3BD55EBC",
    x"3BD54412",
    x"3BD5296B",
    x"3BD50EC8",
    x"3BD4F427",
    x"3BD4D98B",
    x"3BD4BEF1",
    x"3BD4A45B",
    x"3BD489C8",
    x"3BD46F38",
    x"3BD454AC",
    x"3BD43A23",
    x"3BD41F9E",
    x"3BD4051B",
    x"3BD3EA9C",
    x"3BD3D021",
    x"3BD3B5A8",
    x"3BD39B33",
    x"3BD380C1",
    x"3BD36653",
    x"3BD34BE8",
    x"3BD33180",
    x"3BD3171C",
    x"3BD2FCBA",
    x"3BD2E25C",
    x"3BD2C802",
    x"3BD2ADAA",
    x"3BD29356",
    x"3BD27906",
    x"3BD25EB8",
    x"3BD2446E",
    x"3BD22A27",
    x"3BD20FE3",
    x"3BD1F5A3",
    x"3BD1DB66",
    x"3BD1C12C",
    x"3BD1A6F6",
    x"3BD18CC2",
    x"3BD17292",
    x"3BD15866",
    x"3BD13E3C",
    x"3BD12416",
    x"3BD109F3",
    x"3BD0EFD4",
    x"3BD0D5B7",
    x"3BD0BB9E",
    x"3BD0A188",
    x"3BD08776",
    x"3BD06D67",
    x"3BD0535B",
    x"3BD03952",
    x"3BD01F4C",
    x"3BD0054A",
    x"3BCFEB4B",
    x"3BCFD14F",
    x"3BCFB757",
    x"3BCF9D61",
    x"3BCF836F",
    x"3BCF6980",
    x"3BCF4F95",
    x"3BCF35AC",
    x"3BCF1BC7",
    x"3BCF01E6",
    x"3BCEE807",
    x"3BCECE2C",
    x"3BCEB453",
    x"3BCE9A7E",
    x"3BCE80AD",
    x"3BCE66DE",
    x"3BCE4D13",
    x"3BCE334B",
    x"3BCE1986",
    x"3BCDFFC5",
    x"3BCDE606",
    x"3BCDCC4B",
    x"3BCDB293",
    x"3BCD98DE",
    x"3BCD7F2D",
    x"3BCD657F",
    x"3BCD4BD4",
    x"3BCD322C",
    x"3BCD1887",
    x"3BCCFEE6",
    x"3BCCE547",
    x"3BCCCBAC",
    x"3BCCB214",
    x"3BCC9880",
    x"3BCC7EEE",
    x"3BCC6560",
    x"3BCC4BD5",
    x"3BCC324D",
    x"3BCC18C8",
    x"3BCBFF47",
    x"3BCBE5C9",
    x"3BCBCC4D",
    x"3BCBB2D5",
    x"3BCB9961",
    x"3BCB7FEF",
    x"3BCB6681",
    x"3BCB4D15",
    x"3BCB33AD",
    x"3BCB1A49",
    x"3BCB00E7",
    x"3BCAE788",
    x"3BCACE2D",
    x"3BCAB4D5",
    x"3BCA9B80",
    x"3BCA822E",
    x"3BCA68DF",
    x"3BCA4F94",
    x"3BCA364B",
    x"3BCA1D06",
    x"3BCA03C4",
    x"3BC9EA85",
    x"3BC9D149",
    x"3BC9B811",
    x"3BC99EDB",
    x"3BC985A9",
    x"3BC96C7A",
    x"3BC9534E",
    x"3BC93A25",
    x"3BC92100",
    x"3BC907DD",
    x"3BC8EEBE",
    x"3BC8D5A1",
    x"3BC8BC88",
    x"3BC8A372",
    x"3BC88A5F",
    x"3BC87150",
    x"3BC85843",
    x"3BC83F39",
    x"3BC82633",
    x"3BC80D30",
    x"3BC7F430",
    x"3BC7DB33",
    x"3BC7C239",
    x"3BC7A942",
    x"3BC7904F",
    x"3BC7775E",
    x"3BC75E71",
    x"3BC74587",
    x"3BC72C9F",
    x"3BC713BB",
    x"3BC6FADB",
    x"3BC6E1FD",
    x"3BC6C922",
    x"3BC6B04A",
    x"3BC69776",
    x"3BC67EA5",
    x"3BC665D6",
    x"3BC64D0B",
    x"3BC63443",
    x"3BC61B7E",
    x"3BC602BC",
    x"3BC5E9FD",
    x"3BC5D142",
    x"3BC5B889",
    x"3BC59FD4",
    x"3BC58721",
    x"3BC56E72",
    x"3BC555C6",
    x"3BC53D1C",
    x"3BC52476",
    x"3BC50BD3",
    x"3BC4F333",
    x"3BC4DA96",
    x"3BC4C1FD",
    x"3BC4A966",
    x"3BC490D2",
    x"3BC47842",
    x"3BC45FB4",
    x"3BC4472A",
    x"3BC42EA2",
    x"3BC4161E",
    x"3BC3FD9D",
    x"3BC3E51F",
    x"3BC3CCA4",
    x"3BC3B42C",
    x"3BC39BB7",
    x"3BC38345",
    x"3BC36AD6",
    x"3BC3526A",
    x"3BC33A01",
    x"3BC3219B",
    x"3BC30939",
    x"3BC2F0D9",
    x"3BC2D87D",
    x"3BC2C023",
    x"3BC2A7CD",
    x"3BC28F79",
    x"3BC27729",
    x"3BC25EDB",
    x"3BC24691",
    x"3BC22E4A",
    x"3BC21605",
    x"3BC1FDC4",
    x"3BC1E586",
    x"3BC1CD4B",
    x"3BC1B513",
    x"3BC19CDD",
    x"3BC184AB",
    x"3BC16C7C",
    x"3BC15450",
    x"3BC13C27",
    x"3BC12401",
    x"3BC10BDE",
    x"3BC0F3BE",
    x"3BC0DBA1",
    x"3BC0C387",
    x"3BC0AB70",
    x"3BC0935C",
    x"3BC07B4C",
    x"3BC0633E",
    x"3BC04B33",
    x"3BC0332B",
    x"3BC01B26",
    x"3BC00324",
    x"3BBFEB25",
    x"3BBFD329",
    x"3BBFBB30",
    x"3BBFA33A",
    x"3BBF8B48",
    x"3BBF7358",
    x"3BBF5B6B",
    x"3BBF4381",
    x"3BBF2B9A",
    x"3BBF13B6",
    x"3BBEFBD5",
    x"3BBEE3F7",
    x"3BBECC1C",
    x"3BBEB444",
    x"3BBE9C6F",
    x"3BBE849D",
    x"3BBE6CCE",
    x"3BBE5502",
    x"3BBE3D38",
    x"3BBE2572",
    x"3BBE0DAF",
    x"3BBDF5EF",
    x"3BBDDE32",
    x"3BBDC677",
    x"3BBDAEC0",
    x"3BBD970C",
    x"3BBD7F5A",
    x"3BBD67AC",
    x"3BBD5000",
    x"3BBD3858",
    x"3BBD20B2",
    x"3BBD0910",
    x"3BBCF170",
    x"3BBCD9D3",
    x"3BBCC23A",
    x"3BBCAAA3",
    x"3BBC930F",
    x"3BBC7B7E",
    x"3BBC63F0",
    x"3BBC4C65",
    x"3BBC34DD",
    x"3BBC1D58",
    x"3BBC05D6",
    x"3BBBEE56",
    x"3BBBD6DA",
    x"3BBBBF61",
    x"3BBBA7EA",
    x"3BBB9077",
    x"3BBB7906",
    x"3BBB6198",
    x"3BBB4A2E",
    x"3BBB32C6",
    x"3BBB1B61",
    x"3BBB03FF",
    x"3BBAECA0",
    x"3BBAD544",
    x"3BBABDEB",
    x"3BBAA694",
    x"3BBA8F41",
    x"3BBA77F0",
    x"3BBA60A3",
    x"3BBA4958",
    x"3BBA3211",
    x"3BBA1ACC",
    x"3BBA038A",
    x"3BB9EC4B",
    x"3BB9D50F",
    x"3BB9BDD6",
    x"3BB9A69F",
    x"3BB98F6C",
    x"3BB9783C",
    x"3BB9610E",
    x"3BB949E3",
    x"3BB932BB",
    x"3BB91B97",
    x"3BB90475",
    x"3BB8ED55",
    x"3BB8D639",
    x"3BB8BF20",
    x"3BB8A809",
    x"3BB890F6",
    x"3BB879E5",
    x"3BB862D7",
    x"3BB84BCD",
    x"3BB834C4",
    x"3BB81DBF",
    x"3BB806BD",
    x"3BB7EFBE",
    x"3BB7D8C1",
    x"3BB7C1C7",
    x"3BB7AAD1",
    x"3BB793DD",
    x"3BB77CEC",
    x"3BB765FE",
    x"3BB74F12",
    x"3BB7382A",
    x"3BB72144",
    x"3BB70A61",
    x"3BB6F382",
    x"3BB6DCA5",
    x"3BB6C5CA",
    x"3BB6AEF3",
    x"3BB6981F",
    x"3BB6814D",
    x"3BB66A7E",
    x"3BB653B2",
    x"3BB63CE9",
    x"3BB62623",
    x"3BB60F60",
    x"3BB5F89F",
    x"3BB5E1E2",
    x"3BB5CB27",
    x"3BB5B46F",
    x"3BB59DBA",
    x"3BB58708",
    x"3BB57058",
    x"3BB559AB",
    x"3BB54302",
    x"3BB52C5B",
    x"3BB515B7",
    x"3BB4FF15",
    x"3BB4E877",
    x"3BB4D1DB",
    x"3BB4BB42",
    x"3BB4A4AC",
    x"3BB48E19",
    x"3BB47789",
    x"3BB460FB",
    x"3BB44A71",
    x"3BB433E9",
    x"3BB41D64",
    x"3BB406E1",
    x"3BB3F062",
    x"3BB3D9E5",
    x"3BB3C36B",
    x"3BB3ACF4",
    x"3BB39680",
    x"3BB3800F",
    x"3BB369A0",
    x"3BB35334",
    x"3BB33CCB",
    x"3BB32665",
    x"3BB31002",
    x"3BB2F9A1",
    x"3BB2E343",
    x"3BB2CCE8",
    x"3BB2B690",
    x"3BB2A03B",
    x"3BB289E8",
    x"3BB27398",
    x"3BB25D4B",
    x"3BB24701",
    x"3BB230B9",
    x"3BB21A75",
    x"3BB20433",
    x"3BB1EDF4",
    x"3BB1D7B7",
    x"3BB1C17E",
    x"3BB1AB47",
    x"3BB19513",
    x"3BB17EE2",
    x"3BB168B3",
    x"3BB15287",
    x"3BB13C5F",
    x"3BB12638",
    x"3BB11015",
    x"3BB0F9F4",
    x"3BB0E3D6",
    x"3BB0CDBB",
    x"3BB0B7A3",
    x"3BB0A18D",
    x"3BB08B7B",
    x"3BB0756B",
    x"3BB05F5D",
    x"3BB04953",
    x"3BB0334B",
    x"3BB01D46",
    x"3BB00744",
    x"3BAFF144",
    x"3BAFDB47",
    x"3BAFC54D",
    x"3BAFAF56",
    x"3BAF9961",
    x"3BAF8370",
    x"3BAF6D81",
    x"3BAF5794",
    x"3BAF41AB",
    x"3BAF2BC4",
    x"3BAF15E0",
    x"3BAEFFFE",
    x"3BAEEA20",
    x"3BAED444",
    x"3BAEBE6B",
    x"3BAEA894",
    x"3BAE92C1",
    x"3BAE7CF0",
    x"3BAE6721",
    x"3BAE5156",
    x"3BAE3B8D",
    x"3BAE25C7",
    x"3BAE1004",
    x"3BADFA43",
    x"3BADE485",
    x"3BADCECA",
    x"3BADB911",
    x"3BADA35B",
    x"3BAD8DA8",
    x"3BAD77F8",
    x"3BAD624A",
    x"3BAD4CA0",
    x"3BAD36F7",
    x"3BAD2152",
    x"3BAD0BAF",
    x"3BACF60F",
    x"3BACE071",
    x"3BACCAD7",
    x"3BACB53F",
    x"3BAC9FA9",
    x"3BAC8A17",
    x"3BAC7487",
    x"3BAC5EFA",
    x"3BAC496F",
    x"3BAC33E7",
    x"3BAC1E62",
    x"3BAC08E0",
    x"3BABF360",
    x"3BABDDE3",
    x"3BABC868",
    x"3BABB2F1",
    x"3BAB9D7C",
    x"3BAB8809",
    x"3BAB729A",
    x"3BAB5D2D",
    x"3BAB47C2",
    x"3BAB325B",
    x"3BAB1CF6",
    x"3BAB0794",
    x"3BAAF234",
    x"3BAADCD7",
    x"3BAAC77D",
    x"3BAAB225",
    x"3BAA9CD0",
    x"3BAA877E",
    x"3BAA722E",
    x"3BAA5CE1",
    x"3BAA4797",
    x"3BAA3250",
    x"3BAA1D0B",
    x"3BAA07C8",
    x"3BA9F289",
    x"3BA9DD4C",
    x"3BA9C811",
    x"3BA9B2DA",
    x"3BA99DA5",
    x"3BA98872",
    x"3BA97342",
    x"3BA95E15",
    x"3BA948EB",
    x"3BA933C3",
    x"3BA91E9E",
    x"3BA9097B",
    x"3BA8F45C",
    x"3BA8DF3E",
    x"3BA8CA24",
    x"3BA8B50C",
    x"3BA89FF7",
    x"3BA88AE4",
    x"3BA875D4",
    x"3BA860C6",
    x"3BA84BBC",
    x"3BA836B3",
    x"3BA821AE",
    x"3BA80CAB",
    x"3BA7F7AB",
    x"3BA7E2AD",
    x"3BA7CDB2",
    x"3BA7B8BA",
    x"3BA7A3C4",
    x"3BA78ED1",
    x"3BA779E0",
    x"3BA764F2",
    x"3BA75007",
    x"3BA73B1E",
    x"3BA72638",
    x"3BA71155",
    x"3BA6FC74",
    x"3BA6E796",
    x"3BA6D2BA",
    x"3BA6BDE1",
    x"3BA6A90B",
    x"3BA69437",
    x"3BA67F65",
    x"3BA66A97",
    x"3BA655CB",
    x"3BA64101",
    x"3BA62C3B",
    x"3BA61776",
    x"3BA602B5",
    x"3BA5EDF6",
    x"3BA5D939",
    x"3BA5C47F",
    x"3BA5AFC8",
    x"3BA59B13",
    x"3BA58661",
    x"3BA571B2",
    x"3BA55D05",
    x"3BA5485B",
    x"3BA533B3",
    x"3BA51F0E",
    x"3BA50A6B",
    x"3BA4F5CB",
    x"3BA4E12E",
    x"3BA4CC93",
    x"3BA4B7FA",
    x"3BA4A365",
    x"3BA48ED2",
    x"3BA47A41",
    x"3BA465B3",
    x"3BA45128",
    x"3BA43C9F",
    x"3BA42818",
    x"3BA41395",
    x"3BA3FF14",
    x"3BA3EA95",
    x"3BA3D619",
    x"3BA3C19F",
    x"3BA3AD28",
    x"3BA398B4",
    x"3BA38442",
    x"3BA36FD3",
    x"3BA35B66",
    x"3BA346FC",
    x"3BA33295",
    x"3BA31E30",
    x"3BA309CD",
    x"3BA2F56D",
    x"3BA2E110",
    x"3BA2CCB5",
    x"3BA2B85D",
    x"3BA2A407",
    x"3BA28FB4",
    x"3BA27B63",
    x"3BA26715",
    x"3BA252C9",
    x"3BA23E80",
    x"3BA22A39",
    x"3BA215F5",
    x"3BA201B4",
    x"3BA1ED75",
    x"3BA1D939",
    x"3BA1C4FF",
    x"3BA1B0C7",
    x"3BA19C92",
    x"3BA18860",
    x"3BA17430",
    x"3BA16003",
    x"3BA14BD8",
    x"3BA137B0",
    x"3BA1238A",
    x"3BA10F67",
    x"3BA0FB47",
    x"3BA0E728",
    x"3BA0D30D",
    x"3BA0BEF4",
    x"3BA0AADD",
    x"3BA096C9",
    x"3BA082B7",
    x"3BA06EA8",
    x"3BA05A9C",
    x"3BA04692",
    x"3BA0328A",
    x"3BA01E85",
    x"3BA00A82",
    x"3B9FF682",
    x"3B9FE285",
    x"3B9FCE8A",
    x"3B9FBA91",
    x"3B9FA69B",
    x"3B9F92A8",
    x"3B9F7EB6",
    x"3B9F6AC8",
    x"3B9F56DC",
    x"3B9F42F2",
    x"3B9F2F0B",
    x"3B9F1B26",
    x"3B9F0744",
    x"3B9EF365",
    x"3B9EDF87",
    x"3B9ECBAD",
    x"3B9EB7D4",
    x"3B9EA3FF",
    x"3B9E902B",
    x"3B9E7C5B",
    x"3B9E688C",
    x"3B9E54C1",
    x"3B9E40F7",
    x"3B9E2D30",
    x"3B9E196C",
    x"3B9E05AA",
    x"3B9DF1EA",
    x"3B9DDE2D",
    x"3B9DCA73",
    x"3B9DB6BB",
    x"3B9DA305",
    x"3B9D8F52",
    x"3B9D7BA1",
    x"3B9D67F3",
    x"3B9D5447",
    x"3B9D409E",
    x"3B9D2CF7",
    x"3B9D1953",
    x"3B9D05B1",
    x"3B9CF211",
    x"3B9CDE74",
    x"3B9CCADA",
    x"3B9CB742",
    x"3B9CA3AC",
    x"3B9C9019",
    x"3B9C7C88",
    x"3B9C68FA",
    x"3B9C556E",
    x"3B9C41E4",
    x"3B9C2E5D",
    x"3B9C1AD9",
    x"3B9C0757",
    x"3B9BF3D7",
    x"3B9BE05A",
    x"3B9BCCDF",
    x"3B9BB966",
    x"3B9BA5F0",
    x"3B9B927D",
    x"3B9B7F0C",
    x"3B9B6B9D",
    x"3B9B5831",
    x"3B9B44C7",
    x"3B9B3160",
    x"3B9B1DFB",
    x"3B9B0A98",
    x"3B9AF738",
    x"3B9AE3DA",
    x"3B9AD07F",
    x"3B9ABD26",
    x"3B9AA9D0",
    x"3B9A967C",
    x"3B9A832A",
    x"3B9A6FDB",
    x"3B9A5C8E",
    x"3B9A4944",
    x"3B9A35FC",
    x"3B9A22B6",
    x"3B9A0F73",
    x"3B99FC33",
    x"3B99E8F4",
    x"3B99D5B8",
    x"3B99C27F",
    x"3B99AF48",
    x"3B999C13",
    x"3B9988E1",
    x"3B9975B1",
    x"3B996283",
    x"3B994F58",
    x"3B993C2F",
    x"3B992909",
    x"3B9915E5",
    x"3B9902C4",
    x"3B98EFA4",
    x"3B98DC88",
    x"3B98C96D",
    x"3B98B655",
    x"3B98A340",
    x"3B98902D",
    x"3B987D1C",
    x"3B986A0D",
    x"3B985701",
    x"3B9843F8",
    x"3B9830F0",
    x"3B981DEB",
    x"3B980AE9",
    x"3B97F7E9",
    x"3B97E4EB",
    x"3B97D1EF",
    x"3B97BEF6",
    x"3B97AC00",
    x"3B97990B",
    x"3B978619",
    x"3B97732A",
    x"3B97603D",
    x"3B974D52",
    x"3B973A69",
    x"3B972783",
    x"3B97149F",
    x"3B9701BE",
    x"3B96EEDF",
    x"3B96DC02",
    x"3B96C928",
    x"3B96B650",
    x"3B96A37A",
    x"3B9690A7",
    x"3B967DD6",
    x"3B966B08",
    x"3B96583B",
    x"3B964572",
    x"3B9632AA",
    x"3B961FE5",
    x"3B960D22",
    x"3B95FA62",
    x"3B95E7A3",
    x"3B95D4E8",
    x"3B95C22E",
    x"3B95AF77",
    x"3B959CC2",
    x"3B958A10",
    x"3B957760",
    x"3B9564B2",
    x"3B955207",
    x"3B953F5E",
    x"3B952CB7",
    x"3B951A12",
    x"3B950770",
    x"3B94F4D1",
    x"3B94E233",
    x"3B94CF98",
    x"3B94BCFF",
    x"3B94AA69",
    x"3B9497D5",
    x"3B948543",
    x"3B9472B3",
    x"3B946026",
    x"3B944D9B",
    x"3B943B13",
    x"3B94288C",
    x"3B941609",
    x"3B940387",
    x"3B93F108",
    x"3B93DE8B",
    x"3B93CC10",
    x"3B93B998",
    x"3B93A722",
    x"3B9394AE",
    x"3B93823C",
    x"3B936FCD",
    x"3B935D61",
    x"3B934AF6",
    x"3B93388E",
    x"3B932628",
    x"3B9313C4",
    x"3B930163",
    x"3B92EF04",
    x"3B92DCA7",
    x"3B92CA4D",
    x"3B92B7F5",
    x"3B92A59F",
    x"3B92934B",
    x"3B9280FA",
    x"3B926EAB",
    x"3B925C5E",
    x"3B924A14",
    x"3B9237CC",
    x"3B922586",
    x"3B921342",
    x"3B920101",
    x"3B91EEC2",
    x"3B91DC85",
    x"3B91CA4B",
    x"3B91B813",
    x"3B91A5DD",
    x"3B9193A9",
    x"3B918178",
    x"3B916F49",
    x"3B915D1C",
    x"3B914AF2",
    x"3B9138C9",
    x"3B9126A4",
    x"3B911480",
    x"3B91025E",
    x"3B90F03F",
    x"3B90DE22",
    x"3B90CC08",
    x"3B90B9EF",
    x"3B90A7D9",
    x"3B9095C5",
    x"3B9083B4",
    x"3B9071A4",
    x"3B905F97",
    x"3B904D8D",
    x"3B903B84",
    x"3B90297E",
    x"3B90177A",
    x"3B900578",
    x"3B8FF378",
    x"3B8FE17B",
    x"3B8FCF80",
    x"3B8FBD87",
    x"3B8FAB90",
    x"3B8F999C",
    x"3B8F87AA",
    x"3B8F75BA",
    x"3B8F63CD",
    x"3B8F51E1",
    x"3B8F3FF8",
    x"3B8F2E11",
    x"3B8F1C2D",
    x"3B8F0A4A",
    x"3B8EF86A",
    x"3B8EE68C",
    x"3B8ED4B0",
    x"3B8EC2D7",
    x"3B8EB100",
    x"3B8E9F2B",
    x"3B8E8D58",
    x"3B8E7B87",
    x"3B8E69B9",
    x"3B8E57ED",
    x"3B8E4623",
    x"3B8E345B",
    x"3B8E2296",
    x"3B8E10D3",
    x"3B8DFF12",
    x"3B8DED53",
    x"3B8DDB96",
    x"3B8DC9DC",
    x"3B8DB824",
    x"3B8DA66E",
    x"3B8D94BA",
    x"3B8D8309",
    x"3B8D715A",
    x"3B8D5FAD",
    x"3B8D4E02",
    x"3B8D3C59",
    x"3B8D2AB3",
    x"3B8D190E",
    x"3B8D076C",
    x"3B8CF5CD",
    x"3B8CE42F",
    x"3B8CD293",
    x"3B8CC0FA",
    x"3B8CAF63",
    x"3B8C9DCE",
    x"3B8C8C3C",
    x"3B8C7AAB",
    x"3B8C691D",
    x"3B8C5791",
    x"3B8C4607",
    x"3B8C3480",
    x"3B8C22FA",
    x"3B8C1177",
    x"3B8BFFF6",
    x"3B8BEE77",
    x"3B8BDCFA",
    x"3B8BCB80",
    x"3B8BBA07",
    x"3B8BA891",
    x"3B8B971D",
    x"3B8B85AB",
    x"3B8B743C",
    x"3B8B62CE",
    x"3B8B5163",
    x"3B8B3FFA",
    x"3B8B2E93",
    x"3B8B1D2E",
    x"3B8B0BCC",
    x"3B8AFA6B",
    x"3B8AE90D",
    x"3B8AD7B1",
    x"3B8AC657",
    x"3B8AB4FF",
    x"3B8AA3AA",
    x"3B8A9257",
    x"3B8A8105",
    x"3B8A6FB6",
    x"3B8A5E69",
    x"3B8A4D1F",
    x"3B8A3BD6",
    x"3B8A2A90",
    x"3B8A194B",
    x"3B8A0809",
    x"3B89F6C9",
    x"3B89E58C",
    x"3B89D450",
    x"3B89C317",
    x"3B89B1DF",
    x"3B89A0AA",
    x"3B898F77",
    x"3B897E46",
    x"3B896D18",
    x"3B895BEB",
    x"3B894AC1",
    x"3B893998",
    x"3B892872",
    x"3B89174E",
    x"3B89062C",
    x"3B88F50D",
    x"3B88E3EF",
    x"3B88D2D4",
    x"3B88C1BA",
    x"3B88B0A3",
    x"3B889F8E",
    x"3B888E7B",
    x"3B887D6B",
    x"3B886C5C",
    x"3B885B50",
    x"3B884A45",
    x"3B88393D",
    x"3B882837",
    x"3B881733",
    x"3B880631",
    x"3B87F531",
    x"3B87E434",
    x"3B87D338",
    x"3B87C23F",
    x"3B87B148",
    x"3B87A053",
    x"3B878F60",
    x"3B877E6F",
    x"3B876D80",
    x"3B875C93",
    x"3B874BA9",
    x"3B873AC0",
    x"3B8729DA",
    x"3B8718F6",
    x"3B870814",
    x"3B86F734",
    x"3B86E656",
    x"3B86D57A",
    x"3B86C4A1",
    x"3B86B3C9",
    x"3B86A2F4",
    x"3B869221",
    x"3B86814F",
    x"3B867080",
    x"3B865FB3",
    x"3B864EE8",
    x"3B863E1F",
    x"3B862D59",
    x"3B861C94",
    x"3B860BD2",
    x"3B85FB11",
    x"3B85EA53",
    x"3B85D997",
    x"3B85C8DC",
    x"3B85B824",
    x"3B85A76E",
    x"3B8596BB",
    x"3B858609",
    x"3B857559",
    x"3B8564AB",
    x"3B855400",
    x"3B854356",
    x"3B8532AF",
    x"3B85220A",
    x"3B851166",
    x"3B8500C5",
    x"3B84F026",
    x"3B84DF89",
    x"3B84CEEE",
    x"3B84BE56",
    x"3B84ADBF",
    x"3B849D2A",
    x"3B848C98",
    x"3B847C07",
    x"3B846B79",
    x"3B845AEC",
    x"3B844A62",
    x"3B8439DA",
    x"3B842953",
    x"3B8418CF",
    x"3B84084D",
    x"3B83F7CD",
    x"3B83E74F",
    x"3B83D6D3",
    x"3B83C659",
    x"3B83B5E2",
    x"3B83A56C",
    x"3B8394F8",
    x"3B838487",
    x"3B837417",
    x"3B8363AA",
    x"3B83533E",
    x"3B8342D5",
    x"3B83326E",
    x"3B832208",
    x"3B8311A5",
    x"3B830144",
    x"3B82F0E5",
    x"3B82E088",
    x"3B82D02D",
    x"3B82BFD4",
    x"3B82AF7D",
    x"3B829F28",
    x"3B828ED5",
    x"3B827E84",
    x"3B826E35",
    x"3B825DE9",
    x"3B824D9E",
    x"3B823D55",
    x"3B822D0E",
    x"3B821CCA",
    x"3B820C87",
    x"3B81FC47",
    x"3B81EC08",
    x"3B81DBCC",
    x"3B81CB91",
    x"3B81BB59",
    x"3B81AB22",
    x"3B819AEE",
    x"3B818ABC",
    x"3B817A8B",
    x"3B816A5D",
    x"3B815A31",
    x"3B814A06",
    x"3B8139DE",
    x"3B8129B8",
    x"3B811994",
    x"3B810972",
    x"3B80F951",
    x"3B80E933",
    x"3B80D917",
    x"3B80C8FD",
    x"3B80B8E5",
    x"3B80A8CF",
    x"3B8098BB",
    x"3B8088A9",
    x"3B807899",
    x"3B80688A",
    x"3B80587E",
    x"3B804874",
    x"3B80386C",
    x"3B802866",
    x"3B801862",
    x"3B800860",
    x"3B7FF0C0",
    x"3B7FD0C4",
    x"3B7FB0CC",
    x"3B7F90D8",
    x"3B7F70E8",
    x"3B7F50FC",
    x"3B7F3114",
    x"3B7F112F",
    x"3B7EF14F",
    x"3B7ED173",
    x"3B7EB19B",
    x"3B7E91C7",
    x"3B7E71F6",
    x"3B7E522A",
    x"3B7E3262",
    x"3B7E129E",
    x"3B7DF2DD",
    x"3B7DD321",
    x"3B7DB368",
    x"3B7D93B4",
    x"3B7D7404",
    x"3B7D5457",
    x"3B7D34AE",
    x"3B7D150A",
    x"3B7CF569",
    x"3B7CD5CC",
    x"3B7CB634",
    x"3B7C969F",
    x"3B7C770E",
    x"3B7C5781",
    x"3B7C37F8",
    x"3B7C1873",
    x"3B7BF8F2",
    x"3B7BD975",
    x"3B7BB9FC",
    x"3B7B9A86",
    x"3B7B7B15",
    x"3B7B5BA8",
    x"3B7B3C3E",
    x"3B7B1CD9",
    x"3B7AFD77",
    x"3B7ADE19",
    x"3B7ABEBF",
    x"3B7A9F6A",
    x"3B7A8018",
    x"3B7A60CA",
    x"3B7A417F",
    x"3B7A2239",
    x"3B7A02F7",
    x"3B79E3B8",
    x"3B79C47E",
    x"3B79A547",
    x"3B798615",
    x"3B7966E6",
    x"3B7947BB",
    x"3B792894",
    x"3B790971",
    x"3B78EA51",
    x"3B78CB36",
    x"3B78AC1F",
    x"3B788D0B",
    x"3B786DFB",
    x"3B784EF0",
    x"3B782FE8",
    x"3B7810E4",
    x"3B77F1E3",
    x"3B77D2E7",
    x"3B77B3EF",
    x"3B7794FA",
    x"3B777609",
    x"3B77571D",
    x"3B773834",
    x"3B77194F",
    x"3B76FA6D",
    x"3B76DB90",
    x"3B76BCB6",
    x"3B769DE1",
    x"3B767F0F",
    x"3B766041",
    x"3B764177",
    x"3B7622B1",
    x"3B7603EE",
    x"3B75E530",
    x"3B75C675",
    x"3B75A7BE",
    x"3B75890B",
    x"3B756A5C",
    x"3B754BB0",
    x"3B752D09",
    x"3B750E65",
    x"3B74EFC5",
    x"3B74D129",
    x"3B74B291",
    x"3B7493FD",
    x"3B74756C",
    x"3B7456DF",
    x"3B743856",
    x"3B7419D1",
    x"3B73FB50",
    x"3B73DCD2",
    x"3B73BE59",
    x"3B739FE3",
    x"3B738171",
    x"3B736302",
    x"3B734498",
    x"3B732631",
    x"3B7307CE",
    x"3B72E96F",
    x"3B72CB14",
    x"3B72ACBD",
    x"3B728E69",
    x"3B727019",
    x"3B7251CD",
    x"3B723384",
    x"3B721540",
    x"3B71F6FF",
    x"3B71D8C2",
    x"3B71BA89",
    x"3B719C54",
    x"3B717E22",
    x"3B715FF4",
    x"3B7141CA",
    x"3B7123A4",
    x"3B710581",
    x"3B70E762",
    x"3B70C947",
    x"3B70AB30",
    x"3B708D1C",
    x"3B706F0D",
    x"3B705101",
    x"3B7032F8",
    x"3B7014F4",
    x"3B6FF6F3",
    x"3B6FD8F6",
    x"3B6FBAFD",
    x"3B6F9D07",
    x"3B6F7F16",
    x"3B6F6128",
    x"3B6F433D",
    x"3B6F2557",
    x"3B6F0774",
    x"3B6EE995",
    x"3B6ECBBA",
    x"3B6EADE2",
    x"3B6E900E",
    x"3B6E723E",
    x"3B6E5472",
    x"3B6E36A9",
    x"3B6E18E4",
    x"3B6DFB23",
    x"3B6DDD65",
    x"3B6DBFAB",
    x"3B6DA1F5",
    x"3B6D8443",
    x"3B6D6694",
    x"3B6D48E9",
    x"3B6D2B42",
    x"3B6D0D9E",
    x"3B6CEFFE",
    x"3B6CD262",
    x"3B6CB4CA",
    x"3B6C9735",
    x"3B6C79A4",
    x"3B6C5C17",
    x"3B6C3E8D",
    x"3B6C2107",
    x"3B6C0385",
    x"3B6BE606",
    x"3B6BC88B",
    x"3B6BAB14",
    x"3B6B8DA1",
    x"3B6B7031",
    x"3B6B52C4",
    x"3B6B355C",
    x"3B6B17F7",
    x"3B6AFA96",
    x"3B6ADD38",
    x"3B6ABFDF",
    x"3B6AA289",
    x"3B6A8536",
    x"3B6A67E7",
    x"3B6A4A9C",
    x"3B6A2D55",
    x"3B6A1011",
    x"3B69F2D1",
    x"3B69D594",
    x"3B69B85B",
    x"3B699B26",
    x"3B697DF4",
    x"3B6960C6",
    x"3B69439C",
    x"3B692676",
    x"3B690953",
    x"3B68EC33",
    x"3B68CF18",
    x"3B68B1FF",
    x"3B6894EB",
    x"3B6877DA",
    x"3B685ACD",
    x"3B683DC4",
    x"3B6820BE",
    x"3B6803BB",
    x"3B67E6BD",
    x"3B67C9C2",
    x"3B67ACCA",
    x"3B678FD6",
    x"3B6772E6",
    x"3B6755FA",
    x"3B673911",
    x"3B671C2B",
    x"3B66FF4A",
    x"3B66E26C",
    x"3B66C591",
    x"3B66A8BA",
    x"3B668BE7",
    x"3B666F17",
    x"3B66524B",
    x"3B663583",
    x"3B6618BE",
    x"3B65FBFC",
    x"3B65DF3F",
    x"3B65C285",
    x"3B65A5CE",
    x"3B65891B",
    x"3B656C6C",
    x"3B654FC0",
    x"3B653318",
    x"3B651673",
    x"3B64F9D2",
    x"3B64DD35",
    x"3B64C09B",
    x"3B64A405",
    x"3B648772",
    x"3B646AE3",
    x"3B644E57",
    x"3B6431CF",
    x"3B64154B",
    x"3B63F8CA",
    x"3B63DC4D",
    x"3B63BFD3",
    x"3B63A35D",
    x"3B6386EA",
    x"3B636A7B",
    x"3B634E0F",
    x"3B6331A7",
    x"3B631543",
    x"3B62F8E2",
    x"3B62DC85",
    x"3B62C02B",
    x"3B62A3D5",
    x"3B628782",
    x"3B626B33",
    x"3B624EE7",
    x"3B62329F",
    x"3B62165B",
    x"3B61FA1A",
    x"3B61DDDC",
    x"3B61C1A2",
    x"3B61A56C",
    x"3B618939",
    x"3B616D09",
    x"3B6150DD",
    x"3B6134B5",
    x"3B611890",
    x"3B60FC6F",
    x"3B60E051",
    x"3B60C437",
    x"3B60A820",
    x"3B608C0D",
    x"3B606FFD",
    x"3B6053F1",
    x"3B6037E8",
    x"3B601BE3",
    x"3B5FFFE1",
    x"3B5FE3E3",
    x"3B5FC7E8",
    x"3B5FABF1",
    x"3B5F8FFD",
    x"3B5F740D",
    x"3B5F5820",
    x"3B5F3C37",
    x"3B5F2051",
    x"3B5F046F",
    x"3B5EE890",
    x"3B5ECCB5",
    x"3B5EB0DD",
    x"3B5E9508",
    x"3B5E7938",
    x"3B5E5D6A",
    x"3B5E41A0",
    x"3B5E25DA",
    x"3B5E0A17",
    x"3B5DEE57",
    x"3B5DD29B",
    x"3B5DB6E3",
    x"3B5D9B2D",
    x"3B5D7F7C",
    x"3B5D63CE",
    x"3B5D4823",
    x"3B5D2C7C",
    x"3B5D10D8",
    x"3B5CF537",
    x"3B5CD99A",
    x"3B5CBE01",
    x"3B5CA26B",
    x"3B5C86D8",
    x"3B5C6B49",
    x"3B5C4FBE",
    x"3B5C3435",
    x"3B5C18B0",
    x"3B5BFD2F",
    x"3B5BE1B1",
    x"3B5BC637",
    x"3B5BAAC0",
    x"3B5B8F4C",
    x"3B5B73DC",
    x"3B5B586F",
    x"3B5B3D06",
    x"3B5B21A0",
    x"3B5B063D",
    x"3B5AEADE",
    x"3B5ACF83",
    x"3B5AB42A",
    x"3B5A98D6",
    x"3B5A7D84",
    x"3B5A6236",
    x"3B5A46EC",
    x"3B5A2BA4",
    x"3B5A1061",
    x"3B59F520",
    x"3B59D9E3",
    x"3B59BEAA",
    x"3B59A374",
    x"3B598841",
    x"3B596D12",
    x"3B5951E6",
    x"3B5936BD",
    x"3B591B98",
    x"3B590076",
    x"3B58E558",
    x"3B58CA3D",
    x"3B58AF25",
    x"3B589411",
    x"3B587900",
    x"3B585DF3",
    x"3B5842E9",
    x"3B5827E2",
    x"3B580CDF",
    x"3B57F1DF",
    x"3B57D6E2",
    x"3B57BBE9",
    x"3B57A0F3",
    x"3B578601",
    x"3B576B12",
    x"3B575026",
    x"3B57353E",
    x"3B571A59",
    x"3B56FF77",
    x"3B56E499",
    x"3B56C9BE",
    x"3B56AEE7",
    x"3B569412",
    x"3B567942",
    x"3B565E74",
    x"3B5643AA",
    x"3B5628E3",
    x"3B560E20",
    x"3B55F360",
    x"3B55D8A3",
    x"3B55BDEA",
    x"3B55A333",
    x"3B558881",
    x"3B556DD1",
    x"3B555325",
    x"3B55387D",
    x"3B551DD7",
    x"3B550335",
    x"3B54E896",
    x"3B54CDFB",
    x"3B54B363",
    x"3B5498CE",
    x"3B547E3D",
    x"3B5463AF",
    x"3B544924",
    x"3B542E9C",
    x"3B541418",
    x"3B53F997",
    x"3B53DF1A",
    x"3B53C49F",
    x"3B53AA28",
    x"3B538FB5",
    x"3B537545",
    x"3B535AD8",
    x"3B53406E",
    x"3B532607",
    x"3B530BA4",
    x"3B52F145",
    x"3B52D6E8",
    x"3B52BC8F",
    x"3B52A239",
    x"3B5287E6",
    x"3B526D97",
    x"3B52534B",
    x"3B523902",
    x"3B521EBD",
    x"3B52047A",
    x"3B51EA3B",
    x"3B51D000",
    x"3B51B5C7",
    x"3B519B92",
    x"3B518161",
    x"3B516732",
    x"3B514D07",
    x"3B5132DF",
    x"3B5118BA",
    x"3B50FE99",
    x"3B50E47A",
    x"3B50CA60",
    x"3B50B048",
    x"3B509633",
    x"3B507C22",
    x"3B506214",
    x"3B50480A",
    x"3B502E02",
    x"3B5013FE",
    x"3B4FF9FD",
    x"3B4FE000",
    x"3B4FC605",
    x"3B4FAC0E",
    x"3B4F921A",
    x"3B4F782A",
    x"3B4F5E3C",
    x"3B4F4452",
    x"3B4F2A6B",
    x"3B4F1088",
    x"3B4EF6A7",
    x"3B4EDCCA",
    x"3B4EC2F0",
    x"3B4EA919",
    x"3B4E8F46",
    x"3B4E7575",
    x"3B4E5BA8",
    x"3B4E41DE",
    x"3B4E2818",
    x"3B4E0E54",
    x"3B4DF494",
    x"3B4DDAD7",
    x"3B4DC11E",
    x"3B4DA767",
    x"3B4D8DB4",
    x"3B4D7404",
    x"3B4D5A57",
    x"3B4D40AD",
    x"3B4D2706",
    x"3B4D0D63",
    x"3B4CF3C3",
    x"3B4CDA26",
    x"3B4CC08D",
    x"3B4CA6F6",
    x"3B4C8D63",
    x"3B4C73D3",
    x"3B4C5A46",
    x"3B4C40BC",
    x"3B4C2736",
    x"3B4C0DB2",
    x"3B4BF432",
    x"3B4BDAB5",
    x"3B4BC13C",
    x"3B4BA7C5",
    x"3B4B8E52",
    x"3B4B74E1",
    x"3B4B5B74",
    x"3B4B420B",
    x"3B4B28A4",
    x"3B4B0F40",
    x"3B4AF5E0",
    x"3B4ADC83",
    x"3B4AC329",
    x"3B4AA9D2",
    x"3B4A907F",
    x"3B4A772E",
    x"3B4A5DE1",
    x"3B4A4497",
    x"3B4A2B50",
    x"3B4A120C",
    x"3B49F8CB",
    x"3B49DF8E",
    x"3B49C653",
    x"3B49AD1C",
    x"3B4993E8",
    x"3B497AB7",
    x"3B496189",
    x"3B49485F",
    x"3B492F37",
    x"3B491613",
    x"3B48FCF2",
    x"3B48E3D4",
    x"3B48CAB9",
    x"3B48B1A1",
    x"3B48988C",
    x"3B487F7B",
    x"3B48666C",
    x"3B484D61",
    x"3B483459",
    x"3B481B54",
    x"3B480252",
    x"3B47E953",
    x"3B47D058",
    x"3B47B75F",
    x"3B479E6A",
    x"3B478578",
    x"3B476C89",
    x"3B47539D",
    x"3B473AB4",
    x"3B4721CE",
    x"3B4708EB",
    x"3B46F00C",
    x"3B46D72F",
    x"3B46BE56",
    x"3B46A580",
    x"3B468CAD",
    x"3B4673DD",
    x"3B465B10",
    x"3B464246",
    x"3B46297F",
    x"3B4610BB",
    x"3B45F7FB",
    x"3B45DF3D",
    x"3B45C683",
    x"3B45ADCC",
    x"3B459518",
    x"3B457C67",
    x"3B4563B9",
    x"3B454B0E",
    x"3B453266",
    x"3B4519C1",
    x"3B45011F",
    x"3B44E881",
    x"3B44CFE5",
    x"3B44B74D",
    x"3B449EB7",
    x"3B448625",
    x"3B446D96",
    x"3B44550A",
    x"3B443C81",
    x"3B4423FB",
    x"3B440B78",
    x"3B43F2F8",
    x"3B43DA7B",
    x"3B43C201",
    x"3B43A98A",
    x"3B439117",
    x"3B4378A6",
    x"3B436039",
    x"3B4347CE",
    x"3B432F67",
    x"3B431702",
    x"3B42FEA1",
    x"3B42E642",
    x"3B42CDE7",
    x"3B42B58F",
    x"3B429D3A",
    x"3B4284E8",
    x"3B426C99",
    x"3B42544D",
    x"3B423C04",
    x"3B4223BE",
    x"3B420B7B",
    x"3B41F33B",
    x"3B41DAFE",
    x"3B41C2C4",
    x"3B41AA8D",
    x"3B419259",
    x"3B417A29",
    x"3B4161FB",
    x"3B4149D0",
    x"3B4131A8",
    x"3B411984",
    x"3B410162",
    x"3B40E943",
    x"3B40D128",
    x"3B40B90F",
    x"3B40A0F9",
    x"3B4088E7",
    x"3B4070D7",
    x"3B4058CB",
    x"3B4040C1",
    x"3B4028BA",
    x"3B4010B7",
    x"3B3FF8B6",
    x"3B3FE0B9",
    x"3B3FC8BE",
    x"3B3FB0C6",
    x"3B3F98D2",
    x"3B3F80E0",
    x"3B3F68F2",
    x"3B3F5106",
    x"3B3F391D",
    x"3B3F2138",
    x"3B3F0955",
    x"3B3EF175",
    x"3B3ED999",
    x"3B3EC1BF",
    x"3B3EA9E8",
    x"3B3E9214",
    x"3B3E7A44",
    x"3B3E6276",
    x"3B3E4AAB",
    x"3B3E32E3",
    x"3B3E1B1E",
    x"3B3E035C",
    x"3B3DEB9D",
    x"3B3DD3E2",
    x"3B3DBC29",
    x"3B3DA472",
    x"3B3D8CBF",
    x"3B3D750F",
    x"3B3D5D62",
    x"3B3D45B8",
    x"3B3D2E11",
    x"3B3D166C",
    x"3B3CFECB",
    x"3B3CE72D",
    x"3B3CCF91",
    x"3B3CB7F9",
    x"3B3CA063",
    x"3B3C88D1",
    x"3B3C7141",
    x"3B3C59B4",
    x"3B3C422B",
    x"3B3C2AA4",
    x"3B3C1320",
    x"3B3BFB9F",
    x"3B3BE421",
    x"3B3BCCA6",
    x"3B3BB52E",
    x"3B3B9DB9",
    x"3B3B8647",
    x"3B3B6ED7",
    x"3B3B576B",
    x"3B3B4001",
    x"3B3B289B",
    x"3B3B1137",
    x"3B3AF9D7",
    x"3B3AE279",
    x"3B3ACB1E",
    x"3B3AB3C6",
    x"3B3A9C71",
    x"3B3A851F",
    x"3B3A6DD0",
    x"3B3A5683",
    x"3B3A3F3A",
    x"3B3A27F4",
    x"3B3A10B0",
    x"3B39F96F",
    x"3B39E232",
    x"3B39CAF7",
    x"3B39B3BF",
    x"3B399C8A",
    x"3B398558",
    x"3B396E29",
    x"3B3956FC",
    x"3B393FD3",
    x"3B3928AC",
    x"3B391189",
    x"3B38FA68",
    x"3B38E34A",
    x"3B38CC2F",
    x"3B38B517",
    x"3B389E02",
    x"3B3886F0",
    x"3B386FE0",
    x"3B3858D4",
    x"3B3841CA",
    x"3B382AC3",
    x"3B3813BF",
    x"3B37FCBE",
    x"3B37E5C0",
    x"3B37CEC5",
    x"3B37B7CC",
    x"3B37A0D7",
    x"3B3789E4",
    x"3B3772F4",
    x"3B375C07",
    x"3B37451D",
    x"3B372E36",
    x"3B371752",
    x"3B370070",
    x"3B36E992",
    x"3B36D2B6",
    x"3B36BBDD",
    x"3B36A507",
    x"3B368E34",
    x"3B367763",
    x"3B366096",
    x"3B3649CB",
    x"3B363303",
    x"3B361C3E",
    x"3B36057C",
    x"3B35EEBD",
    x"3B35D801",
    x"3B35C147",
    x"3B35AA90",
    x"3B3593DC",
    x"3B357D2B",
    x"3B35667D",
    x"3B354FD2",
    x"3B353929",
    x"3B352283",
    x"3B350BE1",
    x"3B34F540",
    x"3B34DEA3",
    x"3B34C809",
    x"3B34B171",
    x"3B349ADC",
    x"3B34844B",
    x"3B346DBB",
    x"3B34572F",
    x"3B3440A6",
    x"3B342A1F",
    x"3B34139B",
    x"3B33FD1A",
    x"3B33E69C",
    x"3B33D020",
    x"3B33B9A8",
    x"3B33A332",
    x"3B338CBF",
    x"3B33764F",
    x"3B335FE1",
    x"3B334977",
    x"3B33330F",
    x"3B331CAA",
    x"3B330648",
    x"3B32EFE8",
    x"3B32D98C",
    x"3B32C332",
    x"3B32ACDB",
    x"3B329687",
    x"3B328035",
    x"3B3269E7",
    x"3B32539B",
    x"3B323D52",
    x"3B32270C",
    x"3B3210C8",
    x"3B31FA87",
    x"3B31E44A",
    x"3B31CE0E",
    x"3B31B7D6",
    x"3B31A1A0",
    x"3B318B6E",
    x"3B31753E",
    x"3B315F10",
    x"3B3148E6",
    x"3B3132BE",
    x"3B311C99",
    x"3B310677",
    x"3B30F057",
    x"3B30DA3B",
    x"3B30C421",
    x"3B30AE0A",
    x"3B3097F5",
    x"3B3081E4",
    x"3B306BD5",
    x"3B3055C9",
    x"3B303FC0",
    x"3B3029B9",
    x"3B3013B5",
    x"3B2FFDB4",
    x"3B2FE7B6",
    x"3B2FD1BA",
    x"3B2FBBC1",
    x"3B2FA5CB",
    x"3B2F8FD8",
    x"3B2F79E7",
    x"3B2F63F9",
    x"3B2F4E0E",
    x"3B2F3826",
    x"3B2F2240",
    x"3B2F0C5D",
    x"3B2EF67D",
    x"3B2EE0A0",
    x"3B2ECAC5",
    x"3B2EB4ED",
    x"3B2E9F18",
    x"3B2E8945",
    x"3B2E7375",
    x"3B2E5DA8",
    x"3B2E47DE",
    x"3B2E3216",
    x"3B2E1C51",
    x"3B2E068F",
    x"3B2DF0D0",
    x"3B2DDB13",
    x"3B2DC559",
    x"3B2DAFA2",
    x"3B2D99ED",
    x"3B2D843B",
    x"3B2D6E8C",
    x"3B2D58E0",
    x"3B2D4336",
    x"3B2D2D8F",
    x"3B2D17EA",
    x"3B2D0249",
    x"3B2CECAA",
    x"3B2CD70E",
    x"3B2CC174",
    x"3B2CABDD",
    x"3B2C9649",
    x"3B2C80B8",
    x"3B2C6B29",
    x"3B2C559D",
    x"3B2C4014",
    x"3B2C2A8D",
    x"3B2C1509",
    x"3B2BFF88",
    x"3B2BEA09",
    x"3B2BD48D",
    x"3B2BBF14",
    x"3B2BA99D",
    x"3B2B9429",
    x"3B2B7EB8",
    x"3B2B694A",
    x"3B2B53DE",
    x"3B2B3E75",
    x"3B2B290E",
    x"3B2B13AB",
    x"3B2AFE49",
    x"3B2AE8EB",
    x"3B2AD38F",
    x"3B2ABE36",
    x"3B2AA8E0",
    x"3B2A938C",
    x"3B2A7E3B",
    x"3B2A68EC",
    x"3B2A53A1",
    x"3B2A3E57",
    x"3B2A2911",
    x"3B2A13CD",
    x"3B29FE8C",
    x"3B29E94D",
    x"3B29D412",
    x"3B29BED8",
    x"3B29A9A2",
    x"3B29946E",
    x"3B297F3D",
    x"3B296A0E",
    x"3B2954E2",
    x"3B293FB9",
    x"3B292A92",
    x"3B29156E",
    x"3B29004D",
    x"3B28EB2E",
    x"3B28D612",
    x"3B28C0F9",
    x"3B28ABE2",
    x"3B2896CE",
    x"3B2881BC",
    x"3B286CAD",
    x"3B2857A1",
    x"3B284297",
    x"3B282D90",
    x"3B28188C",
    x"3B28038A",
    x"3B27EE8B",
    x"3B27D98F",
    x"3B27C495",
    x"3B27AF9E",
    x"3B279AA9",
    x"3B2785B7",
    x"3B2770C7",
    x"3B275BDB",
    x"3B2746F1",
    x"3B273209",
    x"3B271D24",
    x"3B270842",
    x"3B26F362",
    x"3B26DE85",
    x"3B26C9AA",
    x"3B26B4D2",
    x"3B269FFD",
    x"3B268B2A",
    x"3B26765A",
    x"3B26618D",
    x"3B264CC2",
    x"3B2637FA",
    x"3B262334",
    x"3B260E71",
    x"3B25F9B0",
    x"3B25E4F2",
    x"3B25D037",
    x"3B25BB7E",
    x"3B25A6C8",
    x"3B259215",
    x"3B257D64",
    x"3B2568B5",
    x"3B25540A",
    x"3B253F60",
    x"3B252ABA",
    x"3B251616",
    x"3B250174",
    x"3B24ECD5",
    x"3B24D839",
    x"3B24C39F",
    x"3B24AF08",
    x"3B249A73",
    x"3B2485E1",
    x"3B247152",
    x"3B245CC5",
    x"3B24483B",
    x"3B2433B3",
    x"3B241F2E",
    x"3B240AAB",
    x"3B23F62B",
    x"3B23E1AE",
    x"3B23CD33",
    x"3B23B8BA",
    x"3B23A445",
    x"3B238FD1",
    x"3B237B61",
    x"3B2366F2",
    x"3B235287",
    x"3B233E1E",
    x"3B2329B7",
    x"3B231553",
    x"3B2300F2",
    x"3B22EC93",
    x"3B22D837",
    x"3B22C3DD",
    x"3B22AF86",
    x"3B229B31",
    x"3B2286DF",
    x"3B227290",
    x"3B225E42",
    x"3B2249F8",
    x"3B2235B0",
    x"3B22216B",
    x"3B220D28",
    x"3B21F8E7",
    x"3B21E4A9",
    x"3B21D06E",
    x"3B21BC35",
    x"3B21A7FF",
    x"3B2193CB",
    x"3B217F9A",
    x"3B216B6B",
    x"3B21573F",
    x"3B214316",
    x"3B212EEE",
    x"3B211ACA",
    x"3B2106A8",
    x"3B20F288",
    x"3B20DE6B",
    x"3B20CA51",
    x"3B20B639",
    x"3B20A223",
    x"3B208E10",
    x"3B207A00",
    x"3B2065F2",
    x"3B2051E6",
    x"3B203DDD",
    x"3B2029D7",
    x"3B2015D3",
    x"3B2001D1",
    x"3B1FEDD2",
    x"3B1FD9D6",
    x"3B1FC5DC",
    x"3B1FB1E4",
    x"3B1F9DEF",
    x"3B1F89FD",
    x"3B1F760D",
    x"3B1F621F",
    x"3B1F4E34",
    x"3B1F3A4C",
    x"3B1F2666",
    x"3B1F1282",
    x"3B1EFEA1",
    x"3B1EEAC2",
    x"3B1ED6E6",
    x"3B1EC30D",
    x"3B1EAF36",
    x"3B1E9B61",
    x"3B1E878F",
    x"3B1E73BF",
    x"3B1E5FF2",
    x"3B1E4C27",
    x"3B1E385F",
    x"3B1E2499",
    x"3B1E10D6",
    x"3B1DFD15",
    x"3B1DE956",
    x"3B1DD59A",
    x"3B1DC1E1",
    x"3B1DAE2A",
    x"3B1D9A75",
    x"3B1D86C3",
    x"3B1D7314",
    x"3B1D5F66",
    x"3B1D4BBC",
    x"3B1D3814",
    x"3B1D246E",
    x"3B1D10CA",
    x"3B1CFD2A",
    x"3B1CE98B",
    x"3B1CD5EF",
    x"3B1CC256",
    x"3B1CAEBF",
    x"3B1C9B2A",
    x"3B1C8798",
    x"3B1C7408",
    x"3B1C607B",
    x"3B1C4CF0",
    x"3B1C3968",
    x"3B1C25E2",
    x"3B1C125E",
    x"3B1BFEDD",
    x"3B1BEB5E",
    x"3B1BD7E2",
    x"3B1BC468",
    x"3B1BB0F1",
    x"3B1B9D7C",
    x"3B1B8A0A",
    x"3B1B769A",
    x"3B1B632C",
    x"3B1B4FC1",
    x"3B1B3C58",
    x"3B1B28F2",
    x"3B1B158E",
    x"3B1B022C",
    x"3B1AEECD",
    x"3B1ADB71",
    x"3B1AC816",
    x"3B1AB4BF",
    x"3B1AA169",
    x"3B1A8E16",
    x"3B1A7AC6",
    x"3B1A6778",
    x"3B1A542C",
    x"3B1A40E3",
    x"3B1A2D9C",
    x"3B1A1A57",
    x"3B1A0715",
    x"3B19F3D5",
    x"3B19E098",
    x"3B19CD5D",
    x"3B19BA25",
    x"3B19A6EF",
    x"3B1993BB",
    x"3B19808A",
    x"3B196D5B",
    x"3B195A2E",
    x"3B194704",
    x"3B1933DD",
    x"3B1920B7",
    x"3B190D95",
    x"3B18FA74",
    x"3B18E756",
    x"3B18D43A",
    x"3B18C121",
    x"3B18AE0A",
    x"3B189AF5",
    x"3B1887E3",
    x"3B1874D3",
    x"3B1861C6",
    x"3B184EBB",
    x"3B183BB2",
    x"3B1828AC",
    x"3B1815A8",
    x"3B1802A7",
    x"3B17EFA7",
    x"3B17DCAB",
    x"3B17C9B0",
    x"3B17B6B8",
    x"3B17A3C3",
    x"3B1790CF",
    x"3B177DDE",
    x"3B176AF0",
    x"3B175804",
    x"3B17451A",
    x"3B173232",
    x"3B171F4D",
    x"3B170C6B",
    x"3B16F98A",
    x"3B16E6AC",
    x"3B16D3D1",
    x"3B16C0F7",
    x"3B16AE20",
    x"3B169B4C",
    x"3B168879",
    x"3B1675AA",
    x"3B1662DC",
    x"3B165011",
    x"3B163D48",
    x"3B162A82",
    x"3B1617BD",
    x"3B1604FC",
    x"3B15F23C",
    x"3B15DF7F",
    x"3B15CCC4",
    x"3B15BA0C",
    x"3B15A756",
    x"3B1594A2",
    x"3B1581F1",
    x"3B156F42",
    x"3B155C95",
    x"3B1549EA",
    x"3B153742",
    x"3B15249D",
    x"3B1511F9",
    x"3B14FF58",
    x"3B14ECB9",
    x"3B14DA1D",
    x"3B14C783",
    x"3B14B4EB",
    x"3B14A256",
    x"3B148FC2",
    x"3B147D32",
    x"3B146AA3",
    x"3B145817",
    x"3B14458D",
    x"3B143306",
    x"3B142080",
    x"3B140DFD",
    x"3B13FB7D",
    x"3B13E8FF",
    x"3B13D683",
    x"3B13C409",
    x"3B13B192",
    x"3B139F1D",
    x"3B138CAA",
    x"3B137A39",
    x"3B1367CB",
    x"3B13555F",
    x"3B1342F6",
    x"3B13308F",
    x"3B131E2A",
    x"3B130BC7",
    x"3B12F967",
    x"3B12E709",
    x"3B12D4AD",
    x"3B12C254",
    x"3B12AFFC",
    x"3B129DA8",
    x"3B128B55",
    x"3B127905",
    x"3B1266B7",
    x"3B12546B",
    x"3B124222",
    x"3B122FDB",
    x"3B121D96",
    x"3B120B53",
    x"3B11F913",
    x"3B11E6D5",
    x"3B11D499",
    x"3B11C260",
    x"3B11B029",
    x"3B119DF4",
    x"3B118BC1",
    x"3B117991",
    x"3B116763",
    x"3B115537",
    x"3B11430D",
    x"3B1130E6",
    x"3B111EC1",
    x"3B110C9E",
    x"3B10FA7E",
    x"3B10E860",
    x"3B10D644",
    x"3B10C42A",
    x"3B10B213",
    x"3B109FFE",
    x"3B108DEB",
    x"3B107BDA",
    x"3B1069CC",
    x"3B1057C0",
    x"3B1045B6",
    x"3B1033AE",
    x"3B1021A9",
    x"3B100FA6",
    x"3B0FFDA5",
    x"3B0FEBA7",
    x"3B0FD9AA",
    x"3B0FC7B0",
    x"3B0FB5B8",
    x"3B0FA3C3",
    x"3B0F91CF",
    x"3B0F7FDE",
    x"3B0F6DEF",
    x"3B0F5C03",
    x"3B0F4A18",
    x"3B0F3830",
    x"3B0F264A",
    x"3B0F1467",
    x"3B0F0285",
    x"3B0EF0A6",
    x"3B0EDEC9",
    x"3B0ECCEE",
    x"3B0EBB16",
    x"3B0EA940",
    x"3B0E976C",
    x"3B0E859A",
    x"3B0E73CA",
    x"3B0E61FD",
    x"3B0E5032",
    x"3B0E3E69",
    x"3B0E2CA2",
    x"3B0E1ADE",
    x"3B0E091B",
    x"3B0DF75B",
    x"3B0DE59E",
    x"3B0DD3E2",
    x"3B0DC229",
    x"3B0DB071",
    x"3B0D9EBC",
    x"3B0D8D0A",
    x"3B0D7B59",
    x"3B0D69AB",
    x"3B0D57FF",
    x"3B0D4655",
    x"3B0D34AD",
    x"3B0D2308",
    x"3B0D1164",
    x"3B0CFFC3",
    x"3B0CEE24",
    x"3B0CDC88",
    x"3B0CCAED",
    x"3B0CB955",
    x"3B0CA7BF",
    x"3B0C962B",
    x"3B0C8499",
    x"3B0C730A",
    x"3B0C617D",
    x"3B0C4FF2",
    x"3B0C3E69",
    x"3B0C2CE2",
    x"3B0C1B5E",
    x"3B0C09DB",
    x"3B0BF85B",
    x"3B0BE6DD",
    x"3B0BD561",
    x"3B0BC3E8",
    x"3B0BB270",
    x"3B0BA0FB",
    x"3B0B8F88",
    x"3B0B7E17",
    x"3B0B6CA9",
    x"3B0B5B3C",
    x"3B0B49D2",
    x"3B0B386A",
    x"3B0B2704",
    x"3B0B15A0",
    x"3B0B043E",
    x"3B0AF2DF",
    x"3B0AE182",
    x"3B0AD026",
    x"3B0ABECD",
    x"3B0AAD77",
    x"3B0A9C22",
    x"3B0A8AD0",
    x"3B0A797F",
    x"3B0A6831",
    x"3B0A56E5",
    x"3B0A459C",
    x"3B0A3454",
    x"3B0A230F",
    x"3B0A11CB",
    x"3B0A008A",
    x"3B09EF4B",
    x"3B09DE0E",
    x"3B09CCD4",
    x"3B09BB9B",
    x"3B09AA65",
    x"3B099930",
    x"3B0987FE",
    x"3B0976CE",
    x"3B0965A1",
    x"3B095475",
    x"3B09434C",
    x"3B093224",
    x"3B0920FF",
    x"3B090FDC",
    x"3B08FEBB",
    x"3B08ED9C",
    x"3B08DC80",
    x"3B08CB65",
    x"3B08BA4D",
    x"3B08A937",
    x"3B089822",
    x"3B088711",
    x"3B087601",
    x"3B0864F3",
    x"3B0853E7",
    x"3B0842DE",
    x"3B0831D7",
    x"3B0820D2",
    x"3B080FCF",
    x"3B07FECE",
    x"3B07EDCF",
    x"3B07DCD2",
    x"3B07CBD8",
    x"3B07BADF",
    x"3B07A9E9",
    x"3B0798F5",
    x"3B078803",
    x"3B077713",
    x"3B076625",
    x"3B075539",
    x"3B074450",
    x"3B073368",
    x"3B072283",
    x"3B0711A0",
    x"3B0700BE",
    x"3B06EFDF",
    x"3B06DF02",
    x"3B06CE28",
    x"3B06BD4F",
    x"3B06AC78",
    x"3B069BA4",
    x"3B068AD1",
    x"3B067A01",
    x"3B066933",
    x"3B065867",
    x"3B06479D",
    x"3B0636D5",
    x"3B06260F",
    x"3B06154B",
    x"3B06048A",
    x"3B05F3CA",
    x"3B05E30D",
    x"3B05D251",
    x"3B05C198",
    x"3B05B0E1",
    x"3B05A02C",
    x"3B058F79",
    x"3B057EC8",
    x"3B056E19",
    x"3B055D6D",
    x"3B054CC2",
    x"3B053C19",
    x"3B052B73",
    x"3B051ACF",
    x"3B050A2C",
    x"3B04F98C",
    x"3B04E8EE",
    x"3B04D852",
    x"3B04C7B8",
    x"3B04B720",
    x"3B04A68A",
    x"3B0495F6",
    x"3B048564",
    x"3B0474D5",
    x"3B046447",
    x"3B0453BC",
    x"3B044332",
    x"3B0432AB",
    x"3B042226",
    x"3B0411A2",
    x"3B040121",
    x"3B03F0A2",
    x"3B03E025",
    x"3B03CFAA",
    x"3B03BF31",
    x"3B03AEBA",
    x"3B039E45",
    x"3B038DD3",
    x"3B037D62",
    x"3B036CF3",
    x"3B035C87",
    x"3B034C1C",
    x"3B033BB4",
    x"3B032B4D",
    x"3B031AE9",
    x"3B030A87",
    x"3B02FA26",
    x"3B02E9C8",
    x"3B02D96C",
    x"3B02C912",
    x"3B02B8BA",
    x"3B02A864",
    x"3B02980F",
    x"3B0287BE",
    x"3B02776E",
    x"3B026720",
    x"3B0256D4",
    x"3B02468A",
    x"3B023642",
    x"3B0225FC",
    x"3B0215B9",
    x"3B020577",
    x"3B01F537",
    x"3B01E4FA",
    x"3B01D4BE",
    x"3B01C484",
    x"3B01B44D",
    x"3B01A417",
    x"3B0193E4",
    x"3B0183B2",
    x"3B017383",
    x"3B016356",
    x"3B01532A",
    x"3B014301",
    x"3B0132D9",
    x"3B0122B4",
    x"3B011291",
    x"3B01026F",
    x"3B00F250",
    x"3B00E233",
    x"3B00D218",
    x"3B00C1FE",
    x"3B00B1E7",
    x"3B00A1D2",
    x"3B0091BF",
    x"3B0081AD",
    x"3B00719E",
    x"3B006191",
    x"3B005186",
    x"3B00417D",
    x"3B003175",
    x"3B002170",
    x"3B00116D",
    x"3B00016C",
    x"3AFFE2D9",
    x"3AFFC2DF",
    x"3AFFA2E9",
    x"3AFF82F6",
    x"3AFF6308",
    x"3AFF431E",
    x"3AFF2337",
    x"3AFF0355",
    x"3AFEE376",
    x"3AFEC39C",
    x"3AFEA3C5",
    x"3AFE83F3",
    x"3AFE6424",
    x"3AFE445A",
    x"3AFE2493",
    x"3AFE04D1",
    x"3AFDE512",
    x"3AFDC557",
    x"3AFDA5A1",
    x"3AFD85EE",
    x"3AFD663F",
    x"3AFD4694",
    x"3AFD26EE",
    x"3AFD074B",
    x"3AFCE7AC",
    x"3AFCC811",
    x"3AFCA87A",
    x"3AFC88E7",
    x"3AFC6958",
    x"3AFC49CC",
    x"3AFC2A45",
    x"3AFC0AC2",
    x"3AFBEB42",
    x"3AFBCBC7",
    x"3AFBAC4F",
    x"3AFB8CDC",
    x"3AFB6D6C",
    x"3AFB4E01",
    x"3AFB2E99",
    x"3AFB0F35",
    x"3AFAEFD5",
    x"3AFAD079",
    x"3AFAB121",
    x"3AFA91CD",
    x"3AFA727C",
    x"3AFA5330",
    x"3AFA33E8",
    x"3AFA14A3",
    x"3AF9F562",
    x"3AF9D626",
    x"3AF9B6ED",
    x"3AF997B8",
    x"3AF97887",
    x"3AF9595A",
    x"3AF93A31",
    x"3AF91B0B",
    x"3AF8FBEA",
    x"3AF8DCCC",
    x"3AF8BDB3",
    x"3AF89E9D",
    x"3AF87F8B",
    x"3AF8607D",
    x"3AF84173",
    x"3AF8226D",
    x"3AF8036A",
    x"3AF7E46C",
    x"3AF7C571",
    x"3AF7A67A",
    x"3AF78788",
    x"3AF76899",
    x"3AF749AD",
    x"3AF72AC6",
    x"3AF70BE3",
    x"3AF6ED03",
    x"3AF6CE27",
    x"3AF6AF50",
    x"3AF6907C",
    x"3AF671AC",
    x"3AF652DF",
    x"3AF63417",
    x"3AF61552",
    x"3AF5F691",
    x"3AF5D7D5",
    x"3AF5B91C",
    x"3AF59A66",
    x"3AF57BB5",
    x"3AF55D07",
    x"3AF53E5E",
    x"3AF51FB8",
    x"3AF50116",
    x"3AF4E277",
    x"3AF4C3DD",
    x"3AF4A547",
    x"3AF486B4",
    x"3AF46825",
    x"3AF4499A",
    x"3AF42B12",
    x"3AF40C8F",
    x"3AF3EE0F",
    x"3AF3CF93",
    x"3AF3B11B",
    x"3AF392A7",
    x"3AF37437",
    x"3AF355CA",
    x"3AF33761",
    x"3AF318FC",
    x"3AF2FA9B",
    x"3AF2DC3E",
    x"3AF2BDE4",
    x"3AF29F8E",
    x"3AF2813C",
    x"3AF262EE",
    x"3AF244A3",
    x"3AF2265D",
    x"3AF2081A",
    x"3AF1E9DB",
    x"3AF1CB9F",
    x"3AF1AD68",
    x"3AF18F34",
    x"3AF17104",
    x"3AF152D8",
    x"3AF134AF",
    x"3AF1168B",
    x"3AF0F86A",
    x"3AF0DA4C",
    x"3AF0BC33",
    x"3AF09E1D",
    x"3AF0800C",
    x"3AF061FD",
    x"3AF043F3",
    x"3AF025EC",
    x"3AF007EA",
    x"3AEFE9EA",
    x"3AEFCBEF",
    x"3AEFADF7",
    x"3AEF9004",
    x"3AEF7213",
    x"3AEF5427",
    x"3AEF363E",
    x"3AEF1859",
    x"3AEEFA78",
    x"3AEEDC9B",
    x"3AEEBEC1",
    x"3AEEA0EB",
    x"3AEE8319",
    x"3AEE654A",
    x"3AEE4780",
    x"3AEE29B9",
    x"3AEE0BF5",
    x"3AEDEE36",
    x"3AEDD07A",
    x"3AEDB2C1",
    x"3AED950D",
    x"3AED775C",
    x"3AED59AF",
    x"3AED3C06",
    x"3AED1E60",
    x"3AED00BE",
    x"3AECE320",
    x"3AECC585",
    x"3AECA7EF",
    x"3AEC8A5B",
    x"3AEC6CCC",
    x"3AEC4F40",
    x"3AEC31B8",
    x"3AEC1434",
    x"3AEBF6B3",
    x"3AEBD936",
    x"3AEBBBBD",
    x"3AEB9E47",
    x"3AEB80D5",
    x"3AEB6367",
    x"3AEB45FC",
    x"3AEB2895",
    x"3AEB0B32",
    x"3AEAEDD3",
    x"3AEAD077",
    x"3AEAB31E",
    x"3AEA95CA",
    x"3AEA7879",
    x"3AEA5B2C",
    x"3AEA3DE2",
    x"3AEA209C",
    x"3AEA035A",
    x"3AE9E61C",
    x"3AE9C8E1",
    x"3AE9ABA9",
    x"3AE98E76",
    x"3AE97146",
    x"3AE95419",
    x"3AE936F1",
    x"3AE919CC",
    x"3AE8FCAA",
    x"3AE8DF8C",
    x"3AE8C272",
    x"3AE8A55C",
    x"3AE88849",
    x"3AE86B3A",
    x"3AE84E2E",
    x"3AE83126",
    x"3AE81422",
    x"3AE7F721",
    x"3AE7DA24",
    x"3AE7BD2B",
    x"3AE7A035",
    x"3AE78343",
    x"3AE76654",
    x"3AE74969",
    x"3AE72C82",
    x"3AE70F9E",
    x"3AE6F2BE",
    x"3AE6D5E1",
    x"3AE6B908",
    x"3AE69C33",
    x"3AE67F61",
    x"3AE66293",
    x"3AE645C9",
    x"3AE62902",
    x"3AE60C3E",
    x"3AE5EF7F",
    x"3AE5D2C2",
    x"3AE5B60A",
    x"3AE59955",
    x"3AE57CA4",
    x"3AE55FF6",
    x"3AE5434C",
    x"3AE526A5",
    x"3AE50A02",
    x"3AE4ED62",
    x"3AE4D0C7",
    x"3AE4B42E",
    x"3AE4979A",
    x"3AE47B08",
    x"3AE45E7B",
    x"3AE441F1",
    x"3AE4256A",
    x"3AE408E7",
    x"3AE3EC68",
    x"3AE3CFEC",
    x"3AE3B374",
    x"3AE396FF",
    x"3AE37A8E",
    x"3AE35E21",
    x"3AE341B7",
    x"3AE32550",
    x"3AE308ED",
    x"3AE2EC8E",
    x"3AE2D032",
    x"3AE2B3DA",
    x"3AE29785",
    x"3AE27B34",
    x"3AE25EE7",
    x"3AE2429C",
    x"3AE22656",
    x"3AE20A13",
    x"3AE1EDD3",
    x"3AE1D197",
    x"3AE1B55F",
    x"3AE1992A",
    x"3AE17CF9",
    x"3AE160CB",
    x"3AE144A0",
    x"3AE1287A",
    x"3AE10C56",
    x"3AE0F037",
    x"3AE0D41A",
    x"3AE0B802",
    x"3AE09BEC",
    x"3AE07FDB",
    x"3AE063CC",
    x"3AE047C2",
    x"3AE02BBA",
    x"3AE00FB7",
    x"3ADFF3B6",
    x"3ADFD7BA",
    x"3ADFBBC1",
    x"3ADF9FCB",
    x"3ADF83D9",
    x"3ADF67EA",
    x"3ADF4BFF",
    x"3ADF3017",
    x"3ADF1433",
    x"3ADEF852",
    x"3ADEDC75",
    x"3ADEC09B",
    x"3ADEA4C4",
    x"3ADE88F2",
    x"3ADE6D22",
    x"3ADE5156",
    x"3ADE358E",
    x"3ADE19C9",
    x"3ADDFE07",
    x"3ADDE249",
    x"3ADDC68F",
    x"3ADDAAD8",
    x"3ADD8F24",
    x"3ADD7374",
    x"3ADD57C7",
    x"3ADD3C1E",
    x"3ADD2078",
    x"3ADD04D6",
    x"3ADCE937",
    x"3ADCCD9C",
    x"3ADCB204",
    x"3ADC966F",
    x"3ADC7ADE",
    x"3ADC5F50",
    x"3ADC43C6",
    x"3ADC283F",
    x"3ADC0CBC",
    x"3ADBF13C",
    x"3ADBD5C0",
    x"3ADBBA47",
    x"3ADB9ED1",
    x"3ADB835F",
    x"3ADB67F0",
    x"3ADB4C85",
    x"3ADB311D",
    x"3ADB15B9",
    x"3ADAFA58",
    x"3ADADEFA",
    x"3ADAC3A0",
    x"3ADAA849",
    x"3ADA8CF6",
    x"3ADA71A6",
    x"3ADA565A",
    x"3ADA3B10",
    x"3ADA1FCB",
    x"3ADA0489",
    x"3AD9E94A",
    x"3AD9CE0E",
    x"3AD9B2D6",
    x"3AD997A1",
    x"3AD97C70",
    x"3AD96142",
    x"3AD94618",
    x"3AD92AF1",
    x"3AD90FCD",
    x"3AD8F4AD",
    x"3AD8D990",
    x"3AD8BE76",
    x"3AD8A360",
    x"3AD8884E",
    x"3AD86D3E",
    x"3AD85232",
    x"3AD8372A",
    x"3AD81C25",
    x"3AD80123",
    x"3AD7E624",
    x"3AD7CB29",
    x"3AD7B031",
    x"3AD7953D",
    x"3AD77A4C",
    x"3AD75F5F",
    x"3AD74474",
    x"3AD7298D",
    x"3AD70EAA",
    x"3AD6F3CA",
    x"3AD6D8ED",
    x"3AD6BE14",
    x"3AD6A33D",
    x"3AD6886B",
    x"3AD66D9B",
    x"3AD652CF",
    x"3AD63807",
    x"3AD61D41",
    x"3AD6027F",
    x"3AD5E7C1",
    x"3AD5CD05",
    x"3AD5B24D",
    x"3AD59799",
    x"3AD57CE8",
    x"3AD5623A",
    x"3AD5478F",
    x"3AD52CE8",
    x"3AD51244",
    x"3AD4F7A3",
    x"3AD4DD06",
    x"3AD4C26C",
    x"3AD4A7D5",
    x"3AD48D42",
    x"3AD472B2",
    x"3AD45825",
    x"3AD43D9C",
    x"3AD42316",
    x"3AD40893",
    x"3AD3EE14",
    x"3AD3D398",
    x"3AD3B91F",
    x"3AD39EA9",
    x"3AD38437",
    x"3AD369C8",
    x"3AD34F5D",
    x"3AD334F4",
    x"3AD31A8F",
    x"3AD3002E",
    x"3AD2E5CF",
    x"3AD2CB74",
    x"3AD2B11D",
    x"3AD296C8",
    x"3AD27C77",
    x"3AD26229",
    x"3AD247DE",
    x"3AD22D97",
    x"3AD21353",
    x"3AD1F912",
    x"3AD1DED5",
    x"3AD1C49A",
    x"3AD1AA63",
    x"3AD19030",
    x"3AD175FF",
    x"3AD15BD2",
    x"3AD141A8",
    x"3AD12782",
    x"3AD10D5F",
    x"3AD0F33F",
    x"3AD0D922",
    x"3AD0BF08",
    x"3AD0A4F2",
    x"3AD08ADF",
    x"3AD070CF",
    x"3AD056C3",
    x"3AD03CBA",
    x"3AD022B4",
    x"3AD008B1",
    x"3ACFEEB1",
    x"3ACFD4B5",
    x"3ACFBABC",
    x"3ACFA0C7",
    x"3ACF86D4",
    x"3ACF6CE5",
    x"3ACF52F9",
    x"3ACF3910",
    x"3ACF1F2B",
    x"3ACF0548",
    x"3ACEEB69",
    x"3ACED18E",
    x"3ACEB7B5",
    x"3ACE9DE0",
    x"3ACE840D",
    x"3ACE6A3F",
    x"3ACE5073",
    x"3ACE36AA",
    x"3ACE1CE5",
    x"3ACE0323",
    x"3ACDE964",
    x"3ACDCFA9",
    x"3ACDB5F1",
    x"3ACD9C3B",
    x"3ACD8289",
    x"3ACD68DB",
    x"3ACD4F2F",
    x"3ACD3587",
    x"3ACD1BE2",
    x"3ACD0240",
    x"3ACCE8A1",
    x"3ACCCF06",
    x"3ACCB56E",
    x"3ACC9BD8",
    x"3ACC8247",
    x"3ACC68B8",
    x"3ACC4F2C",
    x"3ACC35A4",
    x"3ACC1C1F",
    x"3ACC029D",
    x"3ACBE91E",
    x"3ACBCFA3",
    x"3ACBB62A",
    x"3ACB9CB5",
    x"3ACB8343",
    x"3ACB69D4",
    x"3ACB5069",
    x"3ACB3700",
    x"3ACB1D9B",
    x"3ACB0439",
    x"3ACAEADA",
    x"3ACAD17E",
    x"3ACAB826",
    x"3ACA9ED0",
    x"3ACA857E",
    x"3ACA6C2F",
    x"3ACA52E3",
    x"3ACA399A",
    x"3ACA2054",
    x"3ACA0712",
    x"3AC9EDD3",
    x"3AC9D497",
    x"3AC9BB5E",
    x"3AC9A228",
    x"3AC988F5",
    x"3AC96FC5",
    x"3AC95699",
    x"3AC93D70",
    x"3AC9244A",
    x"3AC90B27",
    x"3AC8F207",
    x"3AC8D8EA",
    x"3AC8BFD1",
    x"3AC8A6BA",
    x"3AC88DA7",
    x"3AC87497",
    x"3AC85B8A",
    x"3AC84280",
    x"3AC82979",
    x"3AC81076",
    x"3AC7F775",
    x"3AC7DE78",
    x"3AC7C57E",
    x"3AC7AC86",
    x"3AC79392",
    x"3AC77AA1",
    x"3AC761B4",
    x"3AC748C9",
    x"3AC72FE2",
    x"3AC716FD",
    x"3AC6FE1C",
    x"3AC6E53E",
    x"3AC6CC62",
    x"3AC6B38A",
    x"3AC69AB6",
    x"3AC681E4",
    x"3AC66915",
    x"3AC6504A",
    x"3AC63781",
    x"3AC61EBC",
    x"3AC605F9",
    x"3AC5ED3A",
    x"3AC5D47E",
    x"3AC5BBC5",
    x"3AC5A30F",
    x"3AC58A5C",
    x"3AC571AD",
    x"3AC55900",
    x"3AC54056",
    x"3AC527B0",
    x"3AC50F0C",
    x"3AC4F66C",
    x"3AC4DDCF",
    x"3AC4C535",
    x"3AC4AC9D",
    x"3AC49409",
    x"3AC47B78",
    x"3AC462EB",
    x"3AC44A60",
    x"3AC431D8",
    x"3AC41953",
    x"3AC400D2",
    x"3AC3E853",
    x"3AC3CFD8",
    x"3AC3B75F",
    x"3AC39EEA",
    x"3AC38677",
    x"3AC36E08",
    x"3AC3559C",
    x"3AC33D33",
    x"3AC324CD",
    x"3AC30C69",
    x"3AC2F409",
    x"3AC2DBAC",
    x"3AC2C352",
    x"3AC2AAFC",
    x"3AC292A8",
    x"3AC27A57",
    x"3AC26209",
    x"3AC249BE",
    x"3AC23177",
    x"3AC21932",
    x"3AC200F0",
    x"3AC1E8B2",
    x"3AC1D076",
    x"3AC1B83E",
    x"3AC1A008",
    x"3AC187D6",
    x"3AC16FA6",
    x"3AC1577A",
    x"3AC13F50",
    x"3AC1272A",
    x"3AC10F07",
    x"3AC0F6E6",
    x"3AC0DEC9",
    x"3AC0C6AF",
    x"3AC0AE97",
    x"3AC09683",
    x"3AC07E72",
    x"3AC06663",
    x"3AC04E58",
    x"3AC03650",
    x"3AC01E4A",
    x"3AC00648",
    x"3ABFEE49",
    x"3ABFD64D",
    x"3ABFBE53",
    x"3ABFA65D",
    x"3ABF8E6A",
    x"3ABF7679",
    x"3ABF5E8C",
    x"3ABF46A2",
    x"3ABF2EBA",
    x"3ABF16D6",
    x"3ABEFEF5",
    x"3ABEE716",
    x"3ABECF3B",
    x"3ABEB762",
    x"3ABE9F8D",
    x"3ABE87BB",
    x"3ABE6FEB",
    x"3ABE581F",
    x"3ABE4055",
    x"3ABE288F",
    x"3ABE10CB",
    x"3ABDF90A",
    x"3ABDE14D",
    x"3ABDC992",
    x"3ABDB1DA",
    x"3ABD9A26",
    x"3ABD8274",
    x"3ABD6AC5",
    x"3ABD5319",
    x"3ABD3B70",
    x"3ABD23CA",
    x"3ABD0C27",
    x"3ABCF487",
    x"3ABCDCEA",
    x"3ABCC550",
    x"3ABCADB9",
    x"3ABC9624",
    x"3ABC7E93",
    x"3ABC6705",
    x"3ABC4F79",
    x"3ABC37F1",
    x"3ABC206B",
    x"3ABC08E9",
    x"3ABBF169",
    x"3ABBD9ED",
    x"3ABBC273",
    x"3ABBAAFC",
    x"3ABB9388",
    x"3ABB7C17",
    x"3ABB64A9",
    x"3ABB4D3E",
    x"3ABB35D6",
    x"3ABB1E70",
    x"3ABB070E",
    x"3ABAEFAF",
    x"3ABAD852",
    x"3ABAC0F9",
    x"3ABAA9A2",
    x"3ABA924E",
    x"3ABA7AFD",
    x"3ABA63AF",
    x"3ABA4C64",
    x"3ABA351C",
    x"3ABA1DD7",
    x"3ABA0695",
    x"3AB9EF55",
    x"3AB9D819",
    x"3AB9C0DF",
    x"3AB9A9A9",
    x"3AB99275",
    x"3AB97B44",
    x"3AB96416",
    x"3AB94CEB",
    x"3AB935C3",
    x"3AB91E9E",
    x"3AB9077B",
    x"3AB8F05C",
    x"3AB8D93F",
    x"3AB8C226",
    x"3AB8AB0F",
    x"3AB893FB",
    x"3AB87CEA",
    x"3AB865DC",
    x"3AB84ED0",
    x"3AB837C8",
    x"3AB820C2",
    x"3AB809C0",
    x"3AB7F2C0",
    x"3AB7DBC3",
    x"3AB7C4C9",
    x"3AB7ADD2",
    x"3AB796DD",
    x"3AB77FEC",
    x"3AB768FD",
    x"3AB75212",
    x"3AB73B29",
    x"3AB72443",
    x"3AB70D60",
    x"3AB6F680",
    x"3AB6DFA2",
    x"3AB6C8C8",
    x"3AB6B1F0",
    x"3AB69B1B",
    x"3AB68449",
    x"3AB66D7A",
    x"3AB656AE",
    x"3AB63FE5",
    x"3AB6291E",
    x"3AB6125A",
    x"3AB5FB99",
    x"3AB5E4DB",
    x"3AB5CE20",
    x"3AB5B768",
    x"3AB5A0B2",
    x"3AB58A00",
    x"3AB57350",
    x"3AB55CA3",
    x"3AB545F9",
    x"3AB52F51",
    x"3AB518AD",
    x"3AB5020B",
    x"3AB4EB6C",
    x"3AB4D4D0",
    x"3AB4BE37",
    x"3AB4A7A1",
    x"3AB4910D",
    x"3AB47A7C",
    x"3AB463EF",
    x"3AB44D63",
    x"3AB436DB",
    x"3AB42056",
    x"3AB409D3",
    x"3AB3F353",
    x"3AB3DCD6",
    x"3AB3C65C",
    x"3AB3AFE5",
    x"3AB39970",
    x"3AB382FE",
    x"3AB36C8F",
    x"3AB35623",
    x"3AB33FBA",
    x"3AB32953",
    x"3AB312F0",
    x"3AB2FC8F",
    x"3AB2E630",
    x"3AB2CFD5",
    x"3AB2B97C",
    x"3AB2A327",
    x"3AB28CD4",
    x"3AB27683",
    x"3AB26036",
    x"3AB249EB",
    x"3AB233A4",
    x"3AB21D5E",
    x"3AB2071C",
    x"3AB1F0DD",
    x"3AB1DAA0",
    x"3AB1C466",
    x"3AB1AE2F",
    x"3AB197FA",
    x"3AB181C9",
    x"3AB16B9A",
    x"3AB1556E",
    x"3AB13F45",
    x"3AB1291E",
    x"3AB112FA",
    x"3AB0FCD9",
    x"3AB0E6BB",
    x"3AB0D0A0",
    x"3AB0BA87",
    x"3AB0A471",
    x"3AB08E5E",
    x"3AB0784D",
    x"3AB06240",
    x"3AB04C35",
    x"3AB0362D",
    x"3AB02027",
    x"3AB00A25",
    x"3AAFF425",
    x"3AAFDE28",
    x"3AAFC82D",
    x"3AAFB236",
    x"3AAF9C41",
    x"3AAF864F",
    x"3AAF705F",
    x"3AAF5A72",
    x"3AAF4489",
    x"3AAF2EA1",
    x"3AAF18BD",
    x"3AAF02DB",
    x"3AAEECFC",
    x"3AAED720",
    x"3AAEC146",
    x"3AAEAB70",
    x"3AAE959C",
    x"3AAE7FCA",
    x"3AAE69FC",
    x"3AAE5430",
    x"3AAE3E67",
    x"3AAE28A0",
    x"3AAE12DC",
    x"3AADFD1B",
    x"3AADE75D",
    x"3AADD1A2",
    x"3AADBBE9",
    x"3AADA633",
    x"3AAD907F",
    x"3AAD7ACE",
    x"3AAD6520",
    x"3AAD4F75",
    x"3AAD39CD",
    x"3AAD2427",
    x"3AAD0E84",
    x"3AACF8E3",
    x"3AACE345",
    x"3AACCDAA",
    x"3AACB812",
    x"3AACA27C",
    x"3AAC8CE9",
    x"3AAC7759",
    x"3AAC61CB",
    x"3AAC4C41",
    x"3AAC36B8",
    x"3AAC2133",
    x"3AAC0BB0",
    x"3AABF630",
    x"3AABE0B3",
    x"3AABCB38",
    x"3AABB5C0",
    x"3AABA04A",
    x"3AAB8AD8",
    x"3AAB7568",
    x"3AAB5FFA",
    x"3AAB4A90",
    x"3AAB3528",
    x"3AAB1FC2",
    x"3AAB0A60",
    x"3AAAF500",
    x"3AAADFA2",
    x"3AAACA48",
    x"3AAAB4F0",
    x"3AAA9F9B",
    x"3AAA8A48",
    x"3AAA74F8",
    x"3AAA5FAB",
    x"3AAA4A60",
    x"3AAA3518",
    x"3AAA1FD3",
    x"3AAA0A90",
    x"3AA9F550",
    x"3AA9E013",
    x"3AA9CAD8",
    x"3AA9B5A0",
    x"3AA9A06B",
    x"3AA98B38",
    x"3AA97608",
    x"3AA960DB",
    x"3AA94BB0",
    x"3AA93688",
    x"3AA92162",
    x"3AA90C3F",
    x"3AA8F71F",
    x"3AA8E202",
    x"3AA8CCE7",
    x"3AA8B7CE",
    x"3AA8A2B9",
    x"3AA88DA6",
    x"3AA87895",
    x"3AA86387",
    x"3AA84E7C",
    x"3AA83974",
    x"3AA8246E",
    x"3AA80F6B",
    x"3AA7FA6A",
    x"3AA7E56C",
    x"3AA7D071",
    x"3AA7BB78",
    x"3AA7A682",
    x"3AA7918E",
    x"3AA77C9E",
    x"3AA767AF",
    x"3AA752C4",
    x"3AA73DDB",
    x"3AA728F4",
    x"3AA71410",
    x"3AA6FF2F",
    x"3AA6EA51",
    x"3AA6D575",
    x"3AA6C09B",
    x"3AA6ABC4",
    x"3AA696F0",
    x"3AA6821F",
    x"3AA66D50",
    x"3AA65883",
    x"3AA643BA",
    x"3AA62EF2",
    x"3AA61A2E",
    x"3AA6056C",
    x"3AA5F0AC",
    x"3AA5DBF0",
    x"3AA5C735",
    x"3AA5B27E",
    x"3AA59DC9",
    x"3AA58916",
    x"3AA57467",
    x"3AA55FB9",
    x"3AA54B0F",
    x"3AA53667",
    x"3AA521C1",
    x"3AA50D1E",
    x"3AA4F87E",
    x"3AA4E3E0",
    x"3AA4CF45",
    x"3AA4BAAC",
    x"3AA4A616",
    x"3AA49183",
    x"3AA47CF2",
    x"3AA46863",
    x"3AA453D8",
    x"3AA43F4E",
    x"3AA42AC8",
    x"3AA41644",
    x"3AA401C2",
    x"3AA3ED43",
    x"3AA3D8C7",
    x"3AA3C44D",
    x"3AA3AFD6",
    x"3AA39B61",
    x"3AA386EF",
    x"3AA3727F",
    x"3AA35E12",
    x"3AA349A8",
    x"3AA33540",
    x"3AA320DB",
    x"3AA30C78",
    x"3AA2F817",
    x"3AA2E3BA",
    x"3AA2CF5F",
    x"3AA2BB06",
    x"3AA2A6B0",
    x"3AA2925C",
    x"3AA27E0B",
    x"3AA269BD",
    x"3AA25571",
    x"3AA24127",
    x"3AA22CE0",
    x"3AA2189C",
    x"3AA2045A",
    x"3AA1F01B",
    x"3AA1DBDE",
    x"3AA1C7A4",
    x"3AA1B36C",
    x"3AA19F37",
    x"3AA18B05",
    x"3AA176D4",
    x"3AA162A7",
    x"3AA14E7C",
    x"3AA13A53",
    x"3AA1262D",
    x"3AA1120A",
    x"3AA0FDE9",
    x"3AA0E9CA",
    x"3AA0D5AE",
    x"3AA0C195",
    x"3AA0AD7E",
    x"3AA09969",
    x"3AA08558",
    x"3AA07148",
    x"3AA05D3B",
    x"3AA04931",
    x"3AA03529",
    x"3AA02124",
    x"3AA00D21",
    x"3A9FF920",
    x"3A9FE522",
    x"3A9FD127",
    x"3A9FBD2E",
    x"3A9FA938",
    x"3A9F9544",
    x"3A9F8152",
    x"3A9F6D63",
    x"3A9F5977",
    x"3A9F458D",
    x"3A9F31A6",
    x"3A9F1DC1",
    x"3A9F09DE",
    x"3A9EF5FE",
    x"3A9EE221",
    x"3A9ECE46",
    x"3A9EBA6D",
    x"3A9EA697",
    x"3A9E92C3",
    x"3A9E7EF2",
    x"3A9E6B24",
    x"3A9E5758",
    x"3A9E438E",
    x"3A9E2FC7",
    x"3A9E1C02",
    x"3A9E0840",
    x"3A9DF480",
    x"3A9DE0C3",
    x"3A9DCD08",
    x"3A9DB94F",
    x"3A9DA599",
    x"3A9D91E6",
    x"3A9D7E35",
    x"3A9D6A86",
    x"3A9D56DA",
    x"3A9D4331",
    x"3A9D2F89",
    x"3A9D1BE5",
    x"3A9D0842",
    x"3A9CF4A3",
    x"3A9CE105",
    x"3A9CCD6A",
    x"3A9CB9D2",
    x"3A9CA63C",
    x"3A9C92A8",
    x"3A9C7F17",
    x"3A9C6B89",
    x"3A9C57FC",
    x"3A9C4473",
    x"3A9C30EB",
    x"3A9C1D66",
    x"3A9C09E4",
    x"3A9BF664",
    x"3A9BE2E6",
    x"3A9BCF6B",
    x"3A9BBBF2",
    x"3A9BA87C",
    x"3A9B9508",
    x"3A9B8197",
    x"3A9B6E28",
    x"3A9B5ABB",
    x"3A9B4751",
    x"3A9B33EA",
    x"3A9B2084",
    x"3A9B0D21",
    x"3A9AF9C1",
    x"3A9AE663",
    x"3A9AD307",
    x"3A9ABFAE",
    x"3A9AAC57",
    x"3A9A9903",
    x"3A9A85B1",
    x"3A9A7262",
    x"3A9A5F15",
    x"3A9A4BCA",
    x"3A9A3882",
    x"3A9A253C",
    x"3A9A11F8",
    x"3A99FEB7",
    x"3A99EB79",
    x"3A99D83C",
    x"3A99C503",
    x"3A99B1CB",
    x"3A999E96",
    x"3A998B64",
    x"3A997833",
    x"3A996506",
    x"3A9951DA",
    x"3A993EB1",
    x"3A992B8A",
    x"3A991866",
    x"3A990544",
    x"3A98F225",
    x"3A98DF08",
    x"3A98CBED",
    x"3A98B8D5",
    x"3A98A5BF",
    x"3A9892AB",
    x"3A987F9A",
    x"3A986C8B",
    x"3A98597F",
    x"3A984675",
    x"3A98336D",
    x"3A982068",
    x"3A980D65",
    x"3A97FA65",
    x"3A97E767",
    x"3A97D46B",
    x"3A97C172",
    x"3A97AE7B",
    x"3A979B86",
    x"3A978894",
    x"3A9775A4",
    x"3A9762B6",
    x"3A974FCB",
    x"3A973CE2",
    x"3A9729FC",
    x"3A971718",
    x"3A970436",
    x"3A96F157",
    x"3A96DE7A",
    x"3A96CB9F",
    x"3A96B8C7",
    x"3A96A5F1",
    x"3A96931E",
    x"3A96804C",
    x"3A966D7D",
    x"3A965AB1",
    x"3A9647E7",
    x"3A96351F",
    x"3A962259",
    x"3A960F96",
    x"3A95FCD6",
    x"3A95EA17",
    x"3A95D75B",
    x"3A95C4A1",
    x"3A95B1EA",
    x"3A959F35",
    x"3A958C82",
    x"3A9579D2",
    x"3A956724",
    x"3A955478",
    x"3A9541CF",
    x"3A952F27",
    x"3A951C83",
    x"3A9509E0",
    x"3A94F740",
    x"3A94E4A3",
    x"3A94D207",
    x"3A94BF6E",
    x"3A94ACD7",
    x"3A949A43",
    x"3A9487B1",
    x"3A947521",
    x"3A946293",
    x"3A945008",
    x"3A943D7F",
    x"3A942AF9",
    x"3A941875",
    x"3A9405F3",
    x"3A93F373",
    x"3A93E0F6",
    x"3A93CE7B",
    x"3A93BC02",
    x"3A93A98C",
    x"3A939718",
    x"3A9384A6",
    x"3A937237",
    x"3A935FCA",
    x"3A934D5F",
    x"3A933AF6",
    x"3A932890",
    x"3A93162C",
    x"3A9303CA",
    x"3A92F16B",
    x"3A92DF0E",
    x"3A92CCB3",
    x"3A92BA5B",
    x"3A92A805",
    x"3A9295B1",
    x"3A92835F",
    x"3A927110",
    x"3A925EC3",
    x"3A924C78",
    x"3A923A30",
    x"3A9227EA",
    x"3A9215A6",
    x"3A920364",
    x"3A91F125",
    x"3A91DEE8",
    x"3A91CCAD",
    x"3A91BA75",
    x"3A91A83F",
    x"3A91960B",
    x"3A9183D9",
    x"3A9171AA",
    x"3A915F7D",
    x"3A914D52",
    x"3A913B2A",
    x"3A912903",
    x"3A9116DF",
    x"3A9104BE",
    x"3A90F29E",
    x"3A90E081",
    x"3A90CE66",
    x"3A90BC4D",
    x"3A90AA37",
    x"3A909823",
    x"3A908611",
    x"3A907401",
    x"3A9061F4",
    x"3A904FE9",
    x"3A903DE0",
    x"3A902BD9",
    x"3A9019D5",
    x"3A9007D3",
    x"3A8FF5D3",
    x"3A8FE3D5",
    x"3A8FD1DA",
    x"3A8FBFE1",
    x"3A8FADEA",
    x"3A8F9BF5",
    x"3A8F8A03",
    x"3A8F7813",
    x"3A8F6625",
    x"3A8F5439",
    x"3A8F4250",
    x"3A8F3069",
    x"3A8F1E84",
    x"3A8F0CA1",
    x"3A8EFAC1",
    x"3A8EE8E3",
    x"3A8ED707",
    x"3A8EC52D",
    x"3A8EB355",
    x"3A8EA180",
    x"3A8E8FAD",
    x"3A8E7DDC",
    x"3A8E6C0D",
    x"3A8E5A41",
    x"3A8E4877",
    x"3A8E36AF",
    x"3A8E24E9",
    x"3A8E1326",
    x"3A8E0164",
    x"3A8DEFA5",
    x"3A8DDDE8",
    x"3A8DCC2E",
    x"3A8DBA75",
    x"3A8DA8BF",
    x"3A8D970B",
    x"3A8D8559",
    x"3A8D73AA",
    x"3A8D61FD",
    x"3A8D5051",
    x"3A8D3EA8",
    x"3A8D2D02",
    x"3A8D1B5D",
    x"3A8D09BB",
    x"3A8CF81B",
    x"3A8CE67D",
    x"3A8CD4E1",
    x"3A8CC348",
    x"3A8CB1B0",
    x"3A8CA01B",
    x"3A8C8E88",
    x"3A8C7CF8",
    x"3A8C6B69",
    x"3A8C59DD",
    x"3A8C4853",
    x"3A8C36CB",
    x"3A8C2545",
    x"3A8C13C1",
    x"3A8C0240",
    x"3A8BF0C1",
    x"3A8BDF44",
    x"3A8BCDC9",
    x"3A8BBC50",
    x"3A8BAADA",
    x"3A8B9966",
    x"3A8B87F4",
    x"3A8B7684",
    x"3A8B6516",
    x"3A8B53AA",
    x"3A8B4241",
    x"3A8B30DA",
    x"3A8B1F75",
    x"3A8B0E12",
    x"3A8AFCB1",
    x"3A8AEB53",
    x"3A8AD9F6",
    x"3A8AC89C",
    x"3A8AB744",
    x"3A8AA5EE",
    x"3A8A949B",
    x"3A8A8349",
    x"3A8A71FA",
    x"3A8A60AD",
    x"3A8A4F62",
    x"3A8A3E19",
    x"3A8A2CD2",
    x"3A8A1B8E",
    x"3A8A0A4B",
    x"3A89F90B",
    x"3A89E7CD",
    x"3A89D691",
    x"3A89C557",
    x"3A89B420",
    x"3A89A2EA",
    x"3A8991B7",
    x"3A898086",
    x"3A896F57",
    x"3A895E2A",
    x"3A894CFF",
    x"3A893BD7",
    x"3A892AB1",
    x"3A89198C",
    x"3A89086A",
    x"3A88F74A",
    x"3A88E62C",
    x"3A88D511",
    x"3A88C3F7",
    x"3A88B2E0",
    x"3A88A1CA",
    x"3A8890B7",
    x"3A887FA6",
    x"3A886E97",
    x"3A885D8A",
    x"3A884C80",
    x"3A883B77",
    x"3A882A71",
    x"3A88196D",
    x"3A88086B",
    x"3A87F76B",
    x"3A87E66D",
    x"3A87D571",
    x"3A87C477",
    x"3A87B380",
    x"3A87A28B",
    x"3A879197",
    x"3A8780A6",
    x"3A876FB7",
    x"3A875ECA",
    x"3A874DDF",
    x"3A873CF7",
    x"3A872C10",
    x"3A871B2C",
    x"3A870A49",
    x"3A86F969",
    x"3A86E88B",
    x"3A86D7AF",
    x"3A86C6D5",
    x"3A86B5FD",
    x"3A86A528",
    x"3A869454",
    x"3A868383",
    x"3A8672B3",
    x"3A8661E6",
    x"3A86511B",
    x"3A864052",
    x"3A862F8B",
    x"3A861EC6",
    x"3A860E03",
    x"3A85FD42",
    x"3A85EC84",
    x"3A85DBC7",
    x"3A85CB0D",
    x"3A85BA54",
    x"3A85A99E",
    x"3A8598EA",
    x"3A858838",
    x"3A857788",
    x"3A8566DA",
    x"3A85562E",
    x"3A854584",
    x"3A8534DD",
    x"3A852437",
    x"3A851394",
    x"3A8502F2",
    x"3A84F253",
    x"3A84E1B6",
    x"3A84D11B",
    x"3A84C081",
    x"3A84AFEA",
    x"3A849F55",
    x"3A848EC3",
    x"3A847E32",
    x"3A846DA3",
    x"3A845D16",
    x"3A844C8C",
    x"3A843C03",
    x"3A842B7D",
    x"3A841AF8",
    x"3A840A76",
    x"3A83F9F6",
    x"3A83E978",
    x"3A83D8FB",
    x"3A83C881",
    x"3A83B809",
    x"3A83A793",
    x"3A83971F",
    x"3A8386AD",
    x"3A83763E",
    x"3A8365D0",
    x"3A835564",
    x"3A8344FB",
    x"3A833493",
    x"3A83242D",
    x"3A8313CA",
    x"3A830368",
    x"3A82F309",
    x"3A82E2AC",
    x"3A82D250",
    x"3A82C1F7",
    x"3A82B1A0",
    x"3A82A14B",
    x"3A8290F8",
    x"3A8280A6",
    x"3A827057",
    x"3A82600A",
    x"3A824FBF",
    x"3A823F76",
    x"3A822F30",
    x"3A821EEB",
    x"3A820EA8",
    x"3A81FE67",
    x"3A81EE28",
    x"3A81DDEB",
    x"3A81CDB1",
    x"3A81BD78",
    x"3A81AD41",
    x"3A819D0D",
    x"3A818CDA",
    x"3A817CAA",
    x"3A816C7B",
    x"3A815C4E",
    x"3A814C24",
    x"3A813BFB",
    x"3A812BD5",
    x"3A811BB0",
    x"3A810B8E",
    x"3A80FB6E",
    x"3A80EB4F",
    x"3A80DB33",
    x"3A80CB18",
    x"3A80BB00",
    x"3A80AAEA",
    x"3A809AD5",
    x"3A808AC3",
    x"3A807AB3",
    x"3A806AA4",
    x"3A805A98",
    x"3A804A8E",
    x"3A803A85",
    x"3A802A7F",
    x"3A801A7B",
    x"3A800A78",
    x"3A7FF4F0",
    x"3A7FD4F3",
    x"3A7FB4FB",
    x"3A7F9506",
    x"3A7F7515",
    x"3A7F5529",
    x"3A7F3540",
    x"3A7F155B",
    x"3A7EF57B",
    x"3A7ED59E",
    x"3A7EB5C5",
    x"3A7E95F1",
    x"3A7E7620",
    x"3A7E5653",
    x"3A7E368A",
    x"3A7E16C5",
    x"3A7DF705",
    x"3A7DD748",
    x"3A7DB78F",
    x"3A7D97DA",
    x"3A7D7829",
    x"3A7D587C",
    x"3A7D38D3",
    x"3A7D192E",
    x"3A7CF98C",
    x"3A7CD9EF",
    x"3A7CBA56",
    x"3A7C9AC1",
    x"3A7C7B2F",
    x"3A7C5BA2",
    x"3A7C3C18",
    x"3A7C1C93",
    x"3A7BFD11",
    x"3A7BDD94",
    x"3A7BBE1A",
    x"3A7B9EA4",
    x"3A7B7F32",
    x"3A7B5FC4",
    x"3A7B405A",
    x"3A7B20F4",
    x"3A7B0192",
    x"3A7AE234",
    x"3A7AC2D9",
    x"3A7AA383",
    x"3A7A8431",
    x"3A7A64E2",
    x"3A7A4597",
    x"3A7A2651",
    x"3A7A070E",
    x"3A79E7CF",
    x"3A79C894",
    x"3A79A95D",
    x"3A798A29",
    x"3A796AFA",
    x"3A794BCF",
    x"3A792CA7",
    x"3A790D84",
    x"3A78EE64",
    x"3A78CF48",
    x"3A78B030",
    x"3A78911C",
    x"3A78720C",
    x"3A7852FF",
    x"3A7833F7",
    x"3A7814F2",
    x"3A77F5F2",
    x"3A77D6F5",
    x"3A77B7FC",
    x"3A779907",
    x"3A777A16",
    x"3A775B28",
    x"3A773C3F",
    x"3A771D59",
    x"3A76FE78",
    x"3A76DF9A",
    x"3A76C0C0",
    x"3A76A1EA",
    x"3A768317",
    x"3A766449",
    x"3A76457E",
    x"3A7626B7",
    x"3A7607F4",
    x"3A75E935",
    x"3A75CA7A",
    x"3A75ABC3",
    x"3A758D0F",
    x"3A756E5F",
    x"3A754FB4",
    x"3A75310C",
    x"3A751267",
    x"3A74F3C7",
    x"3A74D52A",
    x"3A74B692",
    x"3A7497FD",
    x"3A74796C",
    x"3A745ADE",
    x"3A743C55",
    x"3A741DCF",
    x"3A73FF4E",
    x"3A73E0CF",
    x"3A73C255",
    x"3A73A3DF",
    x"3A73856C",
    x"3A7366FE",
    x"3A734893",
    x"3A732A2B",
    x"3A730BC8",
    x"3A72ED68",
    x"3A72CF0D",
    x"3A72B0B5",
    x"3A729261",
    x"3A727410",
    x"3A7255C3",
    x"3A72377B",
    x"3A721936",
    x"3A71FAF4",
    x"3A71DCB7",
    x"3A71BE7D",
    x"3A71A047",
    x"3A718215",
    x"3A7163E7",
    x"3A7145BC",
    x"3A712795",
    x"3A710972",
    x"3A70EB53",
    x"3A70CD37",
    x"3A70AF20",
    x"3A70910C",
    x"3A7072FB",
    x"3A7054EF",
    x"3A7036E6",
    x"3A7018E1",
    x"3A6FFAE0",
    x"3A6FDCE2",
    x"3A6FBEE9",
    x"3A6FA0F3",
    x"3A6F8300",
    x"3A6F6512",
    x"3A6F4727",
    x"3A6F2940",
    x"3A6F0B5D",
    x"3A6EED7D",
    x"3A6ECFA2",
    x"3A6EB1C9",
    x"3A6E93F5",
    x"3A6E7624",
    x"3A6E5858",
    x"3A6E3A8E",
    x"3A6E1CC9",
    x"3A6DFF07",
    x"3A6DE149",
    x"3A6DC38F",
    x"3A6DA5D8",
    x"3A6D8825",
    x"3A6D6A76",
    x"3A6D4CCB",
    x"3A6D2F23",
    x"3A6D117F",
    x"3A6CF3DF",
    x"3A6CD642",
    x"3A6CB8A9",
    x"3A6C9B14",
    x"3A6C7D82",
    x"3A6C5FF4",
    x"3A6C426A",
    x"3A6C24E4",
    x"3A6C0761",
    x"3A6BE9E2",
    x"3A6BCC67",
    x"3A6BAEEF",
    x"3A6B917B",
    x"3A6B740B",
    x"3A6B569E",
    x"3A6B3935",
    x"3A6B1BD0",
    x"3A6AFE6E",
    x"3A6AE110",
    x"3A6AC3B6",
    x"3A6AA65F",
    x"3A6A890C",
    x"3A6A6BBD",
    x"3A6A4E71",
    x"3A6A3129",
    x"3A6A13E5",
    x"3A69F6A4",
    x"3A69D967",
    x"3A69BC2E",
    x"3A699EF8",
    x"3A6981C6",
    x"3A696498",
    x"3A69476D",
    x"3A692A46",
    x"3A690D22",
    x"3A68F003",
    x"3A68D2E6",
    x"3A68B5CE",
    x"3A6898B9",
    x"3A687BA8",
    x"3A685E9A",
    x"3A684190",
    x"3A68248A",
    x"3A680787",
    x"3A67EA88",
    x"3A67CD8C",
    x"3A67B094",
    x"3A6793A0",
    x"3A6776AF",
    x"3A6759C2",
    x"3A673CD9",
    x"3A671FF3",
    x"3A670311",
    x"3A66E632",
    x"3A66C957",
    x"3A66AC80",
    x"3A668FAC",
    x"3A6672DC",
    x"3A665610",
    x"3A663947",
    x"3A661C81",
    x"3A65FFC0",
    x"3A65E301",
    x"3A65C647",
    x"3A65A990",
    x"3A658CDC",
    x"3A65702D",
    x"3A655380",
    x"3A6536D8",
    x"3A651A33",
    x"3A64FD91",
    x"3A64E0F3",
    x"3A64C459",
    x"3A64A7C2",
    x"3A648B2F",
    x"3A646E9F",
    x"3A645213",
    x"3A64358B",
    x"3A641906",
    x"3A63FC85",
    x"3A63E007",
    x"3A63C38D",
    x"3A63A716",
    x"3A638AA3",
    x"3A636E33",
    x"3A6351C7",
    x"3A63355F",
    x"3A6318FA",
    x"3A62FC99",
    x"3A62E03B",
    x"3A62C3E0",
    x"3A62A78A",
    x"3A628B37",
    x"3A626EE7",
    x"3A62529B",
    x"3A623652",
    x"3A621A0D",
    x"3A61FDCC",
    x"3A61E18E",
    x"3A61C553",
    x"3A61A91D",
    x"3A618CE9",
    x"3A6170B9",
    x"3A61548D",
    x"3A613864",
    x"3A611C3F",
    x"3A61001D",
    x"3A60E3FF",
    x"3A60C7E4",
    x"3A60ABCD",
    x"3A608FB9",
    x"3A6073A9",
    x"3A60579C",
    x"3A603B93",
    x"3A601F8D",
    x"3A60038B",
    x"3A5FE78C",
    x"3A5FCB91",
    x"3A5FAF9A",
    x"3A5F93A5",
    x"3A5F77B5",
    x"3A5F5BC7",
    x"3A5F3FDE",
    x"3A5F23F7",
    x"3A5F0815",
    x"3A5EEC35",
    x"3A5ED05A",
    x"3A5EB481",
    x"3A5E98AD",
    x"3A5E7CDB",
    x"3A5E610D",
    x"3A5E4543",
    x"3A5E297C",
    x"3A5E0DB9",
    x"3A5DF1F9",
    x"3A5DD63C",
    x"3A5DBA83",
    x"3A5D9ECD",
    x"3A5D831B",
    x"3A5D676D",
    x"3A5D4BC1",
    x"3A5D301A",
    x"3A5D1475",
    x"3A5CF8D5",
    x"3A5CDD37",
    x"3A5CC19D",
    x"3A5CA607",
    x"3A5C8A74",
    x"3A5C6EE4",
    x"3A5C5358",
    x"3A5C37CF",
    x"3A5C1C4A",
    x"3A5C00C8",
    x"3A5BE54A",
    x"3A5BC9CF",
    x"3A5BAE57",
    x"3A5B92E3",
    x"3A5B7773",
    x"3A5B5C06",
    x"3A5B409C",
    x"3A5B2535",
    x"3A5B09D2",
    x"3A5AEE73",
    x"3A5AD317",
    x"3A5AB7BE",
    x"3A5A9C69",
    x"3A5A8117",
    x"3A5A65C9",
    x"3A5A4A7E",
    x"3A5A2F36",
    x"3A5A13F2",
    x"3A59F8B1",
    x"3A59DD74",
    x"3A59C23A",
    x"3A59A703",
    x"3A598BD0",
    x"3A5970A0",
    x"3A595574",
    x"3A593A4B",
    x"3A591F25",
    x"3A590403",
    x"3A58E8E4",
    x"3A58CDC9",
    x"3A58B2B1",
    x"3A58979C",
    x"3A587C8B",
    x"3A58617D",
    x"3A584672",
    x"3A582B6B",
    x"3A581068",
    x"3A57F567",
    x"3A57DA6A",
    x"3A57BF71",
    x"3A57A47A",
    x"3A578987",
    x"3A576E98",
    x"3A5753AC",
    x"3A5738C3",
    x"3A571DDE",
    x"3A5702FC",
    x"3A56E81D",
    x"3A56CD42",
    x"3A56B26A",
    x"3A569795",
    x"3A567CC4",
    x"3A5661F6",
    x"3A56472B",
    x"3A562C64",
    x"3A5611A0",
    x"3A55F6E0",
    x"3A55DC22",
    x"3A55C169",
    x"3A55A6B2",
    x"3A558BFF",
    x"3A55714F",
    x"3A5556A3",
    x"3A553BF9",
    x"3A552154",
    x"3A5506B1",
    x"3A54EC12",
    x"3A54D176",
    x"3A54B6DD",
    x"3A549C48",
    x"3A5481B6",
    x"3A546728",
    x"3A544C9D",
    x"3A543215",
    x"3A541790",
    x"3A53FD0F",
    x"3A53E291",
    x"3A53C816",
    x"3A53AD9F",
    x"3A53932B",
    x"3A5378BA",
    x"3A535E4D",
    x"3A5343E2",
    x"3A53297C",
    x"3A530F18",
    x"3A52F4B8",
    x"3A52DA5B",
    x"3A52C001",
    x"3A52A5AB",
    x"3A528B58",
    x"3A527108",
    x"3A5256BC",
    x"3A523C72",
    x"3A52222C",
    x"3A5207EA",
    x"3A51EDAA",
    x"3A51D36E",
    x"3A51B936",
    x"3A519F00",
    x"3A5184CE",
    x"3A516A9F",
    x"3A515073",
    x"3A51364B",
    x"3A511C26",
    x"3A510204",
    x"3A50E7E5",
    x"3A50CDCA",
    x"3A50B3B2",
    x"3A50999D",
    x"3A507F8B",
    x"3A50657D",
    x"3A504B72",
    x"3A50316A",
    x"3A501766",
    x"3A4FFD64",
    x"3A4FE366",
    x"3A4FC96B",
    x"3A4FAF74",
    x"3A4F9580",
    x"3A4F7B8E",
    x"3A4F61A1",
    x"3A4F47B6",
    x"3A4F2DCF",
    x"3A4F13EB",
    x"3A4EFA0A",
    x"3A4EE02C",
    x"3A4EC652",
    x"3A4EAC7B",
    x"3A4E92A7",
    x"3A4E78D6",
    x"3A4E5F08",
    x"3A4E453E",
    x"3A4E2B77",
    x"3A4E11B3",
    x"3A4DF7F3",
    x"3A4DDE35",
    x"3A4DC47B",
    x"3A4DAAC4",
    x"3A4D9110",
    x"3A4D7760",
    x"3A4D5DB3",
    x"3A4D4408",
    x"3A4D2A62",
    x"3A4D10BE",
    x"3A4CF71D",
    x"3A4CDD80",
    x"3A4CC3E6",
    x"3A4CAA4F",
    x"3A4C90BB",
    x"3A4C772B",
    x"3A4C5D9E",
    x"3A4C4414",
    x"3A4C2A8D",
    x"3A4C1109",
    x"3A4BF788",
    x"3A4BDE0B",
    x"3A4BC491",
    x"3A4BAB1A",
    x"3A4B91A6",
    x"3A4B7835",
    x"3A4B5EC8",
    x"3A4B455E",
    x"3A4B2BF7",
    x"3A4B1293",
    x"3A4AF932",
    x"3A4ADFD4",
    x"3A4AC67A",
    x"3A4AAD23",
    x"3A4A93CF",
    x"3A4A7A7E",
    x"3A4A6130",
    x"3A4A47E6",
    x"3A4A2E9E",
    x"3A4A155A",
    x"3A49FC19",
    x"3A49E2DB",
    x"3A49C9A0",
    x"3A49B068",
    x"3A499734",
    x"3A497E03",
    x"3A4964D5",
    x"3A494BA9",
    x"3A493282",
    x"3A49195D",
    x"3A49003B",
    x"3A48E71D",
    x"3A48CE01",
    x"3A48B4E9",
    x"3A489BD4",
    x"3A4882C2",
    x"3A4869B4",
    x"3A4850A8",
    x"3A48379F",
    x"3A481E9A",
    x"3A480598",
    x"3A47EC99",
    x"3A47D39D",
    x"3A47BAA4",
    x"3A47A1AE",
    x"3A4788BB",
    x"3A476FCC",
    x"3A4756DF",
    x"3A473DF6",
    x"3A472510",
    x"3A470C2D",
    x"3A46F34D",
    x"3A46DA70",
    x"3A46C196",
    x"3A46A8C0",
    x"3A468FEC",
    x"3A46771C",
    x"3A465E4E",
    x"3A464584",
    x"3A462CBD",
    x"3A4613F9",
    x"3A45FB38",
    x"3A45E27A",
    x"3A45C9BF",
    x"3A45B108",
    x"3A459853",
    x"3A457FA1",
    x"3A4566F3",
    x"3A454E48",
    x"3A45359F",
    x"3A451CFA",
    x"3A450458",
    x"3A44EBB9",
    x"3A44D31D",
    x"3A44BA84",
    x"3A44A1EF",
    x"3A44895C",
    x"3A4470CC",
    x"3A445840",
    x"3A443FB6",
    x"3A442730",
    x"3A440EAC",
    x"3A43F62C",
    x"3A43DDAF",
    x"3A43C535",
    x"3A43ACBE",
    x"3A43944A",
    x"3A437BD9",
    x"3A43636B",
    x"3A434B00",
    x"3A433298",
    x"3A431A33",
    x"3A4301D1",
    x"3A42E973",
    x"3A42D117",
    x"3A42B8BE",
    x"3A42A069",
    x"3A428816",
    x"3A426FC7",
    x"3A42577A",
    x"3A423F31",
    x"3A4226EA",
    x"3A420EA7",
    x"3A41F667",
    x"3A41DE2A",
    x"3A41C5EF",
    x"3A41ADB8",
    x"3A419584",
    x"3A417D53",
    x"3A416525",
    x"3A414CF9",
    x"3A4134D1",
    x"3A411CAC",
    x"3A41048A",
    x"3A40EC6B",
    x"3A40D44F",
    x"3A40BC36",
    x"3A40A420",
    x"3A408C0D",
    x"3A4073FD",
    x"3A405BF0",
    x"3A4043E6",
    x"3A402BDF",
    x"3A4013DB",
    x"3A3FFBDA",
    x"3A3FE3DC",
    x"3A3FCBE1",
    x"3A3FB3E9",
    x"3A3F9BF4",
    x"3A3F8402",
    x"3A3F6C13",
    x"3A3F5427",
    x"3A3F3C3E",
    x"3A3F2458",
    x"3A3F0C75",
    x"3A3EF495",
    x"3A3EDCB8",
    x"3A3EC4DE",
    x"3A3EAD07",
    x"3A3E9532",
    x"3A3E7D61",
    x"3A3E6593",
    x"3A3E4DC8",
    x"3A3E3600",
    x"3A3E1E3A",
    x"3A3E0678",
    x"3A3DEEB9",
    x"3A3DD6FC",
    x"3A3DBF43",
    x"3A3DA78D",
    x"3A3D8FD9",
    x"3A3D7829",
    x"3A3D607B",
    x"3A3D48D1",
    x"3A3D3129",
    x"3A3D1984",
    x"3A3D01E3",
    x"3A3CEA44",
    x"3A3CD2A8",
    x"3A3CBB0F",
    x"3A3CA379",
    x"3A3C8BE6",
    x"3A3C7456",
    x"3A3C5CC9",
    x"3A3C453F",
    x"3A3C2DB8",
    x"3A3C1634",
    x"3A3BFEB2",
    x"3A3BE734",
    x"3A3BCFB8",
    x"3A3BB840",
    x"3A3BA0CA",
    x"3A3B8958",
    x"3A3B71E8",
    x"3A3B5A7B",
    x"3A3B4311",
    x"3A3B2BAB",
    x"3A3B1447",
    x"3A3AFCE5",
    x"3A3AE587",
    x"3A3ACE2C",
    x"3A3AB6D4",
    x"3A3A9F7E",
    x"3A3A882C",
    x"3A3A70DC",
    x"3A3A5990",
    x"3A3A4246",
    x"3A3A2AFF",
    x"3A3A13BB",
    x"3A39FC7A",
    x"3A39E53C",
    x"3A39CE01",
    x"3A39B6C9",
    x"3A399F93",
    x"3A398861",
    x"3A397131",
    x"3A395A04",
    x"3A3942DB",
    x"3A392BB4",
    x"3A391490",
    x"3A38FD6F",
    x"3A38E650",
    x"3A38CF35",
    x"3A38B81C",
    x"3A38A107",
    x"3A3889F4",
    x"3A3872E4",
    x"3A385BD7",
    x"3A3844CD",
    x"3A382DC6",
    x"3A3816C2",
    x"3A37FFC1",
    x"3A37E8C2",
    x"3A37D1C6",
    x"3A37BACE",
    x"3A37A3D8",
    x"3A378CE5",
    x"3A3775F4",
    x"3A375F07",
    x"3A37481D",
    x"3A373135",
    x"3A371A50",
    x"3A37036F",
    x"3A36EC90",
    x"3A36D5B3",
    x"3A36BEDA",
    x"3A36A804",
    x"3A369130",
    x"3A367A5F",
    x"3A366392",
    x"3A364CC7",
    x"3A3635FE",
    x"3A361F39",
    x"3A360877",
    x"3A35F1B7",
    x"3A35DAFA",
    x"3A35C440",
    x"3A35AD89",
    x"3A3596D5",
    x"3A358023",
    x"3A356975",
    x"3A3552C9",
    x"3A353C20",
    x"3A35257A",
    x"3A350ED7",
    x"3A34F836",
    x"3A34E199",
    x"3A34CAFE",
    x"3A34B466",
    x"3A349DD1",
    x"3A34873E",
    x"3A3470AF",
    x"3A345A22",
    x"3A344398",
    x"3A342D11",
    x"3A34168D",
    x"3A34000C",
    x"3A33E98D",
    x"3A33D311",
    x"3A33BC98",
    x"3A33A622",
    x"3A338FAF",
    x"3A33793E",
    x"3A3362D1",
    x"3A334C66",
    x"3A3335FD",
    x"3A331F98",
    x"3A330936",
    x"3A32F2D6",
    x"3A32DC79",
    x"3A32C61F",
    x"3A32AFC7",
    x"3A329973",
    x"3A328321",
    x"3A326CD2",
    x"3A325686",
    x"3A32403C",
    x"3A3229F6",
    x"3A3213B2",
    x"3A31FD71",
    x"3A31E732",
    x"3A31D0F7",
    x"3A31BABE",
    x"3A31A488",
    x"3A318E55",
    x"3A317825",
    x"3A3161F7",
    x"3A314BCC",
    x"3A3135A4",
    x"3A311F7F",
    x"3A31095C",
    x"3A30F33C",
    x"3A30DD1F",
    x"3A30C705",
    x"3A30B0EE",
    x"3A309AD9",
    x"3A3084C7",
    x"3A306EB8",
    x"3A3058AB",
    x"3A3042A2",
    x"3A302C9B",
    x"3A301696",
    x"3A300095",
    x"3A2FEA96",
    x"3A2FD49A",
    x"3A2FBEA1",
    x"3A2FA8AB",
    x"3A2F92B7",
    x"3A2F7CC6",
    x"3A2F66D8",
    x"3A2F50EC",
    x"3A2F3B03",
    x"3A2F251D",
    x"3A2F0F3A",
    x"3A2EF95A",
    x"3A2EE37C",
    x"3A2ECDA1",
    x"3A2EB7C8",
    x"3A2EA1F3",
    x"3A2E8C20",
    x"3A2E7650",
    x"3A2E6082",
    x"3A2E4AB8",
    x"3A2E34F0",
    x"3A2E1F2A",
    x"3A2E0968",
    x"3A2DF3A8",
    x"3A2DDDEB",
    x"3A2DC831",
    x"3A2DB279",
    x"3A2D9CC4",
    x"3A2D8712",
    x"3A2D7162",
    x"3A2D5BB5",
    x"3A2D460B",
    x"3A2D3064",
    x"3A2D1ABF",
    x"3A2D051D",
    x"3A2CEF7E",
    x"3A2CD9E1",
    x"3A2CC447",
    x"3A2CAEB0",
    x"3A2C991C",
    x"3A2C838A",
    x"3A2C6DFB",
    x"3A2C586F",
    x"3A2C42E5",
    x"3A2C2D5E",
    x"3A2C17D9",
    x"3A2C0258",
    x"3A2BECD9",
    x"3A2BD75D",
    x"3A2BC1E3",
    x"3A2BAC6C",
    x"3A2B96F8",
    x"3A2B8186",
    x"3A2B6C18",
    x"3A2B56AB",
    x"3A2B4142",
    x"3A2B2BDB",
    x"3A2B1677",
    x"3A2B0115",
    x"3A2AEBB7",
    x"3A2AD65B",
    x"3A2AC101",
    x"3A2AABAA",
    x"3A2A9656",
    x"3A2A8105",
    x"3A2A6BB6",
    x"3A2A566A",
    x"3A2A4120",
    x"3A2A2BD9",
    x"3A2A1695",
    x"3A2A0154",
    x"3A29EC15",
    x"3A29D6D9",
    x"3A29C19F",
    x"3A29AC68",
    x"3A299734",
    x"3A298203",
    x"3A296CD4",
    x"3A2957A7",
    x"3A29427E",
    x"3A292D57",
    x"3A291832",
    x"3A290311",
    x"3A28EDF2",
    x"3A28D8D5",
    x"3A28C3BB",
    x"3A28AEA4",
    x"3A289990",
    x"3A28847E",
    x"3A286F6F",
    x"3A285A62",
    x"3A284558",
    x"3A283051",
    x"3A281B4C",
    x"3A28064A",
    x"3A27F14A",
    x"3A27DC4E",
    x"3A27C753",
    x"3A27B25C",
    x"3A279D67",
    x"3A278874",
    x"3A277385",
    x"3A275E97",
    x"3A2749AD",
    x"3A2734C5",
    x"3A271FE0",
    x"3A270AFD",
    x"3A26F61D",
    x"3A26E140",
    x"3A26CC65",
    x"3A26B78C",
    x"3A26A2B7",
    x"3A268DE4",
    x"3A267913",
    x"3A266446",
    x"3A264F7A",
    x"3A263AB2",
    x"3A2625EC",
    x"3A261128",
    x"3A25FC67",
    x"3A25E7A9",
    x"3A25D2ED",
    x"3A25BE34",
    x"3A25A97E",
    x"3A2594CA",
    x"3A258019",
    x"3A256B6A",
    x"3A2556BE",
    x"3A254214",
    x"3A252D6D",
    x"3A2518C9",
    x"3A250427",
    x"3A24EF88",
    x"3A24DAEB",
    x"3A24C651",
    x"3A24B1BA",
    x"3A249D25",
    x"3A248892",
    x"3A247403",
    x"3A245F75",
    x"3A244AEB",
    x"3A243663",
    x"3A2421DD",
    x"3A240D5A",
    x"3A23F8DA",
    x"3A23E45C",
    x"3A23CFE1",
    x"3A23BB68",
    x"3A23A6F2",
    x"3A23927E",
    x"3A237E0D",
    x"3A23699F",
    x"3A235533",
    x"3A2340C9",
    x"3A232C63",
    x"3A2317FE",
    x"3A23039D",
    x"3A22EF3D",
    x"3A22DAE1",
    x"3A22C687",
    x"3A22B22F",
    x"3A229DDA",
    x"3A228988",
    x"3A227538",
    x"3A2260EA",
    x"3A224CA0",
    x"3A223857",
    x"3A222411",
    x"3A220FCE",
    x"3A21FB8D",
    x"3A21E74F",
    x"3A21D314",
    x"3A21BEDB",
    x"3A21AAA4",
    x"3A219670",
    x"3A21823E",
    x"3A216E0F",
    x"3A2159E3",
    x"3A2145B9",
    x"3A213191",
    x"3A211D6C",
    x"3A21094A",
    x"3A20F52A",
    x"3A20E10D",
    x"3A20CCF2",
    x"3A20B8DA",
    x"3A20A4C4",
    x"3A2090B0",
    x"3A207C9F",
    x"3A206891",
    x"3A205485",
    x"3A20407C",
    x"3A202C75",
    x"3A201871",
    x"3A20046F",
    x"3A1FF070",
    x"3A1FDC73",
    x"3A1FC879",
    x"3A1FB481",
    x"3A1FA08C",
    x"3A1F8C99",
    x"3A1F78A8",
    x"3A1F64BB",
    x"3A1F50CF",
    x"3A1F3CE6",
    x"3A1F2900",
    x"3A1F151C",
    x"3A1F013B",
    x"3A1EED5C",
    x"3A1ED97F",
    x"3A1EC5A5",
    x"3A1EB1CE",
    x"3A1E9DF9",
    x"3A1E8A26",
    x"3A1E7656",
    x"3A1E6289",
    x"3A1E4EBE",
    x"3A1E3AF5",
    x"3A1E272F",
    x"3A1E136B",
    x"3A1DFFAA",
    x"3A1DEBEC",
    x"3A1DD82F",
    x"3A1DC475",
    x"3A1DB0BE",
    x"3A1D9D09",
    x"3A1D8957",
    x"3A1D75A7",
    x"3A1D61F9",
    x"3A1D4E4E",
    x"3A1D3AA6",
    x"3A1D2700",
    x"3A1D135C",
    x"3A1CFFBB",
    x"3A1CEC1C",
    x"3A1CD880",
    x"3A1CC4E6",
    x"3A1CB14F",
    x"3A1C9DBA",
    x"3A1C8A27",
    x"3A1C7697",
    x"3A1C630A",
    x"3A1C4F7E",
    x"3A1C3BF6",
    x"3A1C286F",
    x"3A1C14EC",
    x"3A1C016A",
    x"3A1BEDEB",
    x"3A1BDA6F",
    x"3A1BC6F5",
    x"3A1BB37D",
    x"3A1BA008",
    x"3A1B8C95",
    x"3A1B7925",
    x"3A1B65B7",
    x"3A1B524B",
    x"3A1B3EE2",
    x"3A1B2B7B",
    x"3A1B1817",
    x"3A1B04B5",
    x"3A1AF156",
    x"3A1ADDF9",
    x"3A1ACA9F",
    x"3A1AB746",
    x"3A1AA3F1",
    x"3A1A909D",
    x"3A1A7D4D",
    x"3A1A69FE",
    x"3A1A56B2",
    x"3A1A4368",
    x"3A1A3021",
    x"3A1A1CDC",
    x"3A1A099A",
    x"3A19F65A",
    x"3A19E31C",
    x"3A19CFE1",
    x"3A19BCA9",
    x"3A19A972",
    x"3A19963E",
    x"3A19830D",
    x"3A196FDD",
    x"3A195CB1",
    x"3A194986",
    x"3A19365E",
    x"3A192339",
    x"3A191015",
    x"3A18FCF5",
    x"3A18E9D6",
    x"3A18D6BA",
    x"3A18C3A0",
    x"3A18B089",
    x"3A189D74",
    x"3A188A62",
    x"3A187752",
    x"3A186444",
    x"3A185139",
    x"3A183E30",
    x"3A182B29",
    x"3A181825",
    x"3A180523",
    x"3A17F224",
    x"3A17DF27",
    x"3A17CC2C",
    x"3A17B934",
    x"3A17A63E",
    x"3A17934A",
    x"3A178059",
    x"3A176D6A",
    x"3A175A7D",
    x"3A174793",
    x"3A1734AB",
    x"3A1721C6",
    x"3A170EE3",
    x"3A16FC02",
    x"3A16E924",
    x"3A16D648",
    x"3A16C36E",
    x"3A16B097",
    x"3A169DC2",
    x"3A168AF0",
    x"3A167820",
    x"3A166552",
    x"3A165286",
    x"3A163FBD",
    x"3A162CF6",
    x"3A161A32",
    x"3A160770",
    x"3A15F4B0",
    x"3A15E1F3",
    x"3A15CF38",
    x"3A15BC7F",
    x"3A15A9C8",
    x"3A159714",
    x"3A158463",
    x"3A1571B3",
    x"3A155F06",
    x"3A154C5C",
    x"3A1539B3",
    x"3A15270D",
    x"3A151469",
    x"3A1501C8",
    x"3A14EF29",
    x"3A14DC8C",
    x"3A14C9F2",
    x"3A14B75A",
    x"3A14A4C4",
    x"3A149231",
    x"3A147F9F",
    x"3A146D11",
    x"3A145A84",
    x"3A1447FA",
    x"3A143572",
    x"3A1422ED",
    x"3A141069",
    x"3A13FDE9",
    x"3A13EB6A",
    x"3A13D8EE",
    x"3A13C674",
    x"3A13B3FC",
    x"3A13A187",
    x"3A138F14",
    x"3A137CA3",
    x"3A136A34",
    x"3A1357C8",
    x"3A13455F",
    x"3A1332F7",
    x"3A132092",
    x"3A130E2F",
    x"3A12FBCE",
    x"3A12E970",
    x"3A12D714",
    x"3A12C4BA",
    x"3A12B263",
    x"3A12A00E",
    x"3A128DBB",
    x"3A127B6A",
    x"3A12691C",
    x"3A1256D0",
    x"3A124486",
    x"3A12323F",
    x"3A121FFA",
    x"3A120DB7",
    x"3A11FB76",
    x"3A11E938",
    x"3A11D6FC",
    x"3A11C4C2",
    x"3A11B28B",
    x"3A11A055",
    x"3A118E23",
    x"3A117BF2",
    x"3A1169C4",
    x"3A115798",
    x"3A11456E",
    x"3A113346",
    x"3A112121",
    x"3A110EFE",
    x"3A10FCDD",
    x"3A10EABF",
    x"3A10D8A2",
    x"3A10C688",
    x"3A10B471",
    x"3A10A25B",
    x"3A109048",
    x"3A107E37",
    x"3A106C29",
    x"3A105A1C",
    x"3A104812",
    x"3A10360A",
    x"3A102405",
    x"3A101201",
    x"3A100000",
    x"3A0FEE01",
    x"3A0FDC05",
    x"3A0FCA0A",
    x"3A0FB812",
    x"3A0FA61C",
    x"3A0F9429",
    x"3A0F8237",
    x"3A0F7048",
    x"3A0F5E5B",
    x"3A0F4C70",
    x"3A0F3A88",
    x"3A0F28A2",
    x"3A0F16BE",
    x"3A0F04DC",
    x"3A0EF2FD",
    x"3A0EE11F",
    x"3A0ECF44",
    x"3A0EBD6C",
    x"3A0EAB95",
    x"3A0E99C1",
    x"3A0E87EF",
    x"3A0E761F",
    x"3A0E6451",
    x"3A0E5286",
    x"3A0E40BC",
    x"3A0E2EF5",
    x"3A0E1D31",
    x"3A0E0B6E",
    x"3A0DF9AE",
    x"3A0DE7F0",
    x"3A0DD634",
    x"3A0DC47A",
    x"3A0DB2C3",
    x"3A0DA10D",
    x"3A0D8F5A",
    x"3A0D7DAA",
    x"3A0D6BFB",
    x"3A0D5A4F",
    x"3A0D48A4",
    x"3A0D36FC",
    x"3A0D2557",
    x"3A0D13B3",
    x"3A0D0212",
    x"3A0CF073",
    x"3A0CDED6",
    x"3A0CCD3B",
    x"3A0CBBA2",
    x"3A0CAA0C",
    x"3A0C9878",
    x"3A0C86E6",
    x"3A0C7556",
    x"3A0C63C9",
    x"3A0C523D",
    x"3A0C40B4",
    x"3A0C2F2D",
    x"3A0C1DA8",
    x"3A0C0C26",
    x"3A0BFAA5",
    x"3A0BE927",
    x"3A0BD7AB",
    x"3A0BC631",
    x"3A0BB4B9",
    x"3A0BA344",
    x"3A0B91D0",
    x"3A0B805F",
    x"3A0B6EF0",
    x"3A0B5D84",
    x"3A0B4C19",
    x"3A0B3AB1",
    x"3A0B294A",
    x"3A0B17E6",
    x"3A0B0684",
    x"3A0AF525",
    x"3A0AE3C7",
    x"3A0AD26C",
    x"3A0AC112",
    x"3A0AAFBB",
    x"3A0A9E67",
    x"3A0A8D14",
    x"3A0A7BC3",
    x"3A0A6A75",
    x"3A0A5929",
    x"3A0A47DF",
    x"3A0A3697",
    x"3A0A2551",
    x"3A0A140D",
    x"3A0A02CC",
    x"3A09F18D",
    x"3A09E050",
    x"3A09CF15",
    x"3A09BDDC",
    x"3A09ACA5",
    x"3A099B71",
    x"3A098A3E",
    x"3A09790E",
    x"3A0967E0",
    x"3A0956B4",
    x"3A09458A",
    x"3A093463",
    x"3A09233D",
    x"3A09121A",
    x"3A0900F9",
    x"3A08EFDA",
    x"3A08DEBD",
    x"3A08CDA2",
    x"3A08BC89",
    x"3A08AB73",
    x"3A089A5E",
    x"3A08894C",
    x"3A08783C",
    x"3A08672E",
    x"3A085622",
    x"3A084519",
    x"3A083411",
    x"3A08230C",
    x"3A081208",
    x"3A080107",
    x"3A07F008",
    x"3A07DF0B",
    x"3A07CE10",
    x"3A07BD18",
    x"3A07AC21",
    x"3A079B2D",
    x"3A078A3A",
    x"3A07794A",
    x"3A07685C",
    x"3A075770",
    x"3A074686",
    x"3A07359E",
    x"3A0724B9",
    x"3A0713D5",
    x"3A0702F4",
    x"3A06F214",
    x"3A06E137",
    x"3A06D05C",
    x"3A06BF83",
    x"3A06AEAC",
    x"3A069DD7",
    x"3A068D05",
    x"3A067C34",
    x"3A066B66",
    x"3A065A99",
    x"3A0649CF",
    x"3A063907",
    x"3A062841",
    x"3A06177D",
    x"3A0606BB",
    x"3A05F5FB",
    x"3A05E53D",
    x"3A05D482",
    x"3A05C3C8",
    x"3A05B311",
    x"3A05A25C",
    x"3A0591A8",
    x"3A0580F7",
    x"3A057048",
    x"3A055F9B",
    x"3A054EF0",
    x"3A053E47",
    x"3A052DA1",
    x"3A051CFC",
    x"3A050C59",
    x"3A04FBB9",
    x"3A04EB1A",
    x"3A04DA7E",
    x"3A04C9E4",
    x"3A04B94C",
    x"3A04A8B5",
    x"3A049821",
    x"3A04878F",
    x"3A0476FF",
    x"3A046672",
    x"3A0455E6",
    x"3A04455C",
    x"3A0434D5",
    x"3A04244F",
    x"3A0413CB",
    x"3A04034A",
    x"3A03F2CB",
    x"3A03E24D",
    x"3A03D1D2",
    x"3A03C159",
    x"3A03B0E2",
    x"3A03A06D",
    x"3A038FFA",
    x"3A037F89",
    x"3A036F1A",
    x"3A035EAD",
    x"3A034E42",
    x"3A033DD9",
    x"3A032D73",
    x"3A031D0E",
    x"3A030CAB",
    x"3A02FC4B",
    x"3A02EBEC",
    x"3A02DB90",
    x"3A02CB35",
    x"3A02BADD",
    x"3A02AA87",
    x"3A029A32",
    x"3A0289E0",
    x"3A027990",
    x"3A026942",
    x"3A0258F6",
    x"3A0248AB",
    x"3A023863",
    x"3A02281D",
    x"3A0217D9",
    x"3A020797",
    x"3A01F757",
    x"3A01E71A",
    x"3A01D6DE",
    x"3A01C6A4",
    x"3A01B66C",
    x"3A01A636",
    x"3A019602",
    x"3A0185D1",
    x"3A0175A1",
    x"3A016573",
    x"3A015548",
    x"3A01451E",
    x"3A0134F6",
    x"3A0124D1",
    x"3A0114AD",
    x"3A01048C",
    x"3A00F46C",
    x"3A00E44E",
    x"3A00D433",
    x"3A00C419",
    x"3A00B402",
    x"3A00A3EC",
    x"3A0093D9",
    x"3A0083C7",
    x"3A0073B8",
    x"3A0063AB",
    x"3A00539F",
    x"3A004396",
    x"3A00338E",
    x"3A002389",
    x"3A001385",
    x"3A000384",
    x"39FFE709",
    x"39FFC70E",
    x"39FFA717",
    x"39FF8724",
    x"39FF6735",
    x"39FF474A",
    x"39FF2763",
    x"39FF0781",
    x"39FEE7A2",
    x"39FEC7C7",
    x"39FEA7F0",
    x"39FE881D",
    x"39FE684E",
    x"39FE4883",
    x"39FE28BC",
    x"39FE08F8",
    x"39FDE939",
    x"39FDC97E",
    x"39FDA9C7",
    x"39FD8A14",
    x"39FD6A64",
    x"39FD4AB9",
    x"39FD2B12",
    x"39FD0B6E",
    x"39FCEBCF",
    x"39FCCC33",
    x"39FCAC9C",
    x"39FC8D08",
    x"39FC6D79",
    x"39FC4DED",
    x"39FC2E65",
    x"39FC0EE1",
    x"39FBEF61",
    x"39FBCFE5",
    x"39FBB06D",
    x"39FB90F9",
    x"39FB7189",
    x"39FB521D",
    x"39FB32B5",
    x"39FB1350",
    x"39FAF3F0",
    x"39FAD493",
    x"39FAB53B",
    x"39FA95E6",
    x"39FA7695",
    x"39FA5748",
    x"39FA37FF",
    x"39FA18BA",
    x"39F9F979",
    x"39F9DA3C",
    x"39F9BB03",
    x"39F99BCD",
    x"39F97C9C",
    x"39F95D6E",
    x"39F93E44",
    x"39F91F1E",
    x"39F8FFFC",
    x"39F8E0DE",
    x"39F8C1C4",
    x"39F8A2AE",
    x"39F8839C",
    x"39F8648D",
    x"39F84582",
    x"39F8267C",
    x"39F80779",
    x"39F7E87A",
    x"39F7C97F",
    x"39F7AA87",
    x"39F78B94",
    x"39F76CA5",
    x"39F74DB9",
    x"39F72ED1",
    x"39F70FED",
    x"39F6F10D",
    x"39F6D231",
    x"39F6B359",
    x"39F69484",
    x"39F675B3",
    x"39F656E7",
    x"39F6381E",
    x"39F61959",
    x"39F5FA97",
    x"39F5DBDA",
    x"39F5BD20",
    x"39F59E6B",
    x"39F57FB9",
    x"39F5610B",
    x"39F54261",
    x"39F523BA",
    x"39F50518",
    x"39F4E679",
    x"39F4C7DE",
    x"39F4A947",
    x"39F48AB4",
    x"39F46C24",
    x"39F44D99",
    x"39F42F11",
    x"39F4108D",
    x"39F3F20D",
    x"39F3D390",
    x"39F3B518",
    x"39F396A3",
    x"39F37832",
    x"39F359C5",
    x"39F33B5C",
    x"39F31CF6",
    x"39F2FE95",
    x"39F2E037",
    x"39F2C1DC",
    x"39F2A386",
    x"39F28534",
    x"39F266E5",
    x"39F2489A",
    x"39F22A53",
    x"39F20C0F",
    x"39F1EDD0",
    x"39F1CF94",
    x"39F1B15C",
    x"39F19327",
    x"39F174F7",
    x"39F156CA",
    x"39F138A1",
    x"39F11A7C",
    x"39F0FC5B",
    x"39F0DE3D",
    x"39F0C023",
    x"39F0A20D",
    x"39F083FB",
    x"39F065EC",
    x"39F047E1",
    x"39F029DA",
    x"39F00BD7",
    x"39EFEDD7",
    x"39EFCFDB",
    x"39EFB1E3",
    x"39EF93EF",
    x"39EF75FE",
    x"39EF5811",
    x"39EF3A28",
    x"39EF1C43",
    x"39EEFE61",
    x"39EEE083",
    x"39EEC2A9",
    x"39EEA4D2",
    x"39EE8700",
    x"39EE6931",
    x"39EE4B65",
    x"39EE2D9E",
    x"39EE0FDA",
    x"39EDF21A",
    x"39EDD45D",
    x"39EDB6A5",
    x"39ED98F0",
    x"39ED7B3F",
    x"39ED5D91",
    x"39ED3FE7",
    x"39ED2241",
    x"39ED049F",
    x"39ECE700",
    x"39ECC965",
    x"39ECABCD",
    x"39EC8E3A",
    x"39EC70AA",
    x"39EC531E",
    x"39EC3595",
    x"39EC1810",
    x"39EBFA8F",
    x"39EBDD12",
    x"39EBBF98",
    x"39EBA222",
    x"39EB84AF",
    x"39EB6741",
    x"39EB49D6",
    x"39EB2C6E",
    x"39EB0F0A",
    x"39EAF1AA",
    x"39EAD44E",
    x"39EAB6F5",
    x"39EA99A0",
    x"39EA7C4F",
    x"39EA5F01",
    x"39EA41B7",
    x"39EA2471",
    x"39EA072E",
    x"39E9E9EF",
    x"39E9CCB4",
    x"39E9AF7C",
    x"39E99248",
    x"39E97517",
    x"39E957EA",
    x"39E93AC1",
    x"39E91D9C",
    x"39E9007A",
    x"39E8E35C",
    x"39E8C641",
    x"39E8A92A",
    x"39E88C17",
    x"39E86F07",
    x"39E851FB",
    x"39E834F2",
    x"39E817EE",
    x"39E7FAED",
    x"39E7DDEF",
    x"39E7C0F5",
    x"39E7A3FF",
    x"39E7870C",
    x"39E76A1D",
    x"39E74D31",
    x"39E7304A",
    x"39E71365",
    x"39E6F685",
    x"39E6D9A8",
    x"39E6BCCE",
    x"39E69FF9",
    x"39E68326",
    x"39E66658",
    x"39E6498D",
    x"39E62CC5",
    x"39E61002",
    x"39E5F341",
    x"39E5D685",
    x"39E5B9CC",
    x"39E59D16",
    x"39E58065",
    x"39E563B6",
    x"39E5470C",
    x"39E52A64",
    x"39E50DC1",
    x"39E4F121",
    x"39E4D485",
    x"39E4B7EC",
    x"39E49B57",
    x"39E47EC5",
    x"39E46237",
    x"39E445AD",
    x"39E42926",
    x"39E40CA2",
    x"39E3F022",
    x"39E3D3A6",
    x"39E3B72E",
    x"39E39AB8",
    x"39E37E47",
    x"39E361D9",
    x"39E3456E",
    x"39E32907",
    x"39E30CA4",
    x"39E2F044",
    x"39E2D3E8",
    x"39E2B78F",
    x"39E29B3A",
    x"39E27EE9",
    x"39E2629A",
    x"39E24650",
    x"39E22A09",
    x"39E20DC5",
    x"39E1F185",
    x"39E1D549",
    x"39E1B910",
    x"39E19CDB",
    x"39E180A9",
    x"39E1647B",
    x"39E14850",
    x"39E12C28",
    x"39E11005",
    x"39E0F3E4",
    x"39E0D7C8",
    x"39E0BBAF",
    x"39E09F99",
    x"39E08387",
    x"39E06778",
    x"39E04B6D",
    x"39E02F65",
    x"39E01361",
    x"39DFF760",
    x"39DFDB63",
    x"39DFBF69",
    x"39DFA373",
    x"39DF8781",
    x"39DF6B91",
    x"39DF4FA6",
    x"39DF33BD",
    x"39DF17D9",
    x"39DEFBF7",
    x"39DEE01A",
    x"39DEC43F",
    x"39DEA869",
    x"39DE8C95",
    x"39DE70C6",
    x"39DE54F9",
    x"39DE3930",
    x"39DE1D6B",
    x"39DE01A9",
    x"39DDE5EA",
    x"39DDCA2F",
    x"39DDAE78",
    x"39DD92C4",
    x"39DD7713",
    x"39DD5B66",
    x"39DD3FBC",
    x"39DD2416",
    x"39DD0873",
    x"39DCECD4",
    x"39DCD138",
    x"39DCB5A0",
    x"39DC9A0B",
    x"39DC7E79",
    x"39DC62EB",
    x"39DC4760",
    x"39DC2BD9",
    x"39DC1055",
    x"39DBF4D5",
    x"39DBD958",
    x"39DBBDDF",
    x"39DBA269",
    x"39DB86F6",
    x"39DB6B87",
    x"39DB501B",
    x"39DB34B3",
    x"39DB194E",
    x"39DAFDED",
    x"39DAE28F",
    x"39DAC734",
    x"39DAABDD",
    x"39DA9089",
    x"39DA7539",
    x"39DA59EC",
    x"39DA3EA2",
    x"39DA235C",
    x"39DA0819",
    x"39D9ECDA",
    x"39D9D19E",
    x"39D9B666",
    x"39D99B31",
    x"39D97FFF",
    x"39D964D1",
    x"39D949A6",
    x"39D92E7E",
    x"39D9135A",
    x"39D8F839",
    x"39D8DD1C",
    x"39D8C202",
    x"39D8A6EC",
    x"39D88BD8",
    x"39D870C9",
    x"39D855BC",
    x"39D83AB3",
    x"39D81FAD",
    x"39D804AB",
    x"39D7E9AC",
    x"39D7CEB1",
    x"39D7B3B9",
    x"39D798C4",
    x"39D77DD2",
    x"39D762E4",
    x"39D747FA",
    x"39D72D12",
    x"39D7122E",
    x"39D6F74E",
    x"39D6DC71",
    x"39D6C197",
    x"39D6A6C0",
    x"39D68BED",
    x"39D6711D",
    x"39D65651",
    x"39D63B88",
    x"39D620C2",
    x"39D605FF",
    x"39D5EB40",
    x"39D5D085",
    x"39D5B5CC",
    x"39D59B17",
    x"39D58066",
    x"39D565B7",
    x"39D54B0C",
    x"39D53064",
    x"39D515C0",
    x"39D4FB1F",
    x"39D4E081",
    x"39D4C5E7",
    x"39D4AB50",
    x"39D490BC",
    x"39D4762C",
    x"39D45B9E",
    x"39D44115",
    x"39D4268E",
    x"39D40C0B",
    x"39D3F18B",
    x"39D3D70F",
    x"39D3BC95",
    x"39D3A21F",
    x"39D387AD",
    x"39D36D3E",
    x"39D352D2",
    x"39D33869",
    x"39D31E03",
    x"39D303A1",
    x"39D2E943",
    x"39D2CEE7",
    x"39D2B48F",
    x"39D29A3A",
    x"39D27FE8",
    x"39D2659A",
    x"39D24B4F",
    x"39D23107",
    x"39D216C3",
    x"39D1FC81",
    x"39D1E243",
    x"39D1C809",
    x"39D1ADD1",
    x"39D1939D",
    x"39D1796D",
    x"39D15F3F",
    x"39D14515",
    x"39D12AEE",
    x"39D110CA",
    x"39D0F6AA",
    x"39D0DC8C",
    x"39D0C272",
    x"39D0A85C",
    x"39D08E48",
    x"39D07438",
    x"39D05A2B",
    x"39D04022",
    x"39D0261B",
    x"39D00C18",
    x"39CFF218",
    x"39CFD81C",
    x"39CFBE22",
    x"39CFA42C",
    x"39CF8A39",
    x"39CF7049",
    x"39CF565D",
    x"39CF3C74",
    x"39CF228E",
    x"39CF08AB",
    x"39CEEECC",
    x"39CED4F0",
    x"39CEBB17",
    x"39CEA141",
    x"39CE876E",
    x"39CE6D9F",
    x"39CE53D3",
    x"39CE3A0A",
    x"39CE2044",
    x"39CE0682",
    x"39CDECC3",
    x"39CDD307",
    x"39CDB94E",
    x"39CD9F98",
    x"39CD85E6",
    x"39CD6C37",
    x"39CD528B",
    x"39CD38E2",
    x"39CD1F3D",
    x"39CD059A",
    x"39CCEBFB",
    x"39CCD25F",
    x"39CCB8C7",
    x"39CC9F31",
    x"39CC859F",
    x"39CC6C10",
    x"39CC5284",
    x"39CC38FB",
    x"39CC1F76",
    x"39CC05F3",
    x"39CBEC74",
    x"39CBD2F8",
    x"39CBB97F",
    x"39CBA00A",
    x"39CB8697",
    x"39CB6D28",
    x"39CB53BC",
    x"39CB3A53",
    x"39CB20EE",
    x"39CB078B",
    x"39CAEE2C",
    x"39CAD4CF",
    x"39CABB76",
    x"39CAA221",
    x"39CA88CE",
    x"39CA6F7E",
    x"39CA5632",
    x"39CA3CE9",
    x"39CA23A3",
    x"39CA0A60",
    x"39C9F120",
    x"39C9D7E4",
    x"39C9BEAA",
    x"39C9A574",
    x"39C98C41",
    x"39C97311",
    x"39C959E4",
    x"39C940BA",
    x"39C92794",
    x"39C90E71",
    x"39C8F550",
    x"39C8DC33",
    x"39C8C319",
    x"39C8AA02",
    x"39C890EF",
    x"39C877DE",
    x"39C85ED1",
    x"39C845C7",
    x"39C82CBF",
    x"39C813BB",
    x"39C7FABA",
    x"39C7E1BD",
    x"39C7C8C2",
    x"39C7AFCA",
    x"39C796D6",
    x"39C77DE5",
    x"39C764F7",
    x"39C74C0C",
    x"39C73324",
    x"39C71A3F",
    x"39C7015D",
    x"39C6E87E",
    x"39C6CFA3",
    x"39C6B6CB",
    x"39C69DF5",
    x"39C68523",
    x"39C66C54",
    x"39C65388",
    x"39C63ABF",
    x"39C621F9",
    x"39C60937",
    x"39C5F077",
    x"39C5D7BA",
    x"39C5BF01",
    x"39C5A64B",
    x"39C58D97",
    x"39C574E7",
    x"39C55C3A",
    x"39C54390",
    x"39C52AE9",
    x"39C51245",
    x"39C4F9A5",
    x"39C4E107",
    x"39C4C86C",
    x"39C4AFD5",
    x"39C49741",
    x"39C47EAF",
    x"39C46621",
    x"39C44D96",
    x"39C4350D",
    x"39C41C88",
    x"39C40406",
    x"39C3EB87",
    x"39C3D30B",
    x"39C3BA93",
    x"39C3A21D",
    x"39C389AA",
    x"39C3713A",
    x"39C358CE",
    x"39C34064",
    x"39C327FE",
    x"39C30F9A",
    x"39C2F73A",
    x"39C2DEDC",
    x"39C2C682",
    x"39C2AE2B",
    x"39C295D7",
    x"39C27D85",
    x"39C26537",
    x"39C24CEC",
    x"39C234A4",
    x"39C21C5F",
    x"39C2041D",
    x"39C1EBDE",
    x"39C1D3A2",
    x"39C1BB69",
    x"39C1A333",
    x"39C18B00",
    x"39C172D0",
    x"39C15AA3",
    x"39C1427A",
    x"39C12A53",
    x"39C1122F",
    x"39C0FA0E",
    x"39C0E1F0",
    x"39C0C9D6",
    x"39C0B1BE",
    x"39C099A9",
    x"39C08198",
    x"39C06989",
    x"39C0517D",
    x"39C03975",
    x"39C0216F",
    x"39C0096C",
    x"39BFF16C",
    x"39BFD970",
    x"39BFC176",
    x"39BFA97F",
    x"39BF918C",
    x"39BF799B",
    x"39BF61AD",
    x"39BF49C3",
    x"39BF31DB",
    x"39BF19F6",
    x"39BF0214",
    x"39BEEA36",
    x"39BED25A",
    x"39BEBA81",
    x"39BEA2AB",
    x"39BE8AD8",
    x"39BE7309",
    x"39BE5B3C",
    x"39BE4372",
    x"39BE2BAB",
    x"39BE13E7",
    x"39BDFC26",
    x"39BDE468",
    x"39BDCCAD",
    x"39BDB4F5",
    x"39BD9D3F",
    x"39BD858D",
    x"39BD6DDE",
    x"39BD5632",
    x"39BD3E89",
    x"39BD26E2",
    x"39BD0F3F",
    x"39BCF79E",
    x"39BCE001",
    x"39BCC866",
    x"39BCB0CF",
    x"39BC993A",
    x"39BC81A8",
    x"39BC6A1A",
    x"39BC528E",
    x"39BC3B05",
    x"39BC237F",
    x"39BC0BFC",
    x"39BBF47C",
    x"39BBDCFF",
    x"39BBC585",
    x"39BBAE0E",
    x"39BB9699",
    x"39BB7F28",
    x"39BB67BA",
    x"39BB504E",
    x"39BB38E6",
    x"39BB2180",
    x"39BB0A1D",
    x"39BAF2BD",
    x"39BADB61",
    x"39BAC407",
    x"39BAACB0",
    x"39BA955B",
    x"39BA7E0A",
    x"39BA66BC",
    x"39BA4F70",
    x"39BA3828",
    x"39BA20E2",
    x"39BA09A0",
    x"39B9F260",
    x"39B9DB23",
    x"39B9C3E9",
    x"39B9ACB2",
    x"39B9957E",
    x"39B97E4D",
    x"39B9671F",
    x"39B94FF3",
    x"39B938CB",
    x"39B921A5",
    x"39B90A82",
    x"39B8F362",
    x"39B8DC45",
    x"39B8C52B",
    x"39B8AE14",
    x"39B89700",
    x"39B87FEE",
    x"39B868E0",
    x"39B851D4",
    x"39B83ACB",
    x"39B823C5",
    x"39B80CC2",
    x"39B7F5C2",
    x"39B7DEC5",
    x"39B7C7CA",
    x"39B7B0D3",
    x"39B799DE",
    x"39B782EC",
    x"39B76BFD",
    x"39B75511",
    x"39B73E28",
    x"39B72742",
    x"39B7105E",
    x"39B6F97E",
    x"39B6E2A0",
    x"39B6CBC5",
    x"39B6B4ED",
    x"39B69E18",
    x"39B68746",
    x"39B67076",
    x"39B659A9",
    x"39B642E0",
    x"39B62C19",
    x"39B61555",
    x"39B5FE93",
    x"39B5E7D5",
    x"39B5D119",
    x"39B5BA61",
    x"39B5A3AB",
    x"39B58CF8",
    x"39B57648",
    x"39B55F9A",
    x"39B548F0",
    x"39B53248",
    x"39B51BA3",
    x"39B50501",
    x"39B4EE62",
    x"39B4D7C5",
    x"39B4C12C",
    x"39B4AA95",
    x"39B49401",
    x"39B47D70",
    x"39B466E2",
    x"39B45056",
    x"39B439CE",
    x"39B42348",
    x"39B40CC5",
    x"39B3F645",
    x"39B3DFC7",
    x"39B3C94D",
    x"39B3B2D5",
    x"39B39C60",
    x"39B385EE",
    x"39B36F7F",
    x"39B35912",
    x"39B342A8",
    x"39B32C41",
    x"39B315DD",
    x"39B2FF7C",
    x"39B2E91D",
    x"39B2D2C2",
    x"39B2BC69",
    x"39B2A613",
    x"39B28FBF",
    x"39B2796F",
    x"39B26321",
    x"39B24CD6",
    x"39B2368E",
    x"39B22048",
    x"39B20A06",
    x"39B1F3C6",
    x"39B1DD89",
    x"39B1C74E",
    x"39B1B117",
    x"39B19AE2",
    x"39B184B0",
    x"39B16E81",
    x"39B15855",
    x"39B1422B",
    x"39B12C04",
    x"39B115E0",
    x"39B0FFBF",
    x"39B0E9A0",
    x"39B0D384",
    x"39B0BD6B",
    x"39B0A755",
    x"39B09141",
    x"39B07B30",
    x"39B06522",
    x"39B04F17",
    x"39B0390F",
    x"39B02309",
    x"39B00D06",
    x"39AFF706",
    x"39AFE108",
    x"39AFCB0D",
    x"39AFB515",
    x"39AF9F20",
    x"39AF892E",
    x"39AF733E",
    x"39AF5D51",
    x"39AF4766",
    x"39AF317F",
    x"39AF1B9A",
    x"39AF05B8",
    x"39AEEFD9",
    x"39AED9FC",
    x"39AEC422",
    x"39AEAE4B",
    x"39AE9877",
    x"39AE82A5",
    x"39AE6CD6",
    x"39AE570A",
    x"39AE4140",
    x"39AE2B79",
    x"39AE15B5",
    x"39ADFFF4",
    x"39ADEA35",
    x"39ADD479",
    x"39ADBEC0",
    x"39ADA90A",
    x"39AD9356",
    x"39AD7DA5",
    x"39AD67F7",
    x"39AD524B",
    x"39AD3CA2",
    x"39AD26FC",
    x"39AD1158",
    x"39ACFBB7",
    x"39ACE619",
    x"39ACD07E",
    x"39ACBAE5",
    x"39ACA54F",
    x"39AC8FBC",
    x"39AC7A2B",
    x"39AC649D",
    x"39AC4F12",
    x"39AC398A",
    x"39AC2404",
    x"39AC0E81",
    x"39ABF900",
    x"39ABE382",
    x"39ABCE07",
    x"39ABB88F",
    x"39ABA319",
    x"39AB8DA6",
    x"39AB7836",
    x"39AB62C8",
    x"39AB4D5D",
    x"39AB37F5",
    x"39AB228F",
    x"39AB0D2C",
    x"39AAF7CC",
    x"39AAE26E",
    x"39AACD13",
    x"39AAB7BB",
    x"39AAA265",
    x"39AA8D12",
    x"39AA77C2",
    x"39AA6274",
    x"39AA4D29",
    x"39AA37E1",
    x"39AA229B",
    x"39AA0D58",
    x"39A9F818",
    x"39A9E2DA",
    x"39A9CD9F",
    x"39A9B867",
    x"39A9A331",
    x"39A98DFE",
    x"39A978CE",
    x"39A963A0",
    x"39A94E75",
    x"39A9394C",
    x"39A92426",
    x"39A90F03",
    x"39A8F9E3",
    x"39A8E4C5",
    x"39A8CFA9",
    x"39A8BA91",
    x"39A8A57B",
    x"39A89067",
    x"39A87B57",
    x"39A86649",
    x"39A8513D",
    x"39A83C34",
    x"39A8272E",
    x"39A8122A",
    x"39A7FD2A",
    x"39A7E82B",
    x"39A7D32F",
    x"39A7BE36",
    x"39A7A940",
    x"39A7944C",
    x"39A77F5B",
    x"39A76A6C",
    x"39A75580",
    x"39A74097",
    x"39A72BB0",
    x"39A716CC",
    x"39A701EA",
    x"39A6ED0B",
    x"39A6D82F",
    x"39A6C355",
    x"39A6AE7E",
    x"39A699AA",
    x"39A684D8",
    x"39A67009",
    x"39A65B3C",
    x"39A64672",
    x"39A631AA",
    x"39A61CE5",
    x"39A60823",
    x"39A5F363",
    x"39A5DEA6",
    x"39A5C9EC",
    x"39A5B534",
    x"39A5A07E",
    x"39A58BCC",
    x"39A5771B",
    x"39A5626E",
    x"39A54DC3",
    x"39A5391A",
    x"39A52475",
    x"39A50FD1",
    x"39A4FB31",
    x"39A4E692",
    x"39A4D1F7",
    x"39A4BD5E",
    x"39A4A8C8",
    x"39A49434",
    x"39A47FA3",
    x"39A46B14",
    x"39A45688",
    x"39A441FE",
    x"39A42D77",
    x"39A418F3",
    x"39A40471",
    x"39A3EFF2",
    x"39A3DB75",
    x"39A3C6FB",
    x"39A3B283",
    x"39A39E0E",
    x"39A3899C",
    x"39A3752C",
    x"39A360BE",
    x"39A34C54",
    x"39A337EB",
    x"39A32386",
    x"39A30F23",
    x"39A2FAC2",
    x"39A2E664",
    x"39A2D208",
    x"39A2BDAF",
    x"39A2A959",
    x"39A29505",
    x"39A280B4",
    x"39A26C65",
    x"39A25819",
    x"39A243CF",
    x"39A22F88",
    x"39A21B43",
    x"39A20701",
    x"39A1F2C1",
    x"39A1DE84",
    x"39A1CA4A",
    x"39A1B611",
    x"39A1A1DC",
    x"39A18DA9",
    x"39A17979",
    x"39A1654B",
    x"39A1511F",
    x"39A13CF6",
    x"39A128D0",
    x"39A114AC",
    x"39A1008B",
    x"39A0EC6C",
    x"39A0D850",
    x"39A0C436",
    x"39A0B01F",
    x"39A09C0A",
    x"39A087F8",
    x"39A073E8",
    x"39A05FDB",
    x"39A04BD0",
    x"39A037C8",
    x"39A023C2",
    x"39A00FBF",
    x"399FFBBE",
    x"399FE7C0",
    x"399FD3C4",
    x"399FBFCB",
    x"399FABD4",
    x"399F97E0",
    x"399F83EE",
    x"399F6FFF",
    x"399F5C12",
    x"399F4828",
    x"399F3440",
    x"399F205B",
    x"399F0C78",
    x"399EF898",
    x"399EE4BA",
    x"399ED0DF",
    x"399EBD06",
    x"399EA92F",
    x"399E955B",
    x"399E818A",
    x"399E6DBB",
    x"399E59EF",
    x"399E4625",
    x"399E325D",
    x"399E1E98",
    x"399E0AD5",
    x"399DF715",
    x"399DE358",
    x"399DCF9C",
    x"399DBBE4",
    x"399DA82D",
    x"399D947A",
    x"399D80C8",
    x"399D6D19",
    x"399D596D",
    x"399D45C3",
    x"399D321C",
    x"399D1E77",
    x"399D0AD4",
    x"399CF734",
    x"399CE396",
    x"399CCFFB",
    x"399CBC62",
    x"399CA8CC",
    x"399C9538",
    x"399C81A7",
    x"399C6E18",
    x"399C5A8B",
    x"399C4701",
    x"399C3379",
    x"399C1FF4",
    x"399C0C71",
    x"399BF8F1",
    x"399BE573",
    x"399BD1F8",
    x"399BBE7F",
    x"399BAB08",
    x"399B9794",
    x"399B8422",
    x"399B70B3",
    x"399B5D46",
    x"399B49DB",
    x"399B3673",
    x"399B230E",
    x"399B0FAB",
    x"399AFC4A",
    x"399AE8EC",
    x"399AD590",
    x"399AC236",
    x"399AAEDF",
    x"399A9B8B",
    x"399A8838",
    x"399A74E8",
    x"399A619B",
    x"399A4E50",
    x"399A3B07",
    x"399A27C1",
    x"399A147E",
    x"399A013C",
    x"3999EDFD",
    x"3999DAC1",
    x"3999C787",
    x"3999B44F",
    x"3999A119",
    x"39998DE7",
    x"39997AB6",
    x"39996788",
    x"3999545C",
    x"39994133",
    x"39992E0C",
    x"39991AE7",
    x"399907C5",
    x"3998F4A5",
    x"3998E188",
    x"3998CE6D",
    x"3998BB54",
    x"3998A83E",
    x"3998952A",
    x"39988219",
    x"39986F0A",
    x"39985BFD",
    x"399848F3",
    x"399835EB",
    x"399822E5",
    x"39980FE2",
    x"3997FCE1",
    x"3997E9E3",
    x"3997D6E7",
    x"3997C3ED",
    x"3997B0F6",
    x"39979E01",
    x"39978B0E",
    x"3997781E",
    x"39976530",
    x"39975245",
    x"39973F5C",
    x"39972C75",
    x"39971991",
    x"399706AF",
    x"3996F3CF",
    x"3996E0F2",
    x"3996CE17",
    x"3996BB3E",
    x"3996A868",
    x"39969594",
    x"399682C3",
    x"39966FF3",
    x"39965D27",
    x"39964A5C",
    x"39963794",
    x"399624CE",
    x"3996120B",
    x"3995FF4A",
    x"3995EC8B",
    x"3995D9CF",
    x"3995C714",
    x"3995B45D",
    x"3995A1A7",
    x"39958EF4",
    x"39957C44",
    x"39956995",
    x"399556E9",
    x"39954440",
    x"39953198",
    x"39951EF3",
    x"39950C50",
    x"3994F9B0",
    x"3994E712",
    x"3994D476",
    x"3994C1DD",
    x"3994AF46",
    x"39949CB1",
    x"39948A1F",
    x"3994778F",
    x"39946501",
    x"39945275",
    x"39943FEC",
    x"39942D65",
    x"39941AE1",
    x"3994085F",
    x"3993F5DF",
    x"3993E361",
    x"3993D0E6",
    x"3993BE6D",
    x"3993ABF6",
    x"39939982",
    x"39938710",
    x"399374A0",
    x"39936233",
    x"39934FC8",
    x"39933D5F",
    x"39932AF8",
    x"39931894",
    x"39930632",
    x"3992F3D2",
    x"3992E175",
    x"3992CF1A",
    x"3992BCC1",
    x"3992AA6B",
    x"39929817",
    x"399285C5",
    x"39927375",
    x"39926128",
    x"39924EDD",
    x"39923C94",
    x"39922A4E",
    x"3992180A",
    x"399205C8",
    x"3991F388",
    x"3991E14B",
    x"3991CF10",
    x"3991BCD7",
    x"3991AAA1",
    x"3991986D",
    x"3991863B",
    x"3991740B",
    x"399161DE",
    x"39914FB3",
    x"39913D8A",
    x"39912B63",
    x"3991193F",
    x"3991071D",
    x"3990F4FD",
    x"3990E2E0",
    x"3990D0C4",
    x"3990BEAB",
    x"3990AC95",
    x"39909A80",
    x"3990886E",
    x"3990765E",
    x"39906450",
    x"39905245",
    x"3990403C",
    x"39902E35",
    x"39901C30",
    x"39900A2E",
    x"398FF82E",
    x"398FE630",
    x"398FD434",
    x"398FC23B",
    x"398FB044",
    x"398F9E4F",
    x"398F8C5C",
    x"398F7A6C",
    x"398F687E",
    x"398F5692",
    x"398F44A8",
    x"398F32C0",
    x"398F20DB",
    x"398F0EF8",
    x"398EFD17",
    x"398EEB39",
    x"398ED95D",
    x"398EC783",
    x"398EB5AB",
    x"398EA3D5",
    x"398E9202",
    x"398E8031",
    x"398E6E62",
    x"398E5C95",
    x"398E4ACB",
    x"398E3902",
    x"398E273C",
    x"398E1579",
    x"398E03B7",
    x"398DF1F8",
    x"398DE03B",
    x"398DCE80",
    x"398DBCC7",
    x"398DAB10",
    x"398D995C",
    x"398D87AA",
    x"398D75FA",
    x"398D644D",
    x"398D52A1",
    x"398D40F8",
    x"398D2F51",
    x"398D1DAC",
    x"398D0C09",
    x"398CFA69",
    x"398CE8CB",
    x"398CD72F",
    x"398CC595",
    x"398CB3FD",
    x"398CA268",
    x"398C90D5",
    x"398C7F44",
    x"398C6DB5",
    x"398C5C28",
    x"398C4A9E",
    x"398C3916",
    x"398C2790",
    x"398C160C",
    x"398C048A",
    x"398BF30B",
    x"398BE18D",
    x"398BD012",
    x"398BBE99",
    x"398BAD23",
    x"398B9BAE",
    x"398B8A3C",
    x"398B78CC",
    x"398B675E",
    x"398B55F2",
    x"398B4488",
    x"398B3321",
    x"398B21BB",
    x"398B1058",
    x"398AFEF7",
    x"398AED98",
    x"398ADC3C",
    x"398ACAE1",
    x"398AB989",
    x"398AA833",
    x"398A96DF",
    x"398A858D",
    x"398A743E",
    x"398A62F0",
    x"398A51A5",
    x"398A405C",
    x"398A2F15",
    x"398A1DD0",
    x"398A0C8D",
    x"3989FB4D",
    x"3989EA0F",
    x"3989D8D2",
    x"3989C798",
    x"3989B660",
    x"3989A52B",
    x"398993F7",
    x"398982C6",
    x"39897197",
    x"39896069",
    x"39894F3E",
    x"39893E16",
    x"39892CEF",
    x"39891BCA",
    x"39890AA8",
    x"3988F988",
    x"3988E86A",
    x"3988D74E",
    x"3988C634",
    x"3988B51C",
    x"3988A406",
    x"398892F3",
    x"398881E2",
    x"398870D3",
    x"39885FC6",
    x"39884EBB",
    x"39883DB2",
    x"39882CAB",
    x"39881BA7",
    x"39880AA4",
    x"3987F9A4",
    x"3987E8A6",
    x"3987D7AA",
    x"3987C6B0",
    x"3987B5B8",
    x"3987A4C3",
    x"398793CF",
    x"398782DE",
    x"398771EE",
    x"39876101",
    x"39875016",
    x"39873F2D",
    x"39872E46",
    x"39871D61",
    x"39870C7F",
    x"3986FB9E",
    x"3986EAC0",
    x"3986D9E4",
    x"3986C909",
    x"3986B831",
    x"3986A75B",
    x"39869688",
    x"398685B6",
    x"398674E6",
    x"39866419",
    x"3986534D",
    x"39864284",
    x"398631BC",
    x"398620F7",
    x"39861034",
    x"3985FF73",
    x"3985EEB4",
    x"3985DDF8",
    x"3985CD3D",
    x"3985BC84",
    x"3985ABCE",
    x"39859B19",
    x"39858A67",
    x"398579B7",
    x"39856909",
    x"3985585C",
    x"398547B2",
    x"3985370B",
    x"39852665",
    x"398515C1",
    x"3985051F",
    x"3984F480",
    x"3984E3E2",
    x"3984D347",
    x"3984C2AD",
    x"3984B216",
    x"3984A181",
    x"398490EE",
    x"3984805D",
    x"39846FCE",
    x"39845F41",
    x"39844EB6",
    x"39843E2D",
    x"39842DA6",
    x"39841D22",
    x"39840C9F",
    x"3983FC1E",
    x"3983EBA0",
    x"3983DB23",
    x"3983CAA9",
    x"3983BA31",
    x"3983A9BB",
    x"39839946",
    x"398388D4",
    x"39837864",
    x"398367F6",
    x"3983578A",
    x"39834720",
    x"398336B8",
    x"39832653",
    x"398315EF",
    x"3983058D",
    x"3982F52D",
    x"3982E4D0",
    x"3982D474",
    x"3982C41B",
    x"3982B3C3",
    x"3982A36E",
    x"3982931A",
    x"398282C9",
    x"3982727A",
    x"3982622C",
    x"398251E1",
    x"39824198",
    x"39823151",
    x"3982210C",
    x"398210C8",
    x"39820087",
    x"3981F048",
    x"3981E00B",
    x"3981CFD0",
    x"3981BF97",
    x"3981AF60",
    x"39819F2B",
    x"39818EF9",
    x"39817EC8",
    x"39816E99",
    x"39815E6C",
    x"39814E41",
    x"39813E19",
    x"39812DF2",
    x"39811DCD",
    x"39810DAA",
    x"3980FD8A",
    x"3980ED6B",
    x"3980DD4E",
    x"3980CD34",
    x"3980BD1B",
    x"3980AD04",
    x"39809CF0",
    x"39808CDD",
    x"39807CCC",
    x"39806CBE",
    x"39805CB1",
    x"39804CA7",
    x"39803C9E",
    x"39802C98",
    x"39801C93",
    x"39800C90",
    x"397FF920",
    x"397FD923",
    x"397FB929",
    x"397F9934",
    x"397F7943",
    x"397F5956",
    x"397F396D",
    x"397F1988",
    x"397EF9A6",
    x"397ED9C9",
    x"397EB9F0",
    x"397E9A1B",
    x"397E7A49",
    x"397E5A7C",
    x"397E3AB3",
    x"397E1AED",
    x"397DFB2C",
    x"397DDB6F",
    x"397DBBB5",
    x"397D9C00",
    x"397D7C4E",
    x"397D5CA1",
    x"397D3CF7",
    x"397D1D51",
    x"397CFDB0",
    x"397CDE12",
    x"397CBE78",
    x"397C9EE2",
    x"397C7F50",
    x"397C5FC3",
    x"397C4039",
    x"397C20B2",
    x"397C0130",
    x"397BE1B2",
    x"397BC238",
    x"397BA2C2",
    x"397B834F",
    x"397B63E1",
    x"397B4476",
    x"397B2510",
    x"397B05AD",
    x"397AE64E",
    x"397AC6F3",
    x"397AA79D",
    x"397A884A",
    x"397A68FA",
    x"397A49AF",
    x"397A2A68",
    x"397A0B25",
    x"3979EBE5",
    x"3979CCAA",
    x"3979AD72",
    x"39798E3E",
    x"39796F0F",
    x"39794FE3",
    x"397930BB",
    x"39791196",
    x"3978F276",
    x"3978D35A",
    x"3978B441",
    x"3978952D",
    x"3978761C",
    x"3978570F",
    x"39783806",
    x"39781901",
    x"3977FA00",
    x"3977DB03",
    x"3977BC09",
    x"39779D14",
    x"39777E22",
    x"39775F34",
    x"3977404A",
    x"39772164",
    x"39770282",
    x"3976E3A3",
    x"3976C4C9",
    x"3976A5F2",
    x"3976871F",
    x"39766850",
    x"39764985",
    x"39762ABE",
    x"39760BFB",
    x"3975ED3B",
    x"3975CE7F",
    x"3975AFC7",
    x"39759113",
    x"39757263",
    x"397553B7",
    x"3975350E",
    x"3975166A",
    x"3974F7C9",
    x"3974D92C",
    x"3974BA92",
    x"39749BFD",
    x"39747D6B",
    x"39745EDE",
    x"39744054",
    x"397421CE",
    x"3974034B",
    x"3973E4CD",
    x"3973C652",
    x"3973A7DB",
    x"39738968",
    x"39736AF9",
    x"39734C8D",
    x"39732E26",
    x"39730FC2",
    x"3972F162",
    x"3972D305",
    x"3972B4AD",
    x"39729658",
    x"39727807",
    x"397259BA",
    x"39723B71",
    x"39721D2B",
    x"3971FEEA",
    x"3971E0AC",
    x"3971C271",
    x"3971A43B",
    x"39718608",
    x"397167DA",
    x"397149AE",
    x"39712B87",
    x"39710D64",
    x"3970EF44",
    x"3970D128",
    x"3970B30F",
    x"397094FB",
    x"397076EA",
    x"397058DD",
    x"39703AD4",
    x"39701CCF",
    x"396FFECD",
    x"396FE0CF",
    x"396FC2D5",
    x"396FA4DE",
    x"396F86EB",
    x"396F68FC",
    x"396F4B11",
    x"396F2D2A",
    x"396F0F46",
    x"396EF166",
    x"396ED38A",
    x"396EB5B1",
    x"396E97DC",
    x"396E7A0B",
    x"396E5C3E",
    x"396E3E74",
    x"396E20AE",
    x"396E02EC",
    x"396DE52D",
    x"396DC772",
    x"396DA9BB",
    x"396D8C08",
    x"396D6E58",
    x"396D50AC",
    x"396D3304",
    x"396D1560",
    x"396CF7BF",
    x"396CDA22",
    x"396CBC88",
    x"396C9EF3",
    x"396C8161",
    x"396C63D2",
    x"396C4648",
    x"396C28C1",
    x"396C0B3D",
    x"396BEDBE",
    x"396BD042",
    x"396BB2CA",
    x"396B9555",
    x"396B77E4",
    x"396B5A77",
    x"396B3D0E",
    x"396B1FA8",
    x"396B0246",
    x"396AE4E7",
    x"396AC78D",
    x"396AAA36",
    x"396A8CE2",
    x"396A6F92",
    x"396A5246",
    x"396A34FE",
    x"396A17B9",
    x"3969FA78",
    x"3969DD3A",
    x"3969C001",
    x"3969A2CA",
    x"39698598",
    x"39696869",
    x"39694B3E",
    x"39692E16",
    x"396910F2",
    x"3968F3D2",
    x"3968D6B5",
    x"3968B99C",
    x"39689C87",
    x"39687F75",
    x"39686267",
    x"3968455D",
    x"39682856",
    x"39680B52",
    x"3967EE53",
    x"3967D157",
    x"3967B45F",
    x"3967976A",
    x"39677A79",
    x"39675D8B",
    x"396740A1",
    x"396723BB",
    x"396706D8",
    x"3966E9F9",
    x"3966CD1E",
    x"3966B046",
    x"39669372",
    x"396676A1",
    x"396659D4",
    x"39663D0B",
    x"39662045",
    x"39660383",
    x"3965E6C4",
    x"3965CA09",
    x"3965AD51",
    x"3965909E",
    x"396573ED",
    x"39655741",
    x"39653A97",
    x"39651DF2",
    x"39650150",
    x"3964E4B2",
    x"3964C817",
    x"3964AB80",
    x"39648EEC",
    x"3964725C",
    x"396455CF",
    x"39643946",
    x"39641CC1",
    x"3964003F",
    x"3963E3C1",
    x"3963C746",
    x"3963AACF",
    x"39638E5C",
    x"396371EC",
    x"3963557F",
    x"39633916",
    x"39631CB1",
    x"3963004F",
    x"3962E3F1",
    x"3962C796",
    x"3962AB3F",
    x"39628EEB",
    x"3962729B",
    x"3962564F",
    x"39623A06",
    x"39621DC0",
    x"3962017E",
    x"3961E540",
    x"3961C905",
    x"3961ACCD",
    x"3961909A",
    x"39617469",
    x"3961583D",
    x"39613C13",
    x"39611FED",
    x"396103CB",
    x"3960E7AD",
    x"3960CB91",
    x"3960AF7A",
    x"39609365",
    x"39607755",
    x"39605B48",
    x"39603F3E",
    x"39602338",
    x"39600735",
    x"395FEB36",
    x"395FCF3A",
    x"395FB342",
    x"395F974E",
    x"395F7B5C",
    x"395F5F6F",
    x"395F4385",
    x"395F279E",
    x"395F0BBB",
    x"395EEFDB",
    x"395ED3FF",
    x"395EB826",
    x"395E9C51",
    x"395E807F",
    x"395E64B0",
    x"395E48E6",
    x"395E2D1E",
    x"395E115A",
    x"395DF59A",
    x"395DD9DD",
    x"395DBE23",
    x"395DA26D",
    x"395D86BB",
    x"395D6B0C",
    x"395D4F60",
    x"395D33B8",
    x"395D1813",
    x"395CFC72",
    x"395CE0D4",
    x"395CC53A",
    x"395CA9A3",
    x"395C8E0F",
    x"395C727F",
    x"395C56F3",
    x"395C3B69",
    x"395C1FE4",
    x"395C0462",
    x"395BE8E3",
    x"395BCD67",
    x"395BB1EF",
    x"395B967B",
    x"395B7B0A",
    x"395B5F9C",
    x"395B4432",
    x"395B28CB",
    x"395B0D68",
    x"395AF208",
    x"395AD6AB",
    x"395ABB52",
    x"395A9FFC",
    x"395A84AA",
    x"395A695B",
    x"395A4E10",
    x"395A32C8",
    x"395A1783",
    x"3959FC42",
    x"3959E104",
    x"3959C5C9",
    x"3959AA92",
    x"39598F5F",
    x"3959742F",
    x"39595902",
    x"39593DD8",
    x"395922B2",
    x"39590790",
    x"3958EC70",
    x"3958D155",
    x"3958B63C",
    x"39589B27",
    x"39588015",
    x"39586507",
    x"395849FC",
    x"39582EF4",
    x"395813F0",
    x"3957F8EF",
    x"3957DDF2",
    x"3957C2F8",
    x"3957A801",
    x"39578D0E",
    x"3957721E",
    x"39575731",
    x"39573C48",
    x"39572162",
    x"39570680",
    x"3956EBA1",
    x"3956D0C5",
    x"3956B5ED",
    x"39569B18",
    x"39568046",
    x"39566577",
    x"39564AAC",
    x"39562FE5",
    x"39561520",
    x"3955FA60",
    x"3955DFA2",
    x"3955C4E8",
    x"3955AA31",
    x"39558F7D",
    x"395574CD",
    x"39555A20",
    x"39553F76",
    x"395524D0",
    x"39550A2D",
    x"3954EF8D",
    x"3954D4F1",
    x"3954BA58",
    x"39549FC3",
    x"39548530",
    x"39546AA1",
    x"39545016",
    x"3954358D",
    x"39541B08",
    x"39540086",
    x"3953E608",
    x"3953CB8D",
    x"3953B115",
    x"395396A1",
    x"39537C30",
    x"395361C2",
    x"39534757",
    x"39532CF0",
    x"3953128C",
    x"3952F82B",
    x"3952DDCE",
    x"3952C374",
    x"3952A91D",
    x"39528EC9",
    x"39527479",
    x"39525A2C",
    x"39523FE3",
    x"3952259C",
    x"39520B59",
    x"3951F11A",
    x"3951D6DD",
    x"3951BCA4",
    x"3951A26E",
    x"3951883B",
    x"39516E0C",
    x"395153E0",
    x"395139B7",
    x"39511F91",
    x"3951056F",
    x"3950EB50",
    x"3950D134",
    x"3950B71C",
    x"39509D06",
    x"395082F4",
    x"395068E6",
    x"39504EDA",
    x"395034D2",
    x"39501ACD",
    x"395000CB",
    x"394FE6CD",
    x"394FCCD1",
    x"394FB2DA",
    x"394F98E5",
    x"394F7EF3",
    x"394F6505",
    x"394F4B1A",
    x"394F3132",
    x"394F174E",
    x"394EFD6C",
    x"394EE38E",
    x"394EC9B4",
    x"394EAFDC",
    x"394E9608",
    x"394E7C36",
    x"394E6269",
    x"394E489E",
    x"394E2ED6",
    x"394E1512",
    x"394DFB51",
    x"394DE193",
    x"394DC7D9",
    x"394DAE21",
    x"394D946D",
    x"394D7ABC",
    x"394D610F",
    x"394D4764",
    x"394D2DBD",
    x"394D1419",
    x"394CFA78",
    x"394CE0DA",
    x"394CC73F",
    x"394CADA8",
    x"394C9414",
    x"394C7A83",
    x"394C60F5",
    x"394C476B",
    x"394C2DE4",
    x"394C145F",
    x"394BFADE",
    x"394BE161",
    x"394BC7E6",
    x"394BAE6F",
    x"394B94FA",
    x"394B7B89",
    x"394B621C",
    x"394B48B1",
    x"394B2F49",
    x"394B15E5",
    x"394AFC84",
    x"394AE326",
    x"394AC9CB",
    x"394AB074",
    x"394A971F",
    x"394A7DCE",
    x"394A6480",
    x"394A4B35",
    x"394A31ED",
    x"394A18A8",
    x"3949FF67",
    x"3949E628",
    x"3949CCED",
    x"3949B3B5",
    x"39499A80",
    x"3949814E",
    x"39496820",
    x"39494EF4",
    x"394935CC",
    x"39491CA7",
    x"39490385",
    x"3948EA66",
    x"3948D14A",
    x"3948B832",
    x"39489F1C",
    x"3948860A",
    x"39486CFB",
    x"394853EF",
    x"39483AE6",
    x"394821E0",
    x"394808DD",
    x"3947EFDE",
    x"3947D6E1",
    x"3947BDE8",
    x"3947A4F2",
    x"39478BFF",
    x"3947730F",
    x"39475A22",
    x"39474138",
    x"39472852",
    x"39470F6E",
    x"3946F68E",
    x"3946DDB1",
    x"3946C4D6",
    x"3946ABFF",
    x"3946932B",
    x"39467A5B",
    x"3946618D",
    x"394648C2",
    x"39462FFB",
    x"39461736",
    x"3945FE75",
    x"3945E5B7",
    x"3945CCFB",
    x"3945B443",
    x"39459B8E",
    x"394582DC",
    x"39456A2E",
    x"39455182",
    x"394538D9",
    x"39452034",
    x"39450791",
    x"3944EEF2",
    x"3944D655",
    x"3944BDBC",
    x"3944A526",
    x"39448C93",
    x"39447403",
    x"39445B76",
    x"394442EC",
    x"39442A65",
    x"394411E1",
    x"3943F961",
    x"3943E0E3",
    x"3943C869",
    x"3943AFF1",
    x"3943977D",
    x"39437F0B",
    x"3943669D",
    x"39434E31",
    x"394335C9",
    x"39431D64",
    x"39430502",
    x"3942ECA3",
    x"3942D447",
    x"3942BBEE",
    x"3942A398",
    x"39428B45",
    x"394272F5",
    x"39425AA8",
    x"3942425E",
    x"39422A17",
    x"394211D4",
    x"3941F993",
    x"3941E155",
    x"3941C91B",
    x"3941B0E3",
    x"394198AE",
    x"3941807D",
    x"3941684E",
    x"39415023",
    x"394137FA",
    x"39411FD5",
    x"394107B2",
    x"3940EF93",
    x"3940D776",
    x"3940BF5D",
    x"3940A747",
    x"39408F33",
    x"39407723",
    x"39405F15",
    x"3940470B",
    x"39402F04",
    x"394016FF",
    x"393FFEFE",
    x"393FE700",
    x"393FCF04",
    x"393FB70C",
    x"393F9F16",
    x"393F8724",
    x"393F6F35",
    x"393F5748",
    x"393F3F5F",
    x"393F2778",
    x"393F0F95",
    x"393EF7B4",
    x"393EDFD7",
    x"393EC7FD",
    x"393EB025",
    x"393E9850",
    x"393E807F",
    x"393E68B0",
    x"393E50E5",
    x"393E391C",
    x"393E2156",
    x"393E0994",
    x"393DF1D4",
    x"393DDA17",
    x"393DC25E",
    x"393DAAA7",
    x"393D92F3",
    x"393D7B42",
    x"393D6394",
    x"393D4BE9",
    x"393D3441",
    x"393D1C9C",
    x"393D04FA",
    x"393CED5B",
    x"393CD5BF",
    x"393CBE25",
    x"393CA68F",
    x"393C8EFC",
    x"393C776B",
    x"393C5FDE",
    x"393C4853",
    x"393C30CC",
    x"393C1947",
    x"393C01C5",
    x"393BEA47",
    x"393BD2CB",
    x"393BBB52",
    x"393BA3DC",
    x"393B8C69",
    x"393B74F9",
    x"393B5D8C",
    x"393B4622",
    x"393B2EBA",
    x"393B1756",
    x"393AFFF4",
    x"393AE896",
    x"393AD13A",
    x"393AB9E2",
    x"393AA28C",
    x"393A8B39",
    x"393A73E9",
    x"393A5C9C",
    x"393A4552",
    x"393A2E0B",
    x"393A16C6",
    x"3939FF85",
    x"3939E846",
    x"3939D10B",
    x"3939B9D2",
    x"3939A29C",
    x"39398B6A",
    x"3939743A",
    x"39395D0D",
    x"393945E2",
    x"39392EBB",
    x"39391797",
    x"39390075",
    x"3938E957",
    x"3938D23B",
    x"3938BB22",
    x"3938A40C",
    x"39388CF9",
    x"393875E9",
    x"39385EDB",
    x"393847D1",
    x"393830CA",
    x"393819C5",
    x"393802C3",
    x"3937EBC4",
    x"3937D4C8",
    x"3937BDCF",
    x"3937A6D9",
    x"39378FE5",
    x"393778F5",
    x"39376207",
    x"39374B1C",
    x"39373434",
    x"39371D4F",
    x"3937066D",
    x"3936EF8E",
    x"3936D8B1",
    x"3936C1D7",
    x"3936AB01",
    x"3936942D",
    x"39367D5C",
    x"3936668D",
    x"39364FC2",
    x"393638F9",
    x"39362234",
    x"39360B71",
    x"3935F4B1",
    x"3935DDF4",
    x"3935C739",
    x"3935B082",
    x"393599CD",
    x"3935831B",
    x"39356C6C",
    x"393555C0",
    x"39353F17",
    x"39352870",
    x"393511CD",
    x"3934FB2C",
    x"3934E48E",
    x"3934CDF3",
    x"3934B75B",
    x"3934A0C5",
    x"39348A32",
    x"393473A2",
    x"39345D15",
    x"3934468B",
    x"39343004",
    x"3934197F",
    x"393402FD",
    x"3933EC7E",
    x"3933D602",
    x"3933BF89",
    x"3933A912",
    x"3933929F",
    x"39337C2E",
    x"393365C0",
    x"39334F54",
    x"393338EC",
    x"39332286",
    x"39330C23",
    x"3932F5C3",
    x"3932DF66",
    x"3932C90B",
    x"3932B2B3",
    x"39329C5F",
    x"3932860C",
    x"39326FBD",
    x"39325970",
    x"39324327",
    x"39322CE0",
    x"3932169B",
    x"3932005A",
    x"3931EA1B",
    x"3931D3DF",
    x"3931BDA6",
    x"3931A770",
    x"3931913D",
    x"39317B0C",
    x"393164DE",
    x"39314EB3",
    x"3931388A",
    x"39312264",
    x"39310C42",
    x"3930F621",
    x"3930E004",
    x"3930C9E9",
    x"3930B3D1",
    x"39309DBC",
    x"393087AA",
    x"3930719A",
    x"39305B8E",
    x"39304584",
    x"39302F7C",
    x"39301978",
    x"39300376",
    x"392FED77",
    x"392FD77B",
    x"392FC181",
    x"392FAB8A",
    x"392F9596",
    x"392F7FA5",
    x"392F69B6",
    x"392F53CA",
    x"392F3DE1",
    x"392F27FB",
    x"392F1217",
    x"392EFC36",
    x"392EE658",
    x"392ED07D",
    x"392EBAA4",
    x"392EA4CE",
    x"392E8EFB",
    x"392E792A",
    x"392E635D",
    x"392E4D92",
    x"392E37C9",
    x"392E2204",
    x"392E0C41",
    x"392DF681",
    x"392DE0C3",
    x"392DCB08",
    x"392DB550",
    x"392D9F9B",
    x"392D89E8",
    x"392D7439",
    x"392D5E8B",
    x"392D48E1",
    x"392D3339",
    x"392D1D94",
    x"392D07F2",
    x"392CF252",
    x"392CDCB5",
    x"392CC71B",
    x"392CB183",
    x"392C9BEF",
    x"392C865C",
    x"392C70CD",
    x"392C5B40",
    x"392C45B6",
    x"392C302F",
    x"392C1AAA",
    x"392C0528",
    x"392BEFA9",
    x"392BDA2C",
    x"392BC4B2",
    x"392BAF3B",
    x"392B99C6",
    x"392B8455",
    x"392B6EE5",
    x"392B5979",
    x"392B440F",
    x"392B2EA8",
    x"392B1943",
    x"392B03E1",
    x"392AEE82",
    x"392AD926",
    x"392AC3CC",
    x"392AAE75",
    x"392A9920",
    x"392A83CF",
    x"392A6E7F",
    x"392A5933",
    x"392A43E9",
    x"392A2EA2",
    x"392A195E",
    x"392A041C",
    x"3929EEDD",
    x"3929D9A0",
    x"3929C466",
    x"3929AF2F",
    x"392999FA",
    x"392984C8",
    x"39296F99",
    x"39295A6C",
    x"39294543",
    x"3929301B",
    x"39291AF6",
    x"392905D4",
    x"3928F0B5",
    x"3928DB98",
    x"3928C67E",
    x"3928B167",
    x"39289C52",
    x"39288740",
    x"39287230",
    x"39285D23",
    x"39284819",
    x"39283311",
    x"39281E0C",
    x"39280909",
    x"3927F40A",
    x"3927DF0C",
    x"3927CA12",
    x"3927B51A",
    x"3927A025",
    x"39278B32",
    x"39277642",
    x"39276154",
    x"39274C69",
    x"39273781",
    x"3927229C",
    x"39270DB9",
    x"3926F8D8",
    x"3926E3FA",
    x"3926CF1F",
    x"3926BA47",
    x"3926A571",
    x"3926909D",
    x"39267BCC",
    x"392666FE",
    x"39265233",
    x"39263D6A",
    x"392628A3",
    x"392613E0",
    x"3925FF1E",
    x"3925EA60",
    x"3925D5A4",
    x"3925C0EA",
    x"3925AC34",
    x"3925977F",
    x"392582CE",
    x"39256E1F",
    x"39255972",
    x"392544C8",
    x"39253021",
    x"39251B7C",
    x"392506DA",
    x"3924F23B",
    x"3924DD9E",
    x"3924C903",
    x"3924B46B",
    x"39249FD6",
    x"39248B43",
    x"392476B3",
    x"39246226",
    x"39244D9B",
    x"39243912",
    x"3924248C",
    x"39241009",
    x"3923FB88",
    x"3923E70A",
    x"3923D28F",
    x"3923BE16",
    x"3923A99F",
    x"3923952B",
    x"392380BA",
    x"39236C4B",
    x"392357DF",
    x"39234375",
    x"39232F0E",
    x"39231AA9",
    x"39230647",
    x"3922F1E8",
    x"3922DD8B",
    x"3922C930",
    x"3922B4D8",
    x"3922A083",
    x"39228C30",
    x"392277E0",
    x"39226392",
    x"39224F47",
    x"39223AFF",
    x"392226B8",
    x"39221275",
    x"3921FE34",
    x"3921E9F5",
    x"3921D5B9",
    x"3921C180",
    x"3921AD49",
    x"39219915",
    x"392184E3",
    x"392170B3",
    x"39215C86",
    x"3921485C",
    x"39213434",
    x"3921200F",
    x"39210BEC",
    x"3920F7CC",
    x"3920E3AE",
    x"3920CF93",
    x"3920BB7B",
    x"3920A764",
    x"39209351",
    x"39207F40",
    x"39206B31",
    x"39205725",
    x"3920431B",
    x"39202F14",
    x"39201B0F",
    x"3920070D",
    x"391FF30E",
    x"391FDF10",
    x"391FCB16",
    x"391FB71E",
    x"391FA328",
    x"391F8F35",
    x"391F7B44",
    x"391F6756",
    x"391F536A",
    x"391F3F81",
    x"391F2B9A",
    x"391F17B6",
    x"391F03D5",
    x"391EEFF5",
    x"391EDC19",
    x"391EC83E",
    x"391EB467",
    x"391EA091",
    x"391E8CBE",
    x"391E78EE",
    x"391E6520",
    x"391E5155",
    x"391E3D8C",
    x"391E29C5",
    x"391E1601",
    x"391E0240",
    x"391DEE81",
    x"391DDAC4",
    x"391DC70A",
    x"391DB352",
    x"391D9F9D",
    x"391D8BEB",
    x"391D783A",
    x"391D648C",
    x"391D50E1",
    x"391D3D38",
    x"391D2992",
    x"391D15EE",
    x"391D024C",
    x"391CEEAD",
    x"391CDB11",
    x"391CC777",
    x"391CB3DF",
    x"391CA04A",
    x"391C8CB7",
    x"391C7926",
    x"391C6598",
    x"391C520D",
    x"391C3E84",
    x"391C2AFD",
    x"391C1779",
    x"391C03F7",
    x"391BF078",
    x"391BDCFB",
    x"391BC981",
    x"391BB609",
    x"391BA293",
    x"391B8F20",
    x"391B7BB0",
    x"391B6841",
    x"391B54D6",
    x"391B416C",
    x"391B2E05",
    x"391B1AA1",
    x"391B073F",
    x"391AF3DF",
    x"391AE082",
    x"391ACD27",
    x"391AB9CE",
    x"391AA678",
    x"391A9325",
    x"391A7FD4",
    x"391A6C85",
    x"391A5938",
    x"391A45EE",
    x"391A32A7",
    x"391A1F62",
    x"391A0C1F",
    x"3919F8DF",
    x"3919E5A1",
    x"3919D265",
    x"3919BF2C",
    x"3919ABF6",
    x"391998C1",
    x"3919858F",
    x"39197260",
    x"39195F33",
    x"39194C08",
    x"391938E0",
    x"391925BA",
    x"39191296",
    x"3918FF75",
    x"3918EC56",
    x"3918D93A",
    x"3918C620",
    x"3918B309",
    x"39189FF3",
    x"39188CE1",
    x"391879D0",
    x"391866C2",
    x"391853B6",
    x"391840AD",
    x"39182DA6",
    x"39181AA2",
    x"391807A0",
    x"3917F4A0",
    x"3917E1A3",
    x"3917CEA7",
    x"3917BBAF",
    x"3917A8B9",
    x"391795C5",
    x"391782D3",
    x"39176FE4",
    x"39175CF7",
    x"39174A0D",
    x"39173725",
    x"3917243F",
    x"3917115C",
    x"3916FE7B",
    x"3916EB9C",
    x"3916D8C0",
    x"3916C5E6",
    x"3916B30E",
    x"3916A039",
    x"39168D66",
    x"39167A96",
    x"391667C8",
    x"391654FC",
    x"39164232",
    x"39162F6B",
    x"39161CA6",
    x"391609E4",
    x"3915F724",
    x"3915E466",
    x"3915D1AB",
    x"3915BEF2",
    x"3915AC3B",
    x"39159987",
    x"391586D5",
    x"39157425",
    x"39156178",
    x"39154ECD",
    x"39153C24",
    x"3915297E",
    x"391516DA",
    x"39150438",
    x"3914F199",
    x"3914DEFC",
    x"3914CC61",
    x"3914B9C8",
    x"3914A732",
    x"3914949F",
    x"3914820D",
    x"39146F7E",
    x"39145CF1",
    x"39144A67",
    x"391437DF",
    x"39142559",
    x"391412D5",
    x"39140054",
    x"3913EDD5",
    x"3913DB59",
    x"3913C8DE",
    x"3913B667",
    x"3913A3F1",
    x"3913917E",
    x"39137F0D",
    x"39136C9E",
    x"39135A31",
    x"391347C7",
    x"3913355F",
    x"391322FA",
    x"39131097",
    x"3912FE36",
    x"3912EBD7",
    x"3912D97B",
    x"3912C721",
    x"3912B4C9",
    x"3912A274",
    x"39129020",
    x"39127DD0",
    x"39126B81",
    x"39125935",
    x"391246EB",
    x"391234A3",
    x"3912225D",
    x"3912101A",
    x"3911FDD9",
    x"3911EB9B",
    x"3911D95F",
    x"3911C725",
    x"3911B4ED",
    x"3911A2B7",
    x"39119084",
    x"39117E53",
    x"39116C24",
    x"391159F8",
    x"391147CE",
    x"391135A6",
    x"39112381",
    x"3911115D",
    x"3910FF3C",
    x"3910ED1D",
    x"3910DB01",
    x"3910C8E7",
    x"3910B6CF",
    x"3910A4B9",
    x"391092A6",
    x"39108094",
    x"39106E85",
    x"39105C79",
    x"39104A6E",
    x"39103866",
    x"39102660",
    x"3910145D",
    x"3910025B",
    x"390FF05C",
    x"390FDE5F",
    x"390FCC64",
    x"390FBA6C",
    x"390FA876",
    x"390F9682",
    x"390F8490",
    x"390F72A1",
    x"390F60B3",
    x"390F4EC8",
    x"390F3CE0",
    x"390F2AF9",
    x"390F1915",
    x"390F0733",
    x"390EF553",
    x"390EE376",
    x"390ED19A",
    x"390EBFC1",
    x"390EADEA",
    x"390E9C16",
    x"390E8A43",
    x"390E7873",
    x"390E66A5",
    x"390E54DA",
    x"390E4310",
    x"390E3149",
    x"390E1F84",
    x"390E0DC1",
    x"390DFC00",
    x"390DEA42",
    x"390DD886",
    x"390DC6CC",
    x"390DB514",
    x"390DA35F",
    x"390D91AB",
    x"390D7FFA",
    x"390D6E4B",
    x"390D5C9F",
    x"390D4AF4",
    x"390D394C",
    x"390D27A6",
    x"390D1602",
    x"390D0460",
    x"390CF2C1",
    x"390CE124",
    x"390CCF88",
    x"390CBDF0",
    x"390CAC59",
    x"390C9AC5",
    x"390C8932",
    x"390C77A2",
    x"390C6614",
    x"390C5489",
    x"390C42FF",
    x"390C3178",
    x"390C1FF3",
    x"390C0E70",
    x"390BFCEF",
    x"390BEB71",
    x"390BD9F4",
    x"390BC87A",
    x"390BB702",
    x"390BA58D",
    x"390B9419",
    x"390B82A8",
    x"390B7138",
    x"390B5FCB",
    x"390B4E60",
    x"390B3CF8",
    x"390B2B91",
    x"390B1A2D",
    x"390B08CB",
    x"390AF76B",
    x"390AE60D",
    x"390AD4B1",
    x"390AC357",
    x"390AB200",
    x"390AA0AB",
    x"390A8F58",
    x"390A7E07",
    x"390A6CB8",
    x"390A5B6C",
    x"390A4A22",
    x"390A38D9",
    x"390A2793",
    x"390A1650",
    x"390A050E",
    x"3909F3CE",
    x"3909E291",
    x"3909D156",
    x"3909C01D",
    x"3909AEE6",
    x"39099DB1",
    x"39098C7E",
    x"39097B4E",
    x"39096A1F",
    x"390958F3",
    x"390947C9",
    x"390936A1",
    x"3909257B",
    x"39091458",
    x"39090336",
    x"3908F217",
    x"3908E0FA",
    x"3908CFDF",
    x"3908BEC6",
    x"3908ADAF",
    x"39089C9A",
    x"39088B88",
    x"39087A78",
    x"39086969",
    x"3908585D",
    x"39084753",
    x"3908364B",
    x"39082546",
    x"39081442",
    x"39080341",
    x"3907F241",
    x"3907E144",
    x"3907D049",
    x"3907BF50",
    x"3907AE59",
    x"39079D64",
    x"39078C72",
    x"39077B81",
    x"39076A93",
    x"390759A7",
    x"390748BC",
    x"390737D4",
    x"390726EF",
    x"3907160B",
    x"39070529",
    x"3906F449",
    x"3906E36C",
    x"3906D291",
    x"3906C1B7",
    x"3906B0E0",
    x"3906A00B",
    x"39068F38",
    x"39067E67",
    x"39066D99",
    x"39065CCC",
    x"39064C01",
    x"39063B39",
    x"39062A73",
    x"390619AE",
    x"390608EC",
    x"3905F82C",
    x"3905E76E",
    x"3905D6B2",
    x"3905C5F8",
    x"3905B541",
    x"3905A48B",
    x"390593D8",
    x"39058326",
    x"39057277",
    x"390561CA",
    x"3905511E",
    x"39054075",
    x"39052FCE",
    x"39051F29",
    x"39050E86",
    x"3904FDE6",
    x"3904ED47",
    x"3904DCAA",
    x"3904CC10",
    x"3904BB77",
    x"3904AAE1",
    x"39049A4D",
    x"390489BA",
    x"3904792A",
    x"3904689C",
    x"39045810",
    x"39044786",
    x"390436FE",
    x"39042678",
    x"390415F4",
    x"39040573",
    x"3903F4F3",
    x"3903E476",
    x"3903D3FA",
    x"3903C381",
    x"3903B309",
    x"3903A294",
    x"39039221",
    x"390381AF",
    x"39037140",
    x"390360D3",
    x"39035068",
    x"39033FFF",
    x"39032F98",
    x"39031F33",
    x"39030ED0",
    x"3902FE6F",
    x"3902EE10",
    x"3902DDB4",
    x"3902CD59",
    x"3902BD00",
    x"3902ACAA",
    x"39029C55",
    x"39028C03",
    x"39027BB2",
    x"39026B64",
    x"39025B17",
    x"39024ACD",
    x"39023A85",
    x"39022A3E",
    x"390219FA",
    x"390209B8",
    x"3901F978",
    x"3901E93A",
    x"3901D8FD",
    x"3901C8C3",
    x"3901B88B",
    x"3901A855",
    x"39019821",
    x"390187EF",
    x"390177BF",
    x"39016791",
    x"39015765",
    x"3901473B",
    x"39013713",
    x"390126EE",
    x"390116CA",
    x"390106A8",
    x"3900F688",
    x"3900E66A",
    x"3900D64E",
    x"3900C635",
    x"3900B61D",
    x"3900A607",
    x"390095F3",
    x"390085E2",
    x"390075D2",
    x"390065C4",
    x"390055B8",
    x"390045AF",
    x"390035A7",
    x"390025A1",
    x"3900159E",
    x"3900059C",
    x"38FFEB38",
    x"38FFCB3D",
    x"38FFAB46",
    x"38FF8B52",
    x"38FF6B63",
    x"38FF4B77",
    x"38FF2B90",
    x"38FF0BAC",
    x"38FEEBCD",
    x"38FECBF2",
    x"38FEAC1A",
    x"38FE8C46",
    x"38FE6C77",
    x"38FE4CAB",
    x"38FE2CE4",
    x"38FE0D20",
    x"38FDED60",
    x"38FDCDA5",
    x"38FDADED",
    x"38FD8E39",
    x"38FD6E8A",
    x"38FD4EDE",
    x"38FD2F36",
    x"38FD0F92",
    x"38FCEFF2",
    x"38FCD056",
    x"38FCB0BE",
    x"38FC912A",
    x"38FC719A",
    x"38FC520D",
    x"38FC3285",
    x"38FC1301",
    x"38FBF380",
    x"38FBD404",
    x"38FBB48B",
    x"38FB9517",
    x"38FB75A6",
    x"38FB5639",
    x"38FB36D0",
    x"38FB176C",
    x"38FAF80B",
    x"38FAD8AE",
    x"38FAB954",
    x"38FA99FF",
    x"38FA7AAE",
    x"38FA5B61",
    x"38FA3C17",
    x"38FA1CD2",
    x"38F9FD90",
    x"38F9DE52",
    x"38F9BF18",
    x"38F99FE2",
    x"38F980B0",
    x"38F96182",
    x"38F94258",
    x"38F92332",
    x"38F9040F",
    x"38F8E4F1",
    x"38F8C5D6",
    x"38F8A6BF",
    x"38F887AC",
    x"38F8689D",
    x"38F84992",
    x"38F82A8B",
    x"38F80B87",
    x"38F7EC88",
    x"38F7CD8C",
    x"38F7AE95",
    x"38F78FA1",
    x"38F770B1",
    x"38F751C4",
    x"38F732DC",
    x"38F713F8",
    x"38F6F517",
    x"38F6D63A",
    x"38F6B762",
    x"38F6988D",
    x"38F679BB",
    x"38F65AEE",
    x"38F63C25",
    x"38F61D5F",
    x"38F5FE9D",
    x"38F5DFE0",
    x"38F5C125",
    x"38F5A26F",
    x"38F583BD",
    x"38F5650E",
    x"38F54664",
    x"38F527BD",
    x"38F5091A",
    x"38F4EA7A",
    x"38F4CBDF",
    x"38F4AD47",
    x"38F48EB4",
    x"38F47024",
    x"38F45198",
    x"38F4330F",
    x"38F4148B",
    x"38F3F60A",
    x"38F3D78D",
    x"38F3B914",
    x"38F39A9F",
    x"38F37C2E",
    x"38F35DC0",
    x"38F33F56",
    x"38F320F0",
    x"38F3028E",
    x"38F2E430",
    x"38F2C5D5",
    x"38F2A77E",
    x"38F2892B",
    x"38F26ADC",
    x"38F24C90",
    x"38F22E49",
    x"38F21005",
    x"38F1F1C5",
    x"38F1D388",
    x"38F1B550",
    x"38F1971B",
    x"38F178EA",
    x"38F15ABD",
    x"38F13C93",
    x"38F11E6E",
    x"38F1004C",
    x"38F0E22E",
    x"38F0C413",
    x"38F0A5FD",
    x"38F087EA",
    x"38F069DB",
    x"38F04BCF",
    x"38F02DC8",
    x"38F00FC4",
    x"38EFF1C4",
    x"38EFD3C7",
    x"38EFB5CF",
    x"38EF97DA",
    x"38EF79E9",
    x"38EF5BFB",
    x"38EF3E12",
    x"38EF202C",
    x"38EF024A",
    x"38EEE46B",
    x"38EEC691",
    x"38EEA8BA",
    x"38EE8AE6",
    x"38EE6D17",
    x"38EE4F4B",
    x"38EE3183",
    x"38EE13BF",
    x"38EDF5FE",
    x"38EDD841",
    x"38EDBA88",
    x"38ED9CD3",
    x"38ED7F21",
    x"38ED6173",
    x"38ED43C9",
    x"38ED2622",
    x"38ED087F",
    x"38ECEAE0",
    x"38ECCD44",
    x"38ECAFAD",
    x"38EC9218",
    x"38EC7488",
    x"38EC56FB",
    x"38EC3972",
    x"38EC1BED",
    x"38EBFE6B",
    x"38EBE0ED",
    x"38EBC373",
    x"38EBA5FC",
    x"38EB888A",
    x"38EB6B1A",
    x"38EB4DAF",
    x"38EB3047",
    x"38EB12E3",
    x"38EAF582",
    x"38EAD825",
    x"38EABACC",
    x"38EA9D77",
    x"38EA8025",
    x"38EA62D7",
    x"38EA458C",
    x"38EA2845",
    x"38EA0B02",
    x"38E9EDC2",
    x"38E9D087",
    x"38E9B34E",
    x"38E9961A",
    x"38E978E9",
    x"38E95BBB",
    x"38E93E92",
    x"38E9216C",
    x"38E90449",
    x"38E8E72B",
    x"38E8CA10",
    x"38E8ACF8",
    x"38E88FE4",
    x"38E872D4",
    x"38E855C8",
    x"38E838BF",
    x"38E81BBA",
    x"38E7FEB8",
    x"38E7E1BA",
    x"38E7C4BF",
    x"38E7A7C9",
    x"38E78AD6",
    x"38E76DE6",
    x"38E750FA",
    x"38E73412",
    x"38E7172D",
    x"38E6FA4C",
    x"38E6DD6E",
    x"38E6C095",
    x"38E6A3BE",
    x"38E686EC",
    x"38E66A1D",
    x"38E64D51",
    x"38E63089",
    x"38E613C5",
    x"38E5F704",
    x"38E5DA47",
    x"38E5BD8E",
    x"38E5A0D8",
    x"38E58426",
    x"38E56777",
    x"38E54ACC",
    x"38E52E24",
    x"38E51180",
    x"38E4F4E0",
    x"38E4D843",
    x"38E4BBAA",
    x"38E49F14",
    x"38E48282",
    x"38E465F3",
    x"38E44968",
    x"38E42CE1",
    x"38E4105D",
    x"38E3F3DD",
    x"38E3D760",
    x"38E3BAE7",
    x"38E39E71",
    x"38E381FF",
    x"38E36591",
    x"38E34926",
    x"38E32CBF",
    x"38E3105B",
    x"38E2F3FB",
    x"38E2D79E",
    x"38E2BB45",
    x"38E29EEF",
    x"38E2829D",
    x"38E2664E",
    x"38E24A03",
    x"38E22DBC",
    x"38E21178",
    x"38E1F538",
    x"38E1D8FB",
    x"38E1BCC1",
    x"38E1A08B",
    x"38E18459",
    x"38E1682A",
    x"38E14BFF",
    x"38E12FD7",
    x"38E113B3",
    x"38E0F792",
    x"38E0DB75",
    x"38E0BF5C",
    x"38E0A345",
    x"38E08733",
    x"38E06B24",
    x"38E04F18",
    x"38E03310",
    x"38E0170B",
    x"38DFFB0A",
    x"38DFDF0C",
    x"38DFC312",
    x"38DFA71C",
    x"38DF8B29",
    x"38DF6F39",
    x"38DF534D",
    x"38DF3764",
    x"38DF1B7F",
    x"38DEFF9D",
    x"38DEE3BF",
    x"38DEC7E4",
    x"38DEAC0D",
    x"38DE9039",
    x"38DE7469",
    x"38DE589C",
    x"38DE3CD3",
    x"38DE210D",
    x"38DE054B",
    x"38DDE98C",
    x"38DDCDD0",
    x"38DDB218",
    x"38DD9664",
    x"38DD7AB3",
    x"38DD5F05",
    x"38DD435B",
    x"38DD27B4",
    x"38DD0C11",
    x"38DCF071",
    x"38DCD4D5",
    x"38DCB93C",
    x"38DC9DA6",
    x"38DC8214",
    x"38DC6686",
    x"38DC4AFB",
    x"38DC2F73",
    x"38DC13EF",
    x"38DBF86E",
    x"38DBDCF1",
    x"38DBC177",
    x"38DBA601",
    x"38DB8A8D",
    x"38DB6F1E",
    x"38DB53B2",
    x"38DB3849",
    x"38DB1CE4",
    x"38DB0182",
    x"38DAE623",
    x"38DACAC8",
    x"38DAAF71",
    x"38DA941C",
    x"38DA78CC",
    x"38DA5D7E",
    x"38DA4234",
    x"38DA26EE",
    x"38DA0BAA",
    x"38D9F06B",
    x"38D9D52E",
    x"38D9B9F5",
    x"38D99EC0",
    x"38D9838E",
    x"38D9685F",
    x"38D94D34",
    x"38D9320C",
    x"38D916E7",
    x"38D8FBC6",
    x"38D8E0A8",
    x"38D8C58E",
    x"38D8AA77",
    x"38D88F63",
    x"38D87453",
    x"38D85946",
    x"38D83E3D",
    x"38D82336",
    x"38D80834",
    x"38D7ED34",
    x"38D7D238",
    x"38D7B740",
    x"38D79C4B",
    x"38D78159",
    x"38D7666A",
    x"38D74B7F",
    x"38D73097",
    x"38D715B3",
    x"38D6FAD2",
    x"38D6DFF4",
    x"38D6C51A",
    x"38D6AA43",
    x"38D68F6F",
    x"38D6749F",
    x"38D659D2",
    x"38D63F09",
    x"38D62443",
    x"38D60980",
    x"38D5EEC0",
    x"38D5D404",
    x"38D5B94B",
    x"38D59E96",
    x"38D583E4",
    x"38D56935",
    x"38D54E89",
    x"38D533E1",
    x"38D5193C",
    x"38D4FE9B",
    x"38D4E3FD",
    x"38D4C962",
    x"38D4AECA",
    x"38D49436",
    x"38D479A5",
    x"38D45F18",
    x"38D4448D",
    x"38D42A07",
    x"38D40F83",
    x"38D3F503",
    x"38D3DA86",
    x"38D3C00C",
    x"38D3A596",
    x"38D38B23",
    x"38D370B3",
    x"38D35646",
    x"38D33BDD",
    x"38D32177",
    x"38D30715",
    x"38D2ECB6",
    x"38D2D25A",
    x"38D2B801",
    x"38D29DAC",
    x"38D2835A",
    x"38D2690B",
    x"38D24EBF",
    x"38D23477",
    x"38D21A32",
    x"38D1FFF1",
    x"38D1E5B2",
    x"38D1CB77",
    x"38D1B13F",
    x"38D1970B",
    x"38D17CDA",
    x"38D162AC",
    x"38D14881",
    x"38D12E5A",
    x"38D11435",
    x"38D0FA15",
    x"38D0DFF7",
    x"38D0C5DD",
    x"38D0ABC5",
    x"38D091B2",
    x"38D077A1",
    x"38D05D94",
    x"38D0438A",
    x"38D02983",
    x"38D00F7F",
    x"38CFF57F",
    x"38CFDB82",
    x"38CFC188",
    x"38CFA791",
    x"38CF8D9E",
    x"38CF73AE",
    x"38CF59C1",
    x"38CF3FD8",
    x"38CF25F1",
    x"38CF0C0E",
    x"38CEF22E",
    x"38CED852",
    x"38CEBE78",
    x"38CEA4A2",
    x"38CE8ACF",
    x"38CE70FF",
    x"38CE5733",
    x"38CE3D69",
    x"38CE23A3",
    x"38CE09E1",
    x"38CDF021",
    x"38CDD665",
    x"38CDBCAB",
    x"38CDA2F5",
    x"38CD8943",
    x"38CD6F93",
    x"38CD55E7",
    x"38CD3C3E",
    x"38CD2298",
    x"38CD08F5",
    x"38CCEF55",
    x"38CCD5B9",
    x"38CCBC20",
    x"38CCA28A",
    x"38CC88F7",
    x"38CC6F68",
    x"38CC55DC",
    x"38CC3C52",
    x"38CC22CC",
    x"38CC094A",
    x"38CBEFCA",
    x"38CBD64E",
    x"38CBBCD5",
    x"38CBA35F",
    x"38CB89EC",
    x"38CB707C",
    x"38CB5710",
    x"38CB3DA6",
    x"38CB2440",
    x"38CB0ADD",
    x"38CAF17D",
    x"38CAD821",
    x"38CABEC7",
    x"38CAA571",
    x"38CA8C1E",
    x"38CA72CE",
    x"38CA5981",
    x"38CA4038",
    x"38CA26F1",
    x"38CA0DAE",
    x"38C9F46E",
    x"38C9DB31",
    x"38C9C1F7",
    x"38C9A8C0",
    x"38C98F8D",
    x"38C9765D",
    x"38C95D2F",
    x"38C94405",
    x"38C92ADE",
    x"38C911BA",
    x"38C8F89A",
    x"38C8DF7C",
    x"38C8C662",
    x"38C8AD4B",
    x"38C89437",
    x"38C87B26",
    x"38C86218",
    x"38C8490D",
    x"38C83006",
    x"38C81701",
    x"38C7FE00",
    x"38C7E502",
    x"38C7CC07",
    x"38C7B30F",
    x"38C79A1A",
    x"38C78128",
    x"38C7683A",
    x"38C74F4E",
    x"38C73666",
    x"38C71D80",
    x"38C7049E",
    x"38C6EBBF",
    x"38C6D2E3",
    x"38C6BA0B",
    x"38C6A135",
    x"38C68862",
    x"38C66F93",
    x"38C656C6",
    x"38C63DFD",
    x"38C62537",
    x"38C60C74",
    x"38C5F3B4",
    x"38C5DAF7",
    x"38C5C23D",
    x"38C5A986",
    x"38C590D3",
    x"38C57822",
    x"38C55F75",
    x"38C546CA",
    x"38C52E23",
    x"38C5157F",
    x"38C4FCDE",
    x"38C4E43F",
    x"38C4CBA4",
    x"38C4B30D",
    x"38C49A78",
    x"38C481E6",
    x"38C46957",
    x"38C450CC",
    x"38C43843",
    x"38C41FBE",
    x"38C4073B",
    x"38C3EEBC",
    x"38C3D63F",
    x"38C3BDC6",
    x"38C3A550",
    x"38C38CDD",
    x"38C3746D",
    x"38C35C00",
    x"38C34396",
    x"38C32B2F",
    x"38C312CB",
    x"38C2FA6A",
    x"38C2E20C",
    x"38C2C9B2",
    x"38C2B15A",
    x"38C29905",
    x"38C280B4",
    x"38C26865",
    x"38C2501A",
    x"38C237D1",
    x"38C21F8C",
    x"38C20749",
    x"38C1EF0A",
    x"38C1D6CD",
    x"38C1BE94",
    x"38C1A65E",
    x"38C18E2B",
    x"38C175FA",
    x"38C15DCD",
    x"38C145A3",
    x"38C12D7C",
    x"38C11557",
    x"38C0FD36",
    x"38C0E518",
    x"38C0CCFD",
    x"38C0B4E5",
    x"38C09CD0",
    x"38C084BE",
    x"38C06CAF",
    x"38C054A3",
    x"38C03C99",
    x"38C02493",
    x"38C00C90",
    x"38BFF490",
    x"38BFDC93",
    x"38BFC499",
    x"38BFACA2",
    x"38BF94AE",
    x"38BF7CBD",
    x"38BF64CF",
    x"38BF4CE4",
    x"38BF34FC",
    x"38BF1D16",
    x"38BF0534",
    x"38BEED55",
    x"38BED579",
    x"38BEBDA0",
    x"38BEA5CA",
    x"38BE8DF6",
    x"38BE7626",
    x"38BE5E59",
    x"38BE468E",
    x"38BE2EC7",
    x"38BE1703",
    x"38BDFF41",
    x"38BDE783",
    x"38BDCFC7",
    x"38BDB80F",
    x"38BDA059",
    x"38BD88A7",
    x"38BD70F7",
    x"38BD594B",
    x"38BD41A1",
    x"38BD29FA",
    x"38BD1256",
    x"38BCFAB6",
    x"38BCE318",
    x"38BCCB7D",
    x"38BCB3E5",
    x"38BC9C50",
    x"38BC84BE",
    x"38BC6D2F",
    x"38BC55A3",
    x"38BC3E19",
    x"38BC2693",
    x"38BC0F10",
    x"38BBF78F",
    x"38BBE012",
    x"38BBC897",
    x"38BBB120",
    x"38BB99AB",
    x"38BB8239",
    x"38BB6ACA",
    x"38BB535F",
    x"38BB3BF6",
    x"38BB2490",
    x"38BB0D2C",
    x"38BAF5CC",
    x"38BADE6F",
    x"38BAC715",
    x"38BAAFBD",
    x"38BA9869",
    x"38BA8117",
    x"38BA69C8",
    x"38BA527D",
    x"38BA3B34",
    x"38BA23EE",
    x"38BA0CAB",
    x"38B9F56B",
    x"38B9DE2D",
    x"38B9C6F3",
    x"38B9AFBC",
    x"38B99887",
    x"38B98156",
    x"38B96A27",
    x"38B952FB",
    x"38B93BD2",
    x"38B924AC",
    x"38B90D89",
    x"38B8F669",
    x"38B8DF4B",
    x"38B8C831",
    x"38B8B119",
    x"38B89A05",
    x"38B882F3",
    x"38B86BE4",
    x"38B854D8",
    x"38B83DCF",
    x"38B826C8",
    x"38B80FC5",
    x"38B7F8C4",
    x"38B7E1C7",
    x"38B7CACC",
    x"38B7B3D4",
    x"38B79CDF",
    x"38B785ED",
    x"38B76EFE",
    x"38B75811",
    x"38B74128",
    x"38B72A41",
    x"38B7135D",
    x"38B6FC7C",
    x"38B6E59E",
    x"38B6CEC3",
    x"38B6B7EA",
    x"38B6A115",
    x"38B68A42",
    x"38B67372",
    x"38B65CA5",
    x"38B645DB",
    x"38B62F14",
    x"38B6184F",
    x"38B6018D",
    x"38B5EACF",
    x"38B5D413",
    x"38B5BD5A",
    x"38B5A6A3",
    x"38B58FF0",
    x"38B5793F",
    x"38B56292",
    x"38B54BE7",
    x"38B5353F",
    x"38B51E99",
    x"38B507F7",
    x"38B4F158",
    x"38B4DABB",
    x"38B4C421",
    x"38B4AD8A",
    x"38B496F5",
    x"38B48064",
    x"38B469D5",
    x"38B4534A",
    x"38B43CC1",
    x"38B4263A",
    x"38B40FB7",
    x"38B3F936",
    x"38B3E2B9",
    x"38B3CC3E",
    x"38B3B5C6",
    x"38B39F50",
    x"38B388DE",
    x"38B3726E",
    x"38B35C01",
    x"38B34597",
    x"38B32F30",
    x"38B318CB",
    x"38B3026A",
    x"38B2EC0B",
    x"38B2D5AF",
    x"38B2BF55",
    x"38B2A8FF",
    x"38B292AB",
    x"38B27C5A",
    x"38B2660C",
    x"38B24FC1",
    x"38B23978",
    x"38B22332",
    x"38B20CEF",
    x"38B1F6AF",
    x"38B1E071",
    x"38B1CA37",
    x"38B1B3FF",
    x"38B19DCA",
    x"38B18797",
    x"38B17168",
    x"38B15B3B",
    x"38B14511",
    x"38B12EEA",
    x"38B118C5",
    x"38B102A4",
    x"38B0EC85",
    x"38B0D669",
    x"38B0C04F",
    x"38B0AA38",
    x"38B09425",
    x"38B07E13",
    x"38B06805",
    x"38B051F9",
    x"38B03BF1",
    x"38B025EA",
    x"38B00FE7",
    x"38AFF9E6",
    x"38AFE3E9",
    x"38AFCDED",
    x"38AFB7F5",
    x"38AFA1FF",
    x"38AF8C0D",
    x"38AF761C",
    x"38AF602F",
    x"38AF4A44",
    x"38AF345D",
    x"38AF1E77",
    x"38AF0895",
    x"38AEF2B5",
    x"38AEDCD8",
    x"38AEC6FE",
    x"38AEB126",
    x"38AE9B52",
    x"38AE8580",
    x"38AE6FB0",
    x"38AE59E4",
    x"38AE441A",
    x"38AE2E53",
    x"38AE188E",
    x"38AE02CD",
    x"38ADED0E",
    x"38ADD751",
    x"38ADC198",
    x"38ADABE1",
    x"38AD962D",
    x"38AD807B",
    x"38AD6ACD",
    x"38AD5521",
    x"38AD3F77",
    x"38AD29D1",
    x"38AD142D",
    x"38ACFE8C",
    x"38ACE8ED",
    x"38ACD352",
    x"38ACBDB8",
    x"38ACA822",
    x"38AC928E",
    x"38AC7CFD",
    x"38AC676F",
    x"38AC51E4",
    x"38AC3C5B",
    x"38AC26D4",
    x"38AC1151",
    x"38ABFBD0",
    x"38ABE652",
    x"38ABD0D7",
    x"38ABBB5E",
    x"38ABA5E8",
    x"38AB9074",
    x"38AB7B04",
    x"38AB6596",
    x"38AB502A",
    x"38AB3AC2",
    x"38AB255C",
    x"38AB0FF8",
    x"38AAFA98",
    x"38AAE53A",
    x"38AACFDE",
    x"38AABA86",
    x"38AAA530",
    x"38AA8FDC",
    x"38AA7A8C",
    x"38AA653E",
    x"38AA4FF2",
    x"38AA3AAA",
    x"38AA2564",
    x"38AA1020",
    x"38A9FAE0",
    x"38A9E5A2",
    x"38A9D066",
    x"38A9BB2E",
    x"38A9A5F7",
    x"38A990C4",
    x"38A97B93",
    x"38A96665",
    x"38A9513A",
    x"38A93C11",
    x"38A926EB",
    x"38A911C7",
    x"38A8FCA6",
    x"38A8E788",
    x"38A8D26C",
    x"38A8BD53",
    x"38A8A83D",
    x"38A89329",
    x"38A87E18",
    x"38A8690A",
    x"38A853FE",
    x"38A83EF5",
    x"38A829EE",
    x"38A814EA",
    x"38A7FFE9",
    x"38A7EAEA",
    x"38A7D5EE",
    x"38A7C0F5",
    x"38A7ABFE",
    x"38A7970A",
    x"38A78218",
    x"38A76D29",
    x"38A7583D",
    x"38A74353",
    x"38A72E6C",
    x"38A71988",
    x"38A704A6",
    x"38A6EFC6",
    x"38A6DAEA",
    x"38A6C610",
    x"38A6B138",
    x"38A69C63",
    x"38A68791",
    x"38A672C2",
    x"38A65DF4",
    x"38A6492A",
    x"38A63462",
    x"38A61F9D",
    x"38A60ADA",
    x"38A5F61A",
    x"38A5E15D",
    x"38A5CCA2",
    x"38A5B7EA",
    x"38A5A334",
    x"38A58E81",
    x"38A579D0",
    x"38A56522",
    x"38A55077",
    x"38A53BCE",
    x"38A52728",
    x"38A51284",
    x"38A4FDE3",
    x"38A4E945",
    x"38A4D4A9",
    x"38A4C010",
    x"38A4AB79",
    x"38A496E5",
    x"38A48253",
    x"38A46DC4",
    x"38A45938",
    x"38A444AE",
    x"38A43027",
    x"38A41BA2",
    x"38A40720",
    x"38A3F2A0",
    x"38A3DE23",
    x"38A3C9A9",
    x"38A3B531",
    x"38A3A0BB",
    x"38A38C49",
    x"38A377D8",
    x"38A3636B",
    x"38A34EFF",
    x"38A33A97",
    x"38A32631",
    x"38A311CD",
    x"38A2FD6C",
    x"38A2E90E",
    x"38A2D4B2",
    x"38A2C059",
    x"38A2AC02",
    x"38A297AE",
    x"38A2835C",
    x"38A26F0D",
    x"38A25AC0",
    x"38A24676",
    x"38A2322F",
    x"38A21DEA",
    x"38A209A7",
    x"38A1F567",
    x"38A1E12A",
    x"38A1CCEF",
    x"38A1B8B7",
    x"38A1A481",
    x"38A1904E",
    x"38A17C1D",
    x"38A167EE",
    x"38A153C3",
    x"38A13F9A",
    x"38A12B73",
    x"38A1174F",
    x"38A1032D",
    x"38A0EF0E",
    x"38A0DAF1",
    x"38A0C6D7",
    x"38A0B2C0",
    x"38A09EAA",
    x"38A08A98",
    x"38A07688",
    x"38A0627A",
    x"38A04E6F",
    x"38A03A67",
    x"38A02661",
    x"38A0125D",
    x"389FFE5C",
    x"389FEA5D",
    x"389FD661",
    x"389FC268",
    x"389FAE71",
    x"389F9A7C",
    x"389F868A",
    x"389F729B",
    x"389F5EAE",
    x"389F4AC3",
    x"389F36DB",
    x"389F22F5",
    x"389F0F12",
    x"389EFB31",
    x"389EE753",
    x"389ED378",
    x"389EBF9E",
    x"389EABC8",
    x"389E97F3",
    x"389E8422",
    x"389E7052",
    x"389E5C86",
    x"389E48BB",
    x"389E34F3",
    x"389E212E",
    x"389E0D6B",
    x"389DF9AB",
    x"389DE5ED",
    x"389DD231",
    x"389DBE78",
    x"389DAAC2",
    x"389D970E",
    x"389D835C",
    x"389D6FAD",
    x"389D5C00",
    x"389D4856",
    x"389D34AE",
    x"389D2109",
    x"389D0D66",
    x"389CF9C5",
    x"389CE627",
    x"389CD28C",
    x"389CBEF3",
    x"389CAB5C",
    x"389C97C8",
    x"389C8436",
    x"389C70A7",
    x"389C5D1A",
    x"389C498F",
    x"389C3607",
    x"389C2282",
    x"389C0EFF",
    x"389BFB7E",
    x"389BE800",
    x"389BD484",
    x"389BC10B",
    x"389BAD94",
    x"389B9A1F",
    x"389B86AD",
    x"389B733E",
    x"389B5FD1",
    x"389B4C66",
    x"389B38FD",
    x"389B2597",
    x"389B1234",
    x"389AFED3",
    x"389AEB74",
    x"389AD818",
    x"389AC4BE",
    x"389AB167",
    x"389A9E12",
    x"389A8ABF",
    x"389A776F",
    x"389A6422",
    x"389A50D6",
    x"389A3D8D",
    x"389A2A47",
    x"389A1703",
    x"389A03C1",
    x"3899F082",
    x"3899DD45",
    x"3899CA0A",
    x"3899B6D2",
    x"3899A39D",
    x"3899906A",
    x"38997D39",
    x"38996A0A",
    x"389956DE",
    x"389943B4",
    x"3899308D",
    x"38991D68",
    x"38990A46",
    x"3898F726",
    x"3898E408",
    x"3898D0ED",
    x"3898BDD4",
    x"3898AABD",
    x"389897A9",
    x"38988497",
    x"38987188",
    x"38985E7B",
    x"38984B70",
    x"38983868",
    x"38982562",
    x"3898125F",
    x"3897FF5E",
    x"3897EC5F",
    x"3897D963",
    x"3897C669",
    x"3897B371",
    x"3897A07C",
    x"38978D89",
    x"38977A98",
    x"389767AA",
    x"389754BE",
    x"389741D5",
    x"38972EEE",
    x"38971C09",
    x"38970927",
    x"3896F647",
    x"3896E369",
    x"3896D08E",
    x"3896BDB5",
    x"3896AADF",
    x"3896980B",
    x"38968539",
    x"38967269",
    x"38965F9C",
    x"38964CD1",
    x"38963A09",
    x"38962743",
    x"3896147F",
    x"389601BE",
    x"3895EEFF",
    x"3895DC42",
    x"3895C988",
    x"3895B6D0",
    x"3895A41A",
    x"38959167",
    x"38957EB6",
    x"38956C07",
    x"3895595B",
    x"389546B1",
    x"38953409",
    x"38952164",
    x"38950EC1",
    x"3894FC20",
    x"3894E982",
    x"3894D6E5",
    x"3894C44C",
    x"3894B1B4",
    x"38949F1F",
    x"38948C8D",
    x"389479FC",
    x"3894676E",
    x"389454E2",
    x"38944259",
    x"38942FD2",
    x"38941D4D",
    x"38940ACA",
    x"3893F84A",
    x"3893E5CC",
    x"3893D351",
    x"3893C0D8",
    x"3893AE61",
    x"38939BEC",
    x"3893897A",
    x"3893770A",
    x"3893649C",
    x"38935230",
    x"38933FC7",
    x"38932D60",
    x"38931AFC",
    x"3893089A",
    x"3892F63A",
    x"3892E3DC",
    x"3892D181",
    x"3892BF28",
    x"3892ACD1",
    x"38929A7D",
    x"3892882A",
    x"389275DB",
    x"3892638D",
    x"38925142",
    x"38923EF9",
    x"38922CB2",
    x"38921A6D",
    x"3892082B",
    x"3891F5EB",
    x"3891E3AE",
    x"3891D173",
    x"3891BF39",
    x"3891AD03",
    x"38919ACE",
    x"3891889C",
    x"3891766C",
    x"3891643E",
    x"38915213",
    x"38913FEA",
    x"38912DC3",
    x"38911B9E",
    x"3891097C",
    x"3890F75C",
    x"3890E53E",
    x"3890D323",
    x"3890C10A",
    x"3890AEF3",
    x"38909CDE",
    x"38908ACB",
    x"389078BB",
    x"389066AD",
    x"389054A1",
    x"38904298",
    x"38903091",
    x"38901E8C",
    x"38900C89",
    x"388FFA89",
    x"388FE88A",
    x"388FD68F",
    x"388FC495",
    x"388FB29D",
    x"388FA0A8",
    x"388F8EB5",
    x"388F7CC5",
    x"388F6AD6",
    x"388F58EA",
    x"388F4700",
    x"388F3518",
    x"388F2333",
    x"388F114F",
    x"388EFF6E",
    x"388EED8F",
    x"388EDBB3",
    x"388EC9D8",
    x"388EB800",
    x"388EA62A",
    x"388E9457",
    x"388E8285",
    x"388E70B6",
    x"388E5EE9",
    x"388E4D1E",
    x"388E3B56",
    x"388E2990",
    x"388E17CC",
    x"388E060A",
    x"388DF44A",
    x"388DE28D",
    x"388DD0D1",
    x"388DBF18",
    x"388DAD62",
    x"388D9BAD",
    x"388D89FB",
    x"388D784B",
    x"388D669D",
    x"388D54F1",
    x"388D4347",
    x"388D31A0",
    x"388D1FFB",
    x"388D0E58",
    x"388CFCB7",
    x"388CEB19",
    x"388CD97D",
    x"388CC7E3",
    x"388CB64B",
    x"388CA4B5",
    x"388C9321",
    x"388C8190",
    x"388C7001",
    x"388C5E74",
    x"388C4CE9",
    x"388C3B61",
    x"388C29DB",
    x"388C1856",
    x"388C06D5",
    x"388BF555",
    x"388BE3D7",
    x"388BD25C",
    x"388BC0E3",
    x"388BAF6C",
    x"388B9DF7",
    x"388B8C84",
    x"388B7B14",
    x"388B69A5",
    x"388B5839",
    x"388B46CF",
    x"388B3568",
    x"388B2402",
    x"388B129F",
    x"388B013D",
    x"388AEFDE",
    x"388ADE81",
    x"388ACD27",
    x"388ABBCE",
    x"388AAA78",
    x"388A9923",
    x"388A87D1",
    x"388A7681",
    x"388A6534",
    x"388A53E8",
    x"388A429F",
    x"388A3157",
    x"388A2012",
    x"388A0ECF",
    x"3889FD8F",
    x"3889EC50",
    x"3889DB14",
    x"3889C9D9",
    x"3889B8A1",
    x"3889A76B",
    x"38899637",
    x"38898506",
    x"388973D6",
    x"388962A9",
    x"3889517D",
    x"38894054",
    x"38892F2D",
    x"38891E08",
    x"38890CE6",
    x"3888FBC5",
    x"3888EAA7",
    x"3888D98B",
    x"3888C870",
    x"3888B758",
    x"3888A643",
    x"3888952F",
    x"3888841D",
    x"3888730E",
    x"38886201",
    x"388850F5",
    x"38883FEC",
    x"38882EE5",
    x"38881DE1",
    x"38880CDE",
    x"3887FBDD",
    x"3887EADF",
    x"3887D9E3",
    x"3887C8E8",
    x"3887B7F0",
    x"3887A6FA",
    x"38879607",
    x"38878515",
    x"38877425",
    x"38876338",
    x"3887524D",
    x"38874163",
    x"3887307C",
    x"38871F97",
    x"38870EB4",
    x"3886FDD4",
    x"3886ECF5",
    x"3886DC18",
    x"3886CB3E",
    x"3886BA66",
    x"3886A98F",
    x"388698BB",
    x"388687E9",
    x"38867719",
    x"3886664B",
    x"38865580",
    x"388644B6",
    x"388633EE",
    x"38862329",
    x"38861266",
    x"388601A4",
    x"3885F0E5",
    x"3885E028",
    x"3885CF6D",
    x"3885BEB4",
    x"3885ADFD",
    x"38859D49",
    x"38858C96",
    x"38857BE6",
    x"38856B37",
    x"38855A8B",
    x"388549E1",
    x"38853938",
    x"38852892",
    x"388517EE",
    x"3885074C",
    x"3884F6AC",
    x"3884E60F",
    x"3884D573",
    x"3884C4D9",
    x"3884B442",
    x"3884A3AC",
    x"38849319",
    x"38848287",
    x"388471F8",
    x"3884616B",
    x"388450E0",
    x"38844057",
    x"38842FD0",
    x"38841F4B",
    x"38840EC8",
    x"3883FE47",
    x"3883EDC8",
    x"3883DD4C",
    x"3883CCD1",
    x"3883BC58",
    x"3883ABE2",
    x"38839B6D",
    x"38838AFB",
    x"38837A8B",
    x"38836A1C",
    x"388359B0",
    x"38834946",
    x"388338DE",
    x"38832878",
    x"38831814",
    x"388307B2",
    x"3882F752",
    x"3882E6F4",
    x"3882D698",
    x"3882C63E",
    x"3882B5E6",
    x"3882A591",
    x"3882953D",
    x"388284EB",
    x"3882749C",
    x"3882644E",
    x"38825403",
    x"388243B9",
    x"38823372",
    x"3882232C",
    x"388212E9",
    x"388202A8",
    x"3881F268",
    x"3881E22B",
    x"3881D1F0",
    x"3881C1B7",
    x"3881B17F",
    x"3881A14A",
    x"38819117",
    x"388180E6",
    x"388170B7",
    x"3881608A",
    x"3881505F",
    x"38814036",
    x"3881300F",
    x"38811FEA",
    x"38810FC7",
    x"3880FFA6",
    x"3880EF87",
    x"3880DF6A",
    x"3880CF4F",
    x"3880BF36",
    x"3880AF1F",
    x"38809F0A",
    x"38808EF7",
    x"38807EE7",
    x"38806ED8",
    x"38805ECB",
    x"38804EC0",
    x"38803EB7",
    x"38802EB0",
    x"38801EAB",
    x"38800EA9",
    x"387FFD50",
    x"387FDD52",
    x"387FBD58",
    x"387F9D63",
    x"387F7D71",
    x"387F5D83",
    x"387F3D9A",
    x"387F1DB4",
    x"387EFDD2",
    x"387EDDF4",
    x"387EBE1B",
    x"387E9E45",
    x"387E7E73",
    x"387E5EA5",
    x"387E3EDB",
    x"387E1F15",
    x"387DFF54",
    x"387DDF96",
    x"387DBFDC",
    x"387DA026",
    x"387D8074",
    x"387D60C6",
    x"387D411B",
    x"387D2175",
    x"387D01D3",
    x"387CE235",
    x"387CC29B",
    x"387CA304",
    x"387C8372",
    x"387C63E3",
    x"387C4459",
    x"387C24D2",
    x"387C0550",
    x"387BE5D1",
    x"387BC656",
    x"387BA6DF",
    x"387B876C",
    x"387B67FD",
    x"387B4892",
    x"387B292B",
    x"387B09C8",
    x"387AEA69",
    x"387ACB0E",
    x"387AABB6",
    x"387A8C63",
    x"387A6D13",
    x"387A4DC7",
    x"387A2E80",
    x"387A0F3C",
    x"3879EFFC",
    x"3879D0C0",
    x"3879B188",
    x"38799253",
    x"38797323",
    x"387953F7",
    x"387934CE",
    x"387915A9",
    x"3878F689",
    x"3878D76C",
    x"3878B853",
    x"3878993E",
    x"38787A2C",
    x"38785B1F",
    x"38783C16",
    x"38781D10",
    x"3877FE0E",
    x"3877DF11",
    x"3877C017",
    x"3877A121",
    x"3877822E",
    x"38776340",
    x"38774456",
    x"3877256F",
    x"3877068C",
    x"3876E7AD",
    x"3876C8D2",
    x"3876A9FB",
    x"38768B28",
    x"38766C58",
    x"38764D8D",
    x"38762EC5",
    x"38761001",
    x"3875F141",
    x"3875D285",
    x"3875B3CC",
    x"38759518",
    x"38757667",
    x"387557BA",
    x"38753911",
    x"38751A6C",
    x"3874FBCA",
    x"3874DD2D",
    x"3874BE93",
    x"38749FFD",
    x"3874816B",
    x"387462DD",
    x"38744452",
    x"387425CC",
    x"38740749",
    x"3873E8CA",
    x"3873CA4F",
    x"3873ABD7",
    x"38738D64",
    x"38736EF4",
    x"38735088",
    x"38733220",
    x"387313BC",
    x"3872F55B",
    x"3872D6FE",
    x"3872B8A5",
    x"38729A50",
    x"38727BFF",
    x"38725DB1",
    x"38723F67",
    x"38722121",
    x"387202DF",
    x"3871E4A0",
    x"3871C666",
    x"3871A82F",
    x"387189FC",
    x"38716BCC",
    x"38714DA1",
    x"38712F79",
    x"38711155",
    x"3870F335",
    x"3870D518",
    x"3870B6FF",
    x"387098EA",
    x"38707AD9",
    x"38705CCC",
    x"38703EC2",
    x"387020BC",
    x"387002BA",
    x"386FE4BB",
    x"386FC6C1",
    x"386FA8CA",
    x"386F8AD6",
    x"386F6CE7",
    x"386F4EFB",
    x"386F3113",
    x"386F132F",
    x"386EF54E",
    x"386ED772",
    x"386EB998",
    x"386E9BC3",
    x"386E7DF2",
    x"386E6024",
    x"386E425A",
    x"386E2493",
    x"386E06D0",
    x"386DE911",
    x"386DCB56",
    x"386DAD9F",
    x"386D8FEB",
    x"386D723B",
    x"386D548E",
    x"386D36E5",
    x"386D1940",
    x"386CFB9F",
    x"386CDE02",
    x"386CC068",
    x"386CA2D1",
    x"386C853F",
    x"386C67B0",
    x"386C4A25",
    x"386C2C9E",
    x"386C0F1A",
    x"386BF19A",
    x"386BD41D",
    x"386BB6A5",
    x"386B9930",
    x"386B7BBE",
    x"386B5E51",
    x"386B40E7",
    x"386B2381",
    x"386B061E",
    x"386AE8BF",
    x"386ACB64",
    x"386AAE0C",
    x"386A90B8",
    x"386A7368",
    x"386A561B",
    x"386A38D3",
    x"386A1B8D",
    x"3869FE4C",
    x"3869E10E",
    x"3869C3D3",
    x"3869A69D",
    x"3869896A",
    x"38696C3A",
    x"38694F0F",
    x"386931E7",
    x"386914C2",
    x"3868F7A1",
    x"3868DA84",
    x"3868BD6B",
    x"3868A055",
    x"38688343",
    x"38686634",
    x"38684929",
    x"38682C22",
    x"38680F1E",
    x"3867F21E",
    x"3867D522",
    x"3867B829",
    x"38679B34",
    x"38677E42",
    x"38676154",
    x"3867446A",
    x"38672783",
    x"38670AA0",
    x"3866EDC0",
    x"3866D0E4",
    x"3866B40C",
    x"38669737",
    x"38667A66",
    x"38665D99",
    x"386640CF",
    x"38662408",
    x"38660746",
    x"3865EA87",
    x"3865CDCB",
    x"3865B113",
    x"3865945F",
    x"386577AE",
    x"38655B01",
    x"38653E57",
    x"386521B1",
    x"3865050F",
    x"3864E870",
    x"3864CBD5",
    x"3864AF3D",
    x"386492A9",
    x"38647618",
    x"3864598B",
    x"38643D02",
    x"3864207C",
    x"386403FA",
    x"3863E77B",
    x"3863CB00",
    x"3863AE89",
    x"38639214",
    x"386375A4",
    x"38635937",
    x"38633CCE",
    x"38632068",
    x"38630406",
    x"3862E7A7",
    x"3862CB4C",
    x"3862AEF4",
    x"386292A0",
    x"3862764F",
    x"38625A02",
    x"38623DB9",
    x"38622173",
    x"38620530",
    x"3861E8F2",
    x"3861CCB6",
    x"3861B07E",
    x"3861944A",
    x"38617819",
    x"38615BEC",
    x"38613FC2",
    x"3861239C",
    x"38610779",
    x"3860EB5A",
    x"3860CF3F",
    x"3860B326",
    x"38609712",
    x"38607B01",
    x"38605EF3",
    x"386042E9",
    x"386026E2",
    x"38600ADF",
    x"385FEEE0",
    x"385FD2E4",
    x"385FB6EB",
    x"385F9AF6",
    x"385F7F04",
    x"385F6316",
    x"385F472B",
    x"385F2B44",
    x"385F0F61",
    x"385EF380",
    x"385ED7A4",
    x"385EBBCB",
    x"385E9FF5",
    x"385E8423",
    x"385E6854",
    x"385E4C88",
    x"385E30C1",
    x"385E14FC",
    x"385DF93B",
    x"385DDD7E",
    x"385DC1C4",
    x"385DA60D",
    x"385D8A5A",
    x"385D6EAB",
    x"385D52FF",
    x"385D3756",
    x"385D1BB1",
    x"385D000F",
    x"385CE471",
    x"385CC8D6",
    x"385CAD3F",
    x"385C91AB",
    x"385C761A",
    x"385C5A8D",
    x"385C3F04",
    x"385C237E",
    x"385C07FB",
    x"385BEC7C",
    x"385BD100",
    x"385BB587",
    x"385B9A12",
    x"385B7EA1",
    x"385B6333",
    x"385B47C8",
    x"385B2C61",
    x"385B10FD",
    x"385AF59C",
    x"385ADA3F",
    x"385ABEE6",
    x"385AA390",
    x"385A883D",
    x"385A6CEE",
    x"385A51A2",
    x"385A3659",
    x"385A1B14",
    x"3859FFD3",
    x"3859E494",
    x"3859C959",
    x"3859AE22",
    x"385992EE",
    x"385977BD",
    x"38595C90",
    x"38594166",
    x"38592640",
    x"38590B1C",
    x"3858EFFD",
    x"3858D4E0",
    x"3858B9C8",
    x"38589EB2",
    x"385883A0",
    x"38586891",
    x"38584D86",
    x"3858327E",
    x"38581779",
    x"3857FC78",
    x"3857E17A",
    x"3857C67F",
    x"3857AB88",
    x"38579095",
    x"385775A4",
    x"38575AB7",
    x"38573FCE",
    x"385724E7",
    x"38570A04",
    x"3856EF25",
    x"3856D449",
    x"3856B970",
    x"38569E9A",
    x"385683C8",
    x"385668F9",
    x"38564E2E",
    x"38563366",
    x"385618A1",
    x"3855FDE0",
    x"3855E321",
    x"3855C867",
    x"3855ADAF",
    x"385592FB",
    x"3855784B",
    x"38555D9D",
    x"385542F3",
    x"3855284C",
    x"38550DA9",
    x"3854F309",
    x"3854D86C",
    x"3854BDD3",
    x"3854A33D",
    x"385488AA",
    x"38546E1B",
    x"3854538F",
    x"38543906",
    x"38541E80",
    x"385403FE",
    x"3853E97F",
    x"3853CF04",
    x"3853B48C",
    x"38539A17",
    x"38537FA5",
    x"38536537",
    x"38534ACC",
    x"38533064",
    x"38531600",
    x"3852FB9F",
    x"3852E141",
    x"3852C6E6",
    x"3852AC8F",
    x"3852923B",
    x"385277EB",
    x"38525D9D",
    x"38524353",
    x"3852290C",
    x"38520EC9",
    x"3851F489",
    x"3851DA4C",
    x"3851C012",
    x"3851A5DC",
    x"38518BA9",
    x"38517179",
    x"3851574C",
    x"38513D23",
    x"385122FD",
    x"385108DA",
    x"3850EEBB",
    x"3850D49F",
    x"3850BA86",
    x"3850A070",
    x"3850865D",
    x"38506C4E",
    x"38505242",
    x"3850383A",
    x"38501E34",
    x"38500432",
    x"384FEA33",
    x"384FD038",
    x"384FB63F",
    x"384F9C4A",
    x"384F8258",
    x"384F6869",
    x"384F4E7E",
    x"384F3496",
    x"384F1AB1",
    x"384F00CF",
    x"384EE6F1",
    x"384ECD15",
    x"384EB33D",
    x"384E9969",
    x"384E7F97",
    x"384E65C9",
    x"384E4BFE",
    x"384E3236",
    x"384E1871",
    x"384DFEB0",
    x"384DE4F1",
    x"384DCB36",
    x"384DB17F",
    x"384D97CA",
    x"384D7E19",
    x"384D646B",
    x"384D4AC0",
    x"384D3118",
    x"384D1773",
    x"384CFDD2",
    x"384CE434",
    x"384CCA99",
    x"384CB101",
    x"384C976D",
    x"384C7DDB",
    x"384C644D",
    x"384C4AC2",
    x"384C313A",
    x"384C17B6",
    x"384BFE35",
    x"384BE4B6",
    x"384BCB3B",
    x"384BB1C4",
    x"384B984F",
    x"384B7EDD",
    x"384B656F",
    x"384B4C04",
    x"384B329C",
    x"384B1937",
    x"384AFFD6",
    x"384AE678",
    x"384ACD1C",
    x"384AB3C4",
    x"384A9A6F",
    x"384A811E",
    x"384A67CF",
    x"384A4E84",
    x"384A353B",
    x"384A1BF6",
    x"384A02B4",
    x"3849E976",
    x"3849D03A",
    x"3849B702",
    x"38499DCC",
    x"3849849A",
    x"38496B6B",
    x"3849523F",
    x"38493917",
    x"38491FF1",
    x"384906CF",
    x"3848EDAF",
    x"3848D493",
    x"3848BB7A",
    x"3848A264",
    x"38488952",
    x"38487042",
    x"38485736",
    x"38483E2C",
    x"38482526",
    x"38480C23",
    x"3847F323",
    x"3847DA26",
    x"3847C12C",
    x"3847A836",
    x"38478F42",
    x"38477652",
    x"38475D65",
    x"3847447B",
    x"38472B94",
    x"384712B0",
    x"3846F9CF",
    x"3846E0F1",
    x"3846C817",
    x"3846AF3F",
    x"3846966B",
    x"38467D9A",
    x"384664CC",
    x"38464C01",
    x"38463339",
    x"38461A74",
    x"384601B2",
    x"3845E8F3",
    x"3845D038",
    x"3845B77F",
    x"38459ECA",
    x"38458618",
    x"38456D68",
    x"384554BC",
    x"38453C13",
    x"3845236D",
    x"38450ACA",
    x"3844F22A",
    x"3844D98E",
    x"3844C0F4",
    x"3844A85D",
    x"38448FCA",
    x"3844773A",
    x"38445EAC",
    x"38444622",
    x"38442D9B",
    x"38441516",
    x"3843FC95",
    x"3843E417",
    x"3843CB9C",
    x"3843B324",
    x"38439AB0",
    x"3843823E",
    x"384369CF",
    x"38435163",
    x"384338FB",
    x"38432095",
    x"38430833",
    x"3842EFD3",
    x"3842D777",
    x"3842BF1D",
    x"3842A6C7",
    x"38428E73",
    x"38427623",
    x"38425DD6",
    x"3842458C",
    x"38422D45",
    x"38421500",
    x"3841FCBF",
    x"3841E481",
    x"3841CC46",
    x"3841B40E",
    x"38419BD9",
    x"384183A7",
    x"38416B78",
    x"3841534C",
    x"38413B23",
    x"384122FE",
    x"38410ADB",
    x"3840F2BB",
    x"3840DA9E",
    x"3840C284",
    x"3840AA6D",
    x"3840925A",
    x"38407A49",
    x"3840623B",
    x"38404A30",
    x"38403228",
    x"38401A24",
    x"38400222",
    x"383FEA23",
    x"383FD227",
    x"383FBA2F",
    x"383FA239",
    x"383F8A46",
    x"383F7256",
    x"383F5A69",
    x"383F4280",
    x"383F2A99",
    x"383F12B5",
    x"383EFAD4",
    x"383EE2F6",
    x"383ECB1B",
    x"383EB343",
    x"383E9B6F",
    x"383E839D",
    x"383E6BCE",
    x"383E5402",
    x"383E3C39",
    x"383E2473",
    x"383E0CB0",
    x"383DF4EF",
    x"383DDD32",
    x"383DC578",
    x"383DADC1",
    x"383D960D",
    x"383D7E5B",
    x"383D66AD",
    x"383D4F02",
    x"383D3759",
    x"383D1FB4",
    x"383D0811",
    x"383CF072",
    x"383CD8D5",
    x"383CC13C",
    x"383CA9A5",
    x"383C9211",
    x"383C7A81",
    x"383C62F3",
    x"383C4B68",
    x"383C33E0",
    x"383C1C5B",
    x"383C04D9",
    x"383BED5A",
    x"383BD5DD",
    x"383BBE64",
    x"383BA6EE",
    x"383B8F7A",
    x"383B780A",
    x"383B609C",
    x"383B4932",
    x"383B31CA",
    x"383B1A65",
    x"383B0303",
    x"383AEBA5",
    x"383AD449",
    x"383ABCEF",
    x"383AA599",
    x"383A8E46",
    x"383A76F6",
    x"383A5FA8",
    x"383A485E",
    x"383A3116",
    x"383A19D2",
    x"383A0290",
    x"3839EB51",
    x"3839D415",
    x"3839BCDC",
    x"3839A5A6",
    x"38398E73",
    x"38397742",
    x"38396015",
    x"383948EA",
    x"383931C2",
    x"38391A9E",
    x"3839037C",
    x"3838EC5D",
    x"3838D541",
    x"3838BE28",
    x"3838A711",
    x"38388FFE",
    x"383878ED",
    x"383861E0",
    x"38384AD5",
    x"383833CD",
    x"38381CC8",
    x"383805C6",
    x"3837EEC6",
    x"3837D7CA",
    x"3837C0D0",
    x"3837A9DA",
    x"383792E6",
    x"38377BF5",
    x"38376507",
    x"38374E1C",
    x"38373733",
    x"3837204E",
    x"3837096B",
    x"3836F28C",
    x"3836DBAF",
    x"3836C4D5",
    x"3836ADFD",
    x"38369729",
    x"38368058",
    x"38366989",
    x"383652BD",
    x"38363BF4",
    x"3836252E",
    x"38360E6B",
    x"3835F7AB",
    x"3835E0ED",
    x"3835CA32",
    x"3835B37B",
    x"38359CC6",
    x"38358613",
    x"38356F64",
    x"383558B8",
    x"3835420E",
    x"38352B67",
    x"383514C3",
    x"3834FE22",
    x"3834E784",
    x"3834D0E8",
    x"3834BA4F",
    x"3834A3B9",
    x"38348D26",
    x"38347696",
    x"38346009",
    x"3834497E",
    x"383432F6",
    x"38341C71",
    x"383405EF",
    x"3833EF70",
    x"3833D8F3",
    x"3833C27A",
    x"3833AC03",
    x"3833958F",
    x"38337F1D",
    x"383368AF",
    x"38335243",
    x"38333BDA",
    x"38332574",
    x"38330F11",
    x"3832F8B0",
    x"3832E253",
    x"3832CBF8",
    x"3832B5A0",
    x"38329F4A",
    x"383288F8",
    x"383272A8",
    x"38325C5B",
    x"38324611",
    x"38322FCA",
    x"38321985",
    x"38320343",
    x"3831ED04",
    x"3831D6C8",
    x"3831C08F",
    x"3831AA58",
    x"38319424",
    x"38317DF3",
    x"383167C5",
    x"38315199",
    x"38313B70",
    x"3831254A",
    x"38310F27",
    x"3830F906",
    x"3830E2E9",
    x"3830CCCE",
    x"3830B6B5",
    x"3830A0A0",
    x"38308A8D",
    x"3830747D",
    x"38305E70",
    x"38304866",
    x"3830325E",
    x"38301C59",
    x"38300657",
    x"382FF058",
    x"382FDA5B",
    x"382FC461",
    x"382FAE6A",
    x"382F9875",
    x"382F8284",
    x"382F6C95",
    x"382F56A9",
    x"382F40BF",
    x"382F2AD8",
    x"382F14F4",
    x"382EFF13",
    x"382EE935",
    x"382ED359",
    x"382EBD80",
    x"382EA7A9",
    x"382E91D6",
    x"382E7C05",
    x"382E6637",
    x"382E506B",
    x"382E3AA3",
    x"382E24DD",
    x"382E0F19",
    x"382DF959",
    x"382DE39B",
    x"382DCDE0",
    x"382DB828",
    x"382DA272",
    x"382D8CBF",
    x"382D770F",
    x"382D6161",
    x"382D4BB6",
    x"382D360E",
    x"382D2069",
    x"382D0AC6",
    x"382CF526",
    x"382CDF89",
    x"382CC9EE",
    x"382CB456",
    x"382C9EC1",
    x"382C892F",
    x"382C739F",
    x"382C5E12",
    x"382C4887",
    x"382C3300",
    x"382C1D7B",
    x"382C07F8",
    x"382BF279",
    x"382BDCFC",
    x"382BC782",
    x"382BB20A",
    x"382B9C95",
    x"382B8723",
    x"382B71B3",
    x"382B5C46",
    x"382B46DC",
    x"382B3175",
    x"382B1C10",
    x"382B06AE",
    x"382AF14E",
    x"382ADBF1",
    x"382AC697",
    x"382AB140",
    x"382A9BEB",
    x"382A8699",
    x"382A7149",
    x"382A5BFC",
    x"382A46B2",
    x"382A316B",
    x"382A1C26",
    x"382A06E4",
    x"3829F1A4",
    x"3829DC67",
    x"3829C72D",
    x"3829B1F5",
    x"38299CC0",
    x"3829878E",
    x"3829725F",
    x"38295D32",
    x"38294807",
    x"382932E0",
    x"38291DBB",
    x"38290898",
    x"3828F378",
    x"3828DE5B",
    x"3828C941",
    x"3828B429",
    x"38289F14",
    x"38288A01",
    x"382874F1",
    x"38285FE4",
    x"38284AD9",
    x"382835D1",
    x"382820CC",
    x"38280BC9",
    x"3827F6C9",
    x"3827E1CB",
    x"3827CCD0",
    x"3827B7D8",
    x"3827A2E3",
    x"38278DEF",
    x"382778FF",
    x"38276411",
    x"38274F26",
    x"38273A3D",
    x"38272557",
    x"38271074",
    x"3826FB93",
    x"3826E6B5",
    x"3826D1DA",
    x"3826BD01",
    x"3826A82A",
    x"38269357",
    x"38267E86",
    x"382669B7",
    x"382654EB",
    x"38264022",
    x"38262B5B",
    x"38261697",
    x"382601D5",
    x"3825ED17",
    x"3825D85A",
    x"3825C3A0",
    x"3825AEE9",
    x"38259A35",
    x"38258583",
    x"382570D3",
    x"38255C27",
    x"3825477C",
    x"382532D5",
    x"38251E30",
    x"3825098D",
    x"3824F4ED",
    x"3824E050",
    x"3824CBB5",
    x"3824B71D",
    x"3824A287",
    x"38248DF4",
    x"38247964",
    x"382464D6",
    x"3824504B",
    x"38243BC2",
    x"3824273C",
    x"382412B8",
    x"3823FE37",
    x"3823E9B9",
    x"3823D53D",
    x"3823C0C3",
    x"3823AC4C",
    x"382397D8",
    x"38238366",
    x"38236EF7",
    x"38235A8B",
    x"38234621",
    x"382331B9",
    x"38231D54",
    x"382308F2",
    x"3822F492",
    x"3822E035",
    x"3822CBDA",
    x"3822B782",
    x"3822A32C",
    x"38228ED9",
    x"38227A88",
    x"3822663A",
    x"382251EF",
    x"38223DA6",
    x"3822295F",
    x"3822151B",
    x"382200DA",
    x"3821EC9B",
    x"3821D85F",
    x"3821C425",
    x"3821AFEE",
    x"38219BB9",
    x"38218787",
    x"38217357",
    x"38215F2A",
    x"38214B00",
    x"382136D7",
    x"382122B2",
    x"38210E8F",
    x"3820FA6E",
    x"3820E650",
    x"3820D235",
    x"3820BE1C",
    x"3820AA05",
    x"382095F1",
    x"382081E0",
    x"38206DD1",
    x"382059C4",
    x"382045BA",
    x"382031B3",
    x"38201DAE",
    x"382009AB",
    x"381FF5AB",
    x"381FE1AE",
    x"381FCDB3",
    x"381FB9BA",
    x"381FA5C4",
    x"381F91D1",
    x"381F7DE0",
    x"381F69F2",
    x"381F5606",
    x"381F421C",
    x"381F2E35",
    x"381F1A50",
    x"381F066E",
    x"381EF28F",
    x"381EDEB2",
    x"381ECAD7",
    x"381EB6FF",
    x"381EA329",
    x"381E8F56",
    x"381E7B86",
    x"381E67B7",
    x"381E53EC",
    x"381E4022",
    x"381E2C5C",
    x"381E1897",
    x"381E04D5",
    x"381DF116",
    x"381DDD59",
    x"381DC99F",
    x"381DB5E7",
    x"381DA231",
    x"381D8E7E",
    x"381D7ACE",
    x"381D6720",
    x"381D5374",
    x"381D3FCB",
    x"381D2C24",
    x"381D1880",
    x"381D04DE",
    x"381CF13E",
    x"381CDDA2",
    x"381CCA07",
    x"381CB66F",
    x"381CA2D9",
    x"381C8F46",
    x"381C7BB6",
    x"381C6827",
    x"381C549C",
    x"381C4112",
    x"381C2D8B",
    x"381C1A07",
    x"381C0685",
    x"381BF305",
    x"381BDF88",
    x"381BCC0D",
    x"381BB895",
    x"381BA51F",
    x"381B91AC",
    x"381B7E3B",
    x"381B6ACC",
    x"381B5760",
    x"381B43F6",
    x"381B308F",
    x"381B1D2A",
    x"381B09C8",
    x"381AF668",
    x"381AE30A",
    x"381ACFAF",
    x"381ABC56",
    x"381AA900",
    x"381A95AC",
    x"381A825A",
    x"381A6F0B",
    x"381A5BBF",
    x"381A4874",
    x"381A352D",
    x"381A21E7",
    x"381A0EA4",
    x"3819FB64",
    x"3819E825",
    x"3819D4E9",
    x"3819C1B0",
    x"3819AE79",
    x"38199B44",
    x"38198812",
    x"381974E2",
    x"381961B5",
    x"38194E8A",
    x"38193B61",
    x"3819283B",
    x"38191517",
    x"381901F6",
    x"3818EED7",
    x"3818DBBA",
    x"3818C8A0",
    x"3818B588",
    x"3818A273",
    x"38188F5F",
    x"38187C4F",
    x"38186940",
    x"38185634",
    x"3818432B",
    x"38183024",
    x"38181D1F",
    x"38180A1C",
    x"3817F71C",
    x"3817E41F",
    x"3817D123",
    x"3817BE2A",
    x"3817AB34",
    x"3817983F",
    x"3817854E",
    x"3817725E",
    x"38175F71",
    x"38174C86",
    x"3817399E",
    x"381726B8",
    x"381713D4",
    x"381700F3",
    x"3816EE14",
    x"3816DB37",
    x"3816C85D",
    x"3816B585",
    x"3816A2B0",
    x"38168FDD",
    x"38167D0C",
    x"38166A3D",
    x"38165771",
    x"381644A7",
    x"381631E0",
    x"38161F1B",
    x"38160C58",
    x"3815F998",
    x"3815E6DA",
    x"3815D41E",
    x"3815C165",
    x"3815AEAE",
    x"38159BF9",
    x"38158947",
    x"38157697",
    x"381563E9",
    x"3815513E",
    x"38153E95",
    x"38152BEE",
    x"3815194A",
    x"381506A8",
    x"3814F408",
    x"3814E16B",
    x"3814CED0",
    x"3814BC37",
    x"3814A9A1",
    x"3814970D",
    x"3814847B",
    x"381471EC",
    x"38145F5F",
    x"38144CD4",
    x"38143A4B",
    x"381427C5",
    x"38141541",
    x"381402C0",
    x"3813F041",
    x"3813DDC4",
    x"3813CB49",
    x"3813B8D1",
    x"3813A65B",
    x"381393E7",
    x"38138176",
    x"38136F07",
    x"38135C9A",
    x"38134A30",
    x"381337C8",
    x"38132562",
    x"381312FE",
    x"3813009D",
    x"3812EE3E",
    x"3812DBE2",
    x"3812C987",
    x"3812B72F",
    x"3812A4DA",
    x"38129286",
    x"38128035",
    x"38126DE6",
    x"38125B99",
    x"3812494F",
    x"38123707",
    x"381224C1",
    x"3812127E",
    x"3812003D",
    x"3811EDFE",
    x"3811DBC1",
    x"3811C987",
    x"3811B74F",
    x"3811A519",
    x"381192E6",
    x"381180B4",
    x"38116E85",
    x"38115C59",
    x"38114A2E",
    x"38113806",
    x"381125E0",
    x"381113BD",
    x"3811019B",
    x"3810EF7C",
    x"3810DD60",
    x"3810CB45",
    x"3810B92D",
    x"3810A717",
    x"38109503",
    x"381082F1",
    x"381070E2",
    x"38105ED5",
    x"38104CCA",
    x"38103AC2",
    x"381028BC",
    x"381016B8",
    x"381004B6",
    x"380FF2B7",
    x"380FE0B9",
    x"380FCEBE",
    x"380FBCC6",
    x"380FAACF",
    x"380F98DB",
    x"380F86E9",
    x"380F74F9",
    x"380F630C",
    x"380F5121",
    x"380F3F38",
    x"380F2D51",
    x"380F1B6C",
    x"380F098A",
    x"380EF7AA",
    x"380EE5CC",
    x"380ED3F0",
    x"380EC217",
    x"380EB040",
    x"380E9E6B",
    x"380E8C98",
    x"380E7AC8",
    x"380E68FA",
    x"380E572E",
    x"380E4564",
    x"380E339C",
    x"380E21D7",
    x"380E1014",
    x"380DFE53",
    x"380DEC94",
    x"380DDAD8",
    x"380DC91D",
    x"380DB765",
    x"380DA5B0",
    x"380D93FC",
    x"380D824B",
    x"380D709B",
    x"380D5EEE",
    x"380D4D44",
    x"380D3B9B",
    x"380D29F5",
    x"380D1851",
    x"380D06AF",
    x"380CF50F",
    x"380CE371",
    x"380CD1D6",
    x"380CC03D",
    x"380CAEA6",
    x"380C9D11",
    x"380C8B7F",
    x"380C79EE",
    x"380C6860",
    x"380C56D4",
    x"380C454B",
    x"380C33C3",
    x"380C223E",
    x"380C10BA",
    x"380BFF39",
    x"380BEDBB",
    x"380BDC3E",
    x"380BCAC4",
    x"380BB94B",
    x"380BA7D5",
    x"380B9661",
    x"380B84F0",
    x"380B7380",
    x"380B6213",
    x"380B50A8",
    x"380B3F3F",
    x"380B2DD8",
    x"380B1C73",
    x"380B0B11",
    x"380AF9B0",
    x"380AE852",
    x"380AD6F6",
    x"380AC59D",
    x"380AB445",
    x"380AA2EF",
    x"380A919C",
    x"380A804B",
    x"380A6EFC",
    x"380A5DAF",
    x"380A4C65",
    x"380A3B1C",
    x"380A29D6",
    x"380A1892",
    x"380A0750",
    x"3809F610",
    x"3809E4D2",
    x"3809D397",
    x"3809C25D",
    x"3809B126",
    x"38099FF1",
    x"38098EBE",
    x"38097D8D",
    x"38096C5F",
    x"38095B32",
    x"38094A08",
    x"380938E0",
    x"380927BA",
    x"38091696",
    x"38090574",
    x"3808F454",
    x"3808E337",
    x"3808D21C",
    x"3808C103",
    x"3808AFEB",
    x"38089ED7",
    x"38088DC4",
    x"38087CB3",
    x"38086BA5",
    x"38085A98",
    x"3808498E",
    x"38083886",
    x"38082780",
    x"3808167C",
    x"3808057A",
    x"3807F47B",
    x"3807E37D",
    x"3807D282",
    x"3807C188",
    x"3807B091",
    x"38079F9C",
    x"38078EA9",
    x"38077DB9",
    x"38076CCA",
    x"38075BDD",
    x"38074AF3",
    x"38073A0B",
    x"38072924",
    x"38071840",
    x"3807075E",
    x"3806F67F",
    x"3806E5A1",
    x"3806D4C5",
    x"3806C3EC",
    x"3806B314",
    x"3806A23F",
    x"3806916C",
    x"3806809A",
    x"38066FCB",
    x"38065EFF",
    x"38064E34",
    x"38063D6B",
    x"38062CA4",
    x"38061BE0",
    x"38060B1D",
    x"3805FA5D",
    x"3805E99F",
    x"3805D8E3",
    x"3805C829",
    x"3805B771",
    x"3805A6BB",
    x"38059607",
    x"38058555",
    x"380574A6",
    x"380563F8",
    x"3805534D",
    x"380542A3",
    x"380531FC",
    x"38052157",
    x"380510B4",
    x"38050013",
    x"3804EF74",
    x"3804DED7",
    x"3804CE3C",
    x"3804BDA3",
    x"3804AD0C",
    x"38049C78",
    x"38048BE5",
    x"38047B55",
    x"38046AC6",
    x"38045A3A",
    x"380449B0",
    x"38043928",
    x"380428A2",
    x"3804181E",
    x"3804079C",
    x"3803F71C",
    x"3803E69E",
    x"3803D622",
    x"3803C5A8",
    x"3803B531",
    x"3803A4BB",
    x"38039447",
    x"380383D6",
    x"38037366",
    x"380362F9",
    x"3803528E",
    x"38034224",
    x"380331BD",
    x"38032158",
    x"380310F5",
    x"38030094",
    x"3802F035",
    x"3802DFD8",
    x"3802CF7D",
    x"3802BF24",
    x"3802AECD",
    x"38029E78",
    x"38028E25",
    x"38027DD5",
    x"38026D86",
    x"38025D39",
    x"38024CEF",
    x"38023CA6",
    x"38022C5F",
    x"38021C1B",
    x"38020BD8",
    x"3801FB98",
    x"3801EB5A",
    x"3801DB1D",
    x"3801CAE3",
    x"3801BAAA",
    x"3801AA74",
    x"38019A40",
    x"38018A0D",
    x"380179DD",
    x"380169AF",
    x"38015983",
    x"38014959",
    x"38013930",
    x"3801290A",
    x"380118E6",
    x"380108C4",
    x"3800F8A4",
    x"3800E886",
    x"3800D86A",
    x"3800C850",
    x"3800B838",
    x"3800A822",
    x"3800980E",
    x"380087FC",
    x"380077EC",
    x"380067DE",
    x"380057D2",
    x"380047C8",
    x"380037C0",
    x"380027BA",
    x"380017B6",
    x"380007B4",
    x"37FFEF68",
    x"37FFCF6C",
    x"37FFAF74",
    x"37FF8F80",
    x"37FF6F90",
    x"37FF4FA4",
    x"37FF2FBC",
    x"37FF0FD8",
    x"37FEEFF8",
    x"37FED01C",
    x"37FEB044",
    x"37FE9070",
    x"37FE70A0",
    x"37FE50D4",
    x"37FE310C",
    x"37FE1148",
    x"37FDF188",
    x"37FDD1CC",
    x"37FDB213",
    x"37FD925F",
    x"37FD72AF",
    x"37FD5302",
    x"37FD335A",
    x"37FD13B6",
    x"37FCF415",
    x"37FCD479",
    x"37FCB4E0",
    x"37FC954B",
    x"37FC75BB",
    x"37FC562E",
    x"37FC36A5",
    x"37FC1720",
    x"37FBF79F",
    x"37FBD822",
    x"37FBB8A9",
    x"37FB9934",
    x"37FB79C3",
    x"37FB5A56",
    x"37FB3AEC",
    x"37FB1B87",
    x"37FAFC25",
    x"37FADCC8",
    x"37FABD6E",
    x"37FA9E19",
    x"37FA7EC7",
    x"37FA5F79",
    x"37FA402F",
    x"37FA20E9",
    x"37FA01A7",
    x"37F9E268",
    x"37F9C32E",
    x"37F9A3F8",
    x"37F984C5",
    x"37F96596",
    x"37F9466C",
    x"37F92745",
    x"37F90822",
    x"37F8E903",
    x"37F8C9E8",
    x"37F8AAD0",
    x"37F88BBD",
    x"37F86CAD",
    x"37F84DA2",
    x"37F82E9A",
    x"37F80F96",
    x"37F7F096",
    x"37F7D19A",
    x"37F7B2A2",
    x"37F793AD",
    x"37F774BD",
    x"37F755D0",
    x"37F736E7",
    x"37F71802",
    x"37F6F921",
    x"37F6DA44",
    x"37F6BB6B",
    x"37F69C95",
    x"37F67DC4",
    x"37F65EF6",
    x"37F6402C",
    x"37F62166",
    x"37F602A3",
    x"37F5E3E5",
    x"37F5C52B",
    x"37F5A674",
    x"37F587C1",
    x"37F56912",
    x"37F54A67",
    x"37F52BBF",
    x"37F50D1C",
    x"37F4EE7C",
    x"37F4CFE0",
    x"37F4B148",
    x"37F492B4",
    x"37F47423",
    x"37F45597",
    x"37F4370E",
    x"37F41889",
    x"37F3FA08",
    x"37F3DB8A",
    x"37F3BD11",
    x"37F39E9B",
    x"37F38029",
    x"37F361BB",
    x"37F34351",
    x"37F324EA",
    x"37F30688",
    x"37F2E829",
    x"37F2C9CE",
    x"37F2AB76",
    x"37F28D23",
    x"37F26ED3",
    x"37F25087",
    x"37F2323F",
    x"37F213FA",
    x"37F1F5BA",
    x"37F1D77D",
    x"37F1B944",
    x"37F19B0F",
    x"37F17CDD",
    x"37F15EAF",
    x"37F14086",
    x"37F1225F",
    x"37F1043D",
    x"37F0E61E",
    x"37F0C803",
    x"37F0A9EC",
    x"37F08BD9",
    x"37F06DC9",
    x"37F04FBD",
    x"37F031B5",
    x"37F013B1",
    x"37EFF5B0",
    x"37EFD7B4",
    x"37EFB9BB",
    x"37EF9BC5",
    x"37EF7DD4",
    x"37EF5FE6",
    x"37EF41FC",
    x"37EF2415",
    x"37EF0633",
    x"37EEE854",
    x"37EECA78",
    x"37EEACA1",
    x"37EE8ECD",
    x"37EE70FD",
    x"37EE5331",
    x"37EE3569",
    x"37EE17A4",
    x"37EDF9E3",
    x"37EDDC25",
    x"37EDBE6C",
    x"37EDA0B6",
    x"37ED8303",
    x"37ED6555",
    x"37ED47AA",
    x"37ED2A03",
    x"37ED0C60",
    x"37ECEEC0",
    x"37ECD124",
    x"37ECB38C",
    x"37EC95F7",
    x"37EC7866",
    x"37EC5AD9",
    x"37EC3D4F",
    x"37EC1FCA",
    x"37EC0247",
    x"37EBE4C9",
    x"37EBC74E",
    x"37EBA9D7",
    x"37EB8C64",
    x"37EB6EF4",
    x"37EB5188",
    x"37EB3420",
    x"37EB16BB",
    x"37EAF95A",
    x"37EADBFD",
    x"37EABEA3",
    x"37EAA14D",
    x"37EA83FB",
    x"37EA66AC",
    x"37EA4961",
    x"37EA2C1A",
    x"37EA0ED6",
    x"37E9F196",
    x"37E9D45A",
    x"37E9B721",
    x"37E999EC",
    x"37E97CBA",
    x"37E95F8D",
    x"37E94263",
    x"37E9253C",
    x"37E90819",
    x"37E8EAFA",
    x"37E8CDDE",
    x"37E8B0C7",
    x"37E893B2",
    x"37E876A2",
    x"37E85995",
    x"37E83C8B",
    x"37E81F85",
    x"37E80283",
    x"37E7E585",
    x"37E7C88A",
    x"37E7AB93",
    x"37E78E9F",
    x"37E771AF",
    x"37E754C3",
    x"37E737DA",
    x"37E71AF5",
    x"37E6FE13",
    x"37E6E135",
    x"37E6C45B",
    x"37E6A784",
    x"37E68AB1",
    x"37E66DE1",
    x"37E65115",
    x"37E6344D",
    x"37E61788",
    x"37E5FAC7",
    x"37E5DE0A",
    x"37E5C150",
    x"37E5A499",
    x"37E587E7",
    x"37E56B37",
    x"37E54E8C",
    x"37E531E4",
    x"37E5153F",
    x"37E4F89E",
    x"37E4DC01",
    x"37E4BF67",
    x"37E4A2D1",
    x"37E4863F",
    x"37E469B0",
    x"37E44D24",
    x"37E4309C",
    x"37E41418",
    x"37E3F797",
    x"37E3DB1A",
    x"37E3BEA1",
    x"37E3A22B",
    x"37E385B8",
    x"37E36949",
    x"37E34CDE",
    x"37E33076",
    x"37E31412",
    x"37E2F7B1",
    x"37E2DB54",
    x"37E2BEFA",
    x"37E2A2A4",
    x"37E28651",
    x"37E26A02",
    x"37E24DB7",
    x"37E2316F",
    x"37E2152B",
    x"37E1F8EA",
    x"37E1DCAC",
    x"37E1C073",
    x"37E1A43C",
    x"37E18809",
    x"37E16BDA",
    x"37E14FAF",
    x"37E13386",
    x"37E11762",
    x"37E0FB40",
    x"37E0DF23",
    x"37E0C309",
    x"37E0A6F2",
    x"37E08ADF",
    x"37E06ECF",
    x"37E052C3",
    x"37E036BB",
    x"37E01AB6",
    x"37DFFEB4",
    x"37DFE2B6",
    x"37DFC6BB",
    x"37DFAAC4",
    x"37DF8ED1",
    x"37DF72E0",
    x"37DF56F4",
    x"37DF3B0B",
    x"37DF1F25",
    x"37DF0343",
    x"37DEE764",
    x"37DECB89",
    x"37DEAFB1",
    x"37DE93DD",
    x"37DE780C",
    x"37DE5C3F",
    x"37DE4075",
    x"37DE24AF",
    x"37DE08EC",
    x"37DDED2D",
    x"37DDD171",
    x"37DDB5B8",
    x"37DD9A03",
    x"37DD7E52",
    x"37DD62A4",
    x"37DD46F9",
    x"37DD2B52",
    x"37DD0FAE",
    x"37DCF40E",
    x"37DCD871",
    x"37DCBCD8",
    x"37DCA142",
    x"37DC85B0",
    x"37DC6A21",
    x"37DC4E95",
    x"37DC330D",
    x"37DC1789",
    x"37DBFC07",
    x"37DBE08A",
    x"37DBC50F",
    x"37DBA998",
    x"37DB8E25",
    x"37DB72B5",
    x"37DB5748",
    x"37DB3BDF",
    x"37DB2079",
    x"37DB0517",
    x"37DAE9B8",
    x"37DACE5C",
    x"37DAB304",
    x"37DA97B0",
    x"37DA7C5E",
    x"37DA6111",
    x"37DA45C6",
    x"37DA2A7F",
    x"37DA0F3B",
    x"37D9F3FB",
    x"37D9D8BE",
    x"37D9BD85",
    x"37D9A24F",
    x"37D9871C",
    x"37D96BED",
    x"37D950C2",
    x"37D93599",
    x"37D91A74",
    x"37D8FF52",
    x"37D8E434",
    x"37D8C919",
    x"37D8AE02",
    x"37D892EE",
    x"37D877DD",
    x"37D85CD0",
    x"37D841C6",
    x"37D826C0",
    x"37D80BBC",
    x"37D7F0BD",
    x"37D7D5C0",
    x"37D7BAC7",
    x"37D79FD1",
    x"37D784DF",
    x"37D769F0",
    x"37D74F05",
    x"37D7341D",
    x"37D71938",
    x"37D6FE56",
    x"37D6E378",
    x"37D6C89D",
    x"37D6ADC6",
    x"37D692F2",
    x"37D67821",
    x"37D65D54",
    x"37D6428A",
    x"37D627C3",
    x"37D60D00",
    x"37D5F240",
    x"37D5D783",
    x"37D5BCCA",
    x"37D5A214",
    x"37D58762",
    x"37D56CB2",
    x"37D55206",
    x"37D5375E",
    x"37D51CB9",
    x"37D50217",
    x"37D4E778",
    x"37D4CCDD",
    x"37D4B245",
    x"37D497B0",
    x"37D47D1F",
    x"37D46291",
    x"37D44806",
    x"37D42D7F",
    x"37D412FB",
    x"37D3F87A",
    x"37D3DDFD",
    x"37D3C383",
    x"37D3A90C",
    x"37D38E98",
    x"37D37428",
    x"37D359BB",
    x"37D33F52",
    x"37D324EC",
    x"37D30A89",
    x"37D2F029",
    x"37D2D5CD",
    x"37D2BB73",
    x"37D2A11E",
    x"37D286CB",
    x"37D26C7C",
    x"37D25230",
    x"37D237E7",
    x"37D21DA2",
    x"37D20360",
    x"37D1E921",
    x"37D1CEE6",
    x"37D1B4AE",
    x"37D19A79",
    x"37D18047",
    x"37D16618",
    x"37D14BED",
    x"37D131C6",
    x"37D117A1",
    x"37D0FD80",
    x"37D0E362",
    x"37D0C947",
    x"37D0AF2F",
    x"37D0951B",
    x"37D07B0A",
    x"37D060FC",
    x"37D046F2",
    x"37D02CEA",
    x"37D012E6",
    x"37CFF8E6",
    x"37CFDEE8",
    x"37CFC4EE",
    x"37CFAAF7",
    x"37CF9103",
    x"37CF7713",
    x"37CF5D26",
    x"37CF433B",
    x"37CF2955",
    x"37CF0F71",
    x"37CEF591",
    x"37CEDBB4",
    x"37CEC1DA",
    x"37CEA803",
    x"37CE8E30",
    x"37CE7460",
    x"37CE5A93",
    x"37CE40C9",
    x"37CE2703",
    x"37CE0D3F",
    x"37CDF37F",
    x"37CDD9C2",
    x"37CDC009",
    x"37CDA652",
    x"37CD8C9F",
    x"37CD72EF",
    x"37CD5943",
    x"37CD3F99",
    x"37CD25F3",
    x"37CD0C50",
    x"37CCF2B0",
    x"37CCD913",
    x"37CCBF79",
    x"37CCA5E3",
    x"37CC8C50",
    x"37CC72C0",
    x"37CC5933",
    x"37CC3FAA",
    x"37CC2623",
    x"37CC0CA0",
    x"37CBF320",
    x"37CBD9A3",
    x"37CBC02A",
    x"37CBA6B3",
    x"37CB8D40",
    x"37CB73D0",
    x"37CB5A63",
    x"37CB40F9",
    x"37CB2793",
    x"37CB0E2F",
    x"37CAF4CF",
    x"37CADB72",
    x"37CAC218",
    x"37CAA8C2",
    x"37CA8F6E",
    x"37CA761E",
    x"37CA5CD1",
    x"37CA4387",
    x"37CA2A40",
    x"37CA10FC",
    x"37C9F7BC",
    x"37C9DE7E",
    x"37C9C544",
    x"37C9AC0D",
    x"37C992D9",
    x"37C979A8",
    x"37C9607A",
    x"37C94750",
    x"37C92E29",
    x"37C91504",
    x"37C8FBE3",
    x"37C8E2C5",
    x"37C8C9AB",
    x"37C8B093",
    x"37C8977F",
    x"37C87E6D",
    x"37C8655F",
    x"37C84C54",
    x"37C8334C",
    x"37C81A47",
    x"37C80145",
    x"37C7E847",
    x"37C7CF4B",
    x"37C7B653",
    x"37C79D5E",
    x"37C7846C",
    x"37C76B7D",
    x"37C75291",
    x"37C739A8",
    x"37C720C2",
    x"37C707E0",
    x"37C6EF00",
    x"37C6D624",
    x"37C6BD4B",
    x"37C6A475",
    x"37C68BA2",
    x"37C672D2",
    x"37C65A05",
    x"37C6413B",
    x"37C62875",
    x"37C60FB1",
    x"37C5F6F1",
    x"37C5DE33",
    x"37C5C579",
    x"37C5ACC2",
    x"37C5940E",
    x"37C57B5D",
    x"37C562AF",
    x"37C54A04",
    x"37C5315D",
    x"37C518B8",
    x"37C50016",
    x"37C4E778",
    x"37C4CEDD",
    x"37C4B644",
    x"37C49DAF",
    x"37C4851D",
    x"37C46C8E",
    x"37C45402",
    x"37C43B79",
    x"37C422F3",
    x"37C40A70",
    x"37C3F1F0",
    x"37C3D973",
    x"37C3C0FA",
    x"37C3A883",
    x"37C39010",
    x"37C3779F",
    x"37C35F32",
    x"37C346C7",
    x"37C32E60",
    x"37C315FC",
    x"37C2FD9B",
    x"37C2E53C",
    x"37C2CCE1",
    x"37C2B489",
    x"37C29C34",
    x"37C283E2",
    x"37C26B93",
    x"37C25347",
    x"37C23AFE",
    x"37C222B9",
    x"37C20A76",
    x"37C1F236",
    x"37C1D9F9",
    x"37C1C1BF",
    x"37C1A989",
    x"37C19155",
    x"37C17924",
    x"37C160F7",
    x"37C148CC",
    x"37C130A5",
    x"37C11880",
    x"37C1005E",
    x"37C0E840",
    x"37C0D024",
    x"37C0B80C",
    x"37C09FF6",
    x"37C087E4",
    x"37C06FD4",
    x"37C057C8",
    x"37C03FBE",
    x"37C027B8",
    x"37C00FB4",
    x"37BFF7B4",
    x"37BFDFB7",
    x"37BFC7BC",
    x"37BFAFC5",
    x"37BF97D0",
    x"37BF7FDF",
    x"37BF67F0",
    x"37BF5005",
    x"37BF381C",
    x"37BF2037",
    x"37BF0854",
    x"37BEF075",
    x"37BED898",
    x"37BEC0BE",
    x"37BEA8E8",
    x"37BE9114",
    x"37BE7944",
    x"37BE6176",
    x"37BE49AB",
    x"37BE31E3",
    x"37BE1A1F",
    x"37BE025D",
    x"37BDEA9E",
    x"37BDD2E2",
    x"37BDBB29",
    x"37BDA373",
    x"37BD8BC1",
    x"37BD7411",
    x"37BD5C64",
    x"37BD44B9",
    x"37BD2D12",
    x"37BD156E",
    x"37BCFDCD",
    x"37BCE62F",
    x"37BCCE93",
    x"37BCB6FB",
    x"37BC9F66",
    x"37BC87D3",
    x"37BC7044",
    x"37BC58B7",
    x"37BC412E",
    x"37BC29A7",
    x"37BC1223",
    x"37BBFAA2",
    x"37BBE324",
    x"37BBCBAA",
    x"37BBB432",
    x"37BB9CBD",
    x"37BB854A",
    x"37BB6DDB",
    x"37BB566F",
    x"37BB3F06",
    x"37BB279F",
    x"37BB103C",
    x"37BAF8DB",
    x"37BAE17D",
    x"37BACA23",
    x"37BAB2CB",
    x"37BA9B76",
    x"37BA8424",
    x"37BA6CD5",
    x"37BA5589",
    x"37BA3E40",
    x"37BA26F9",
    x"37BA0FB6",
    x"37B9F875",
    x"37B9E138",
    x"37B9C9FD",
    x"37B9B2C5",
    x"37B99B90",
    x"37B9845E",
    x"37B96D2F",
    x"37B95603",
    x"37B93EDA",
    x"37B927B3",
    x"37B91090",
    x"37B8F96F",
    x"37B8E251",
    x"37B8CB37",
    x"37B8B41F",
    x"37B89D0A",
    x"37B885F7",
    x"37B86EE8",
    x"37B857DC",
    x"37B840D2",
    x"37B829CB",
    x"37B812C8",
    x"37B7FBC7",
    x"37B7E4C9",
    x"37B7CDCE",
    x"37B7B6D5",
    x"37B79FE0",
    x"37B788ED",
    x"37B771FE",
    x"37B75B11",
    x"37B74427",
    x"37B72D40",
    x"37B7165C",
    x"37B6FF7A",
    x"37B6E89C",
    x"37B6D1C0",
    x"37B6BAE7",
    x"37B6A411",
    x"37B68D3E",
    x"37B6766E",
    x"37B65FA1",
    x"37B648D6",
    x"37B6320E",
    x"37B61B4A",
    x"37B60488",
    x"37B5EDC8",
    x"37B5D70C",
    x"37B5C053",
    x"37B5A99C",
    x"37B592E8",
    x"37B57C37",
    x"37B56589",
    x"37B54EDE",
    x"37B53836",
    x"37B52190",
    x"37B50AED",
    x"37B4F44D",
    x"37B4DDB0",
    x"37B4C716",
    x"37B4B07E",
    x"37B499EA",
    x"37B48358",
    x"37B46CC9",
    x"37B4563D",
    x"37B43FB3",
    x"37B4292D",
    x"37B412A9",
    x"37B3FC28",
    x"37B3E5AA",
    x"37B3CF2F",
    x"37B3B8B6",
    x"37B3A240",
    x"37B38BCE",
    x"37B3755D",
    x"37B35EF0",
    x"37B34886",
    x"37B3321E",
    x"37B31BB9",
    x"37B30557",
    x"37B2EEF8",
    x"37B2D89B",
    x"37B2C242",
    x"37B2ABEB",
    x"37B29597",
    x"37B27F45",
    x"37B268F7",
    x"37B252AB",
    x"37B23C62",
    x"37B2261C",
    x"37B20FD9",
    x"37B1F998",
    x"37B1E35A",
    x"37B1CD1F",
    x"37B1B6E7",
    x"37B1A0B2",
    x"37B18A7F",
    x"37B1744F",
    x"37B15E22",
    x"37B147F7",
    x"37B131D0",
    x"37B11BAB",
    x"37B10589",
    x"37B0EF6A",
    x"37B0D94D",
    x"37B0C333",
    x"37B0AD1C",
    x"37B09708",
    x"37B080F6",
    x"37B06AE8",
    x"37B054DC",
    x"37B03ED3",
    x"37B028CC",
    x"37B012C8",
    x"37AFFCC7",
    x"37AFE6C9",
    x"37AFD0CE",
    x"37AFBAD5",
    x"37AFA4DF",
    x"37AF8EEC",
    x"37AF78FB",
    x"37AF630D",
    x"37AF4D22",
    x"37AF373A",
    x"37AF2155",
    x"37AF0B72",
    x"37AEF592",
    x"37AEDFB4",
    x"37AEC9DA",
    x"37AEB402",
    x"37AE9E2D",
    x"37AE885A",
    x"37AE728B",
    x"37AE5CBE",
    x"37AE46F4",
    x"37AE312C",
    x"37AE1B67",
    x"37AE05A5",
    x"37ADEFE6",
    x"37ADDA29",
    x"37ADC46F",
    x"37ADAEB8",
    x"37AD9904",
    x"37AD8352",
    x"37AD6DA3",
    x"37AD57F6",
    x"37AD424D",
    x"37AD2CA6",
    x"37AD1702",
    x"37AD0160",
    x"37ACEBC1",
    x"37ACD625",
    x"37ACC08C",
    x"37ACAAF5",
    x"37AC9561",
    x"37AC7FD0",
    x"37AC6A41",
    x"37AC54B5",
    x"37AC3F2C",
    x"37AC29A5",
    x"37AC1421",
    x"37ABFEA0",
    x"37ABE922",
    x"37ABD3A6",
    x"37ABBE2D",
    x"37ABA8B6",
    x"37AB9343",
    x"37AB7DD2",
    x"37AB6863",
    x"37AB52F8",
    x"37AB3D8F",
    x"37AB2828",
    x"37AB12C5",
    x"37AAFD64",
    x"37AAE805",
    x"37AAD2A9",
    x"37AABD50",
    x"37AAA7FA",
    x"37AA92A7",
    x"37AA7D56",
    x"37AA6807",
    x"37AA52BB",
    x"37AA3D72",
    x"37AA282C",
    x"37AA12E8",
    x"37A9FDA7",
    x"37A9E869",
    x"37A9D32D",
    x"37A9BDF4",
    x"37A9A8BE",
    x"37A9938A",
    x"37A97E59",
    x"37A9692A",
    x"37A953FF",
    x"37A93ED5",
    x"37A929AF",
    x"37A9148B",
    x"37A8FF6A",
    x"37A8EA4B",
    x"37A8D52F",
    x"37A8C016",
    x"37A8AAFF",
    x"37A895EB",
    x"37A880DA",
    x"37A86BCB",
    x"37A856BF",
    x"37A841B5",
    x"37A82CAE",
    x"37A817AA",
    x"37A802A8",
    x"37A7EDA9",
    x"37A7D8AD",
    x"37A7C3B3",
    x"37A7AEBC",
    x"37A799C8",
    x"37A784D6",
    x"37A76FE6",
    x"37A75AFA",
    x"37A74610",
    x"37A73128",
    x"37A71C43",
    x"37A70761",
    x"37A6F281",
    x"37A6DDA4",
    x"37A6C8CA",
    x"37A6B3F2",
    x"37A69F1D",
    x"37A68A4A",
    x"37A6757A",
    x"37A660AD",
    x"37A64BE2",
    x"37A6371A",
    x"37A62255",
    x"37A60D92",
    x"37A5F8D1",
    x"37A5E413",
    x"37A5CF58",
    x"37A5BAA0",
    x"37A5A5E9",
    x"37A59136",
    x"37A57C85",
    x"37A567D7",
    x"37A5532B",
    x"37A53E82",
    x"37A529DC",
    x"37A51538",
    x"37A50096",
    x"37A4EBF7",
    x"37A4D75B",
    x"37A4C2C2",
    x"37A4AE2B",
    x"37A49996",
    x"37A48504",
    x"37A47075",
    x"37A45BE8",
    x"37A4475E",
    x"37A432D6",
    x"37A41E51",
    x"37A409CF",
    x"37A3F54F",
    x"37A3E0D1",
    x"37A3CC57",
    x"37A3B7DE",
    x"37A3A369",
    x"37A38EF5",
    x"37A37A85",
    x"37A36617",
    x"37A351AB",
    x"37A33D42",
    x"37A328DC",
    x"37A31478",
    x"37A30017",
    x"37A2EBB8",
    x"37A2D75C",
    x"37A2C302",
    x"37A2AEAB",
    x"37A29A57",
    x"37A28605",
    x"37A271B5",
    x"37A25D68",
    x"37A2491E",
    x"37A234D6",
    x"37A22091",
    x"37A20C4E",
    x"37A1F80D",
    x"37A1E3D0",
    x"37A1CF95",
    x"37A1BB5C",
    x"37A1A726",
    x"37A192F2",
    x"37A17EC1",
    x"37A16A92",
    x"37A15666",
    x"37A1423D",
    x"37A12E16",
    x"37A119F1",
    x"37A105CF",
    x"37A0F1B0",
    x"37A0DD93",
    x"37A0C978",
    x"37A0B560",
    x"37A0A14B",
    x"37A08D38",
    x"37A07928",
    x"37A0651A",
    x"37A0510E",
    x"37A03D06",
    x"37A028FF",
    x"37A014FB",
    x"37A000FA",
    x"379FECFB",
    x"379FD8FF",
    x"379FC505",
    x"379FB10D",
    x"379F9D19",
    x"379F8926",
    x"379F7536",
    x"379F6149",
    x"379F4D5E",
    x"379F3976",
    x"379F2590",
    x"379F11AC",
    x"379EFDCB",
    x"379EE9ED",
    x"379ED611",
    x"379EC237",
    x"379EAE60",
    x"379E9A8C",
    x"379E86BA",
    x"379E72EA",
    x"379E5F1D",
    x"379E4B52",
    x"379E378A",
    x"379E23C4",
    x"379E1001",
    x"379DFC40",
    x"379DE882",
    x"379DD4C6",
    x"379DC10D",
    x"379DAD56",
    x"379D99A1",
    x"379D85EF",
    x"379D7240",
    x"379D5E93",
    x"379D4AE8",
    x"379D3740",
    x"379D239A",
    x"379D0FF7",
    x"379CFC56",
    x"379CE8B8",
    x"379CD51C",
    x"379CC183",
    x"379CADEC",
    x"379C9A57",
    x"379C86C5",
    x"379C7336",
    x"379C5FA9",
    x"379C4C1E",
    x"379C3896",
    x"379C2510",
    x"379C118C",
    x"379BFE0B",
    x"379BEA8D",
    x"379BD711",
    x"379BC397",
    x"379BB020",
    x"379B9CAB",
    x"379B8939",
    x"379B75C9",
    x"379B625B",
    x"379B4EF0",
    x"379B3B87",
    x"379B2821",
    x"379B14BD",
    x"379B015C",
    x"379AEDFD",
    x"379ADAA0",
    x"379AC746",
    x"379AB3EF",
    x"379AA099",
    x"379A8D47",
    x"379A79F6",
    x"379A66A8",
    x"379A535C",
    x"379A4013",
    x"379A2CCC",
    x"379A1988",
    x"379A0646",
    x"3799F306",
    x"3799DFC9",
    x"3799CC8E",
    x"3799B956",
    x"3799A620",
    x"379992ED",
    x"37997FBB",
    x"37996C8D",
    x"37995960",
    x"37994636",
    x"3799330F",
    x"37991FEA",
    x"37990CC7",
    x"3798F9A6",
    x"3798E688",
    x"3798D36D",
    x"3798C053",
    x"3798AD3D",
    x"37989A28",
    x"37988716",
    x"37987406",
    x"379860F9",
    x"37984DEE",
    x"37983AE6",
    x"379827DF",
    x"379814DC",
    x"379801DA",
    x"3797EEDB",
    x"3797DBDE",
    x"3797C8E4",
    x"3797B5EC",
    x"3797A2F7",
    x"37979004",
    x"37977D13",
    x"37976A24",
    x"37975738",
    x"3797444E",
    x"37973167",
    x"37971E82",
    x"37970B9F",
    x"3796F8BF",
    x"3796E5E1",
    x"3796D306",
    x"3796C02D",
    x"3796AD56",
    x"37969A81",
    x"379687AF",
    x"379674DF",
    x"37966212",
    x"37964F47",
    x"37963C7E",
    x"379629B8",
    x"379616F4",
    x"37960432",
    x"3795F173",
    x"3795DEB6",
    x"3795CBFB",
    x"3795B943",
    x"3795A68D",
    x"379593D9",
    x"37958128",
    x"37956E79",
    x"37955BCC",
    x"37954922",
    x"3795367A",
    x"379523D4",
    x"37951131",
    x"3794FE90",
    x"3794EBF1",
    x"3794D955",
    x"3794C6BB",
    x"3794B423",
    x"3794A18E",
    x"37948EFB",
    x"37947C6A",
    x"379469DC",
    x"3794574F",
    x"379444C6",
    x"3794323E",
    x"37941FB9",
    x"37940D36",
    x"3793FAB6",
    x"3793E838",
    x"3793D5BC",
    x"3793C342",
    x"3793B0CB",
    x"37939E56",
    x"37938BE3",
    x"37937973",
    x"37936705",
    x"37935499",
    x"37934230",
    x"37932FC9",
    x"37931D64",
    x"37930B01",
    x"3792F8A1",
    x"3792E643",
    x"3792D3E8",
    x"3792C18E",
    x"3792AF37",
    x"37929CE2",
    x"37928A90",
    x"37927840",
    x"379265F2",
    x"379253A6",
    x"3792415D",
    x"37922F16",
    x"37921CD1",
    x"37920A8F",
    x"3791F84F",
    x"3791E611",
    x"3791D3D5",
    x"3791C19C",
    x"3791AF65",
    x"37919D30",
    x"37918AFD",
    x"379178CD",
    x"3791669F",
    x"37915474",
    x"3791424A",
    x"37913023",
    x"37911DFE",
    x"37910BDB",
    x"3790F9BB",
    x"3790E79D",
    x"3790D581",
    x"3790C368",
    x"3790B150",
    x"37909F3B",
    x"37908D29",
    x"37907B18",
    x"3790690A",
    x"379056FE",
    x"379044F4",
    x"379032ED",
    x"379020E7",
    x"37900EE4",
    x"378FFCE4",
    x"378FEAE5",
    x"378FD8E9",
    x"378FC6EF",
    x"378FB4F7",
    x"378FA302",
    x"378F910E",
    x"378F7F1D",
    x"378F6D2F",
    x"378F5B42",
    x"378F4958",
    x"378F3770",
    x"378F258A",
    x"378F13A6",
    x"378F01C5",
    x"378EEFE6",
    x"378EDE09",
    x"378ECC2E",
    x"378EBA56",
    x"378EA880",
    x"378E96AC",
    x"378E84DA",
    x"378E730B",
    x"378E613D",
    x"378E4F72",
    x"378E3DAA",
    x"378E2BE3",
    x"378E1A1F",
    x"378E085C",
    x"378DF69C",
    x"378DE4DF",
    x"378DD323",
    x"378DC16A",
    x"378DAFB3",
    x"378D9DFE",
    x"378D8C4B",
    x"378D7A9B",
    x"378D68ED",
    x"378D5741",
    x"378D4597",
    x"378D33EF",
    x"378D224A",
    x"378D10A7",
    x"378CFF06",
    x"378CED67",
    x"378CDBCA",
    x"378CCA30",
    x"378CB898",
    x"378CA702",
    x"378C956E",
    x"378C83DD",
    x"378C724D",
    x"378C60C0",
    x"378C4F35",
    x"378C3DAC",
    x"378C2C26",
    x"378C1AA1",
    x"378C091F",
    x"378BF79F",
    x"378BE621",
    x"378BD4A5",
    x"378BC32C",
    x"378BB1B5",
    x"378BA03F",
    x"378B8ECC",
    x"378B7D5C",
    x"378B6BED",
    x"378B5A81",
    x"378B4916",
    x"378B37AE",
    x"378B2649",
    x"378B14E5",
    x"378B0383",
    x"378AF224",
    x"378AE0C7",
    x"378ACF6C",
    x"378ABE13",
    x"378AACBC",
    x"378A9B68",
    x"378A8A15",
    x"378A78C5",
    x"378A6777",
    x"378A562B",
    x"378A44E2",
    x"378A339A",
    x"378A2255",
    x"378A1112",
    x"3789FFD1",
    x"3789EE92",
    x"3789DD55",
    x"3789CC1A",
    x"3789BAE2",
    x"3789A9AC",
    x"37899877",
    x"37898745",
    x"37897616",
    x"378964E8",
    x"378953BC",
    x"37894293",
    x"3789316C",
    x"37892047",
    x"37890F24",
    x"3788FE03",
    x"3788ECE4",
    x"3788DBC8",
    x"3788CAAD",
    x"3788B995",
    x"3788A87F",
    x"3788976B",
    x"37888659",
    x"37887549",
    x"3788643C",
    x"37885330",
    x"37884227",
    x"37883120",
    x"3788201B",
    x"37880F18",
    x"3787FE17",
    x"3787ED18",
    x"3787DC1C",
    x"3787CB21",
    x"3787BA29",
    x"3787A933",
    x"3787983E",
    x"3787874C",
    x"3787765D",
    x"3787656F",
    x"37875483",
    x"3787439A",
    x"378732B2",
    x"378721CD",
    x"378710EA",
    x"37870009",
    x"3786EF2A",
    x"3786DE4D",
    x"3786CD72",
    x"3786BC9A",
    x"3786ABC3",
    x"37869AEF",
    x"37868A1C",
    x"3786794C",
    x"3786687E",
    x"378657B2",
    x"378646E8",
    x"37863620",
    x"3786255B",
    x"37861497",
    x"378603D6",
    x"3785F316",
    x"3785E259",
    x"3785D19D",
    x"3785C0E4",
    x"3785B02D",
    x"37859F78",
    x"37858EC5",
    x"37857E15",
    x"37856D66",
    x"37855CB9",
    x"37854C0F",
    x"37853B66",
    x"37852AC0",
    x"37851A1C",
    x"37850979",
    x"3784F8D9",
    x"3784E83B",
    x"3784D79F",
    x"3784C705",
    x"3784B66D",
    x"3784A5D8",
    x"37849544",
    x"378484B2",
    x"37847423",
    x"37846395",
    x"3784530A",
    x"37844280",
    x"378431F9",
    x"37842174",
    x"378410F1",
    x"37840070",
    x"3783EFF1",
    x"3783DF74",
    x"3783CEF9",
    x"3783BE80",
    x"3783AE09",
    x"37839D95",
    x"37838D22",
    x"37837CB1",
    x"37836C43",
    x"37835BD6",
    x"37834B6C",
    x"37833B03",
    x"37832A9D",
    x"37831A39",
    x"378309D6",
    x"3782F976",
    x"3782E918",
    x"3782D8BC",
    x"3782C862",
    x"3782B80A",
    x"3782A7B4",
    x"37829760",
    x"3782870E",
    x"378276BE",
    x"37826670",
    x"37825625",
    x"378245DB",
    x"37823593",
    x"3782254D",
    x"3782150A",
    x"378204C8",
    x"3781F489",
    x"3781E44B",
    x"3781D40F",
    x"3781C3D6",
    x"3781B39F",
    x"3781A369",
    x"37819336",
    x"37818304",
    x"378172D5",
    x"378162A8",
    x"3781527C",
    x"37814253",
    x"3781322C",
    x"37812206",
    x"378111E3",
    x"378101C2",
    x"3780F1A3",
    x"3780E186",
    x"3780D16A",
    x"3780C151",
    x"3780B13A",
    x"3780A125",
    x"37809112",
    x"37808101",
    x"378070F1",
    x"378060E4",
    x"378050D9",
    x"378040D0",
    x"378030C9",
    x"378020C4",
    x"378010C1",
    x"378000C0",
    x"377FE181",
    x"377FC187",
    x"377FA191",
    x"377F819F",
    x"377F61B1",
    x"377F41C6",
    x"377F21E0",
    x"377F01FE",
    x"377EE220",
    x"377EC245",
    x"377EA26F",
    x"377E829D",
    x"377E62CE",
    x"377E4304",
    x"377E233E",
    x"377E037B",
    x"377DE3BD",
    x"377DC402",
    x"377DA44C",
    x"377D8499",
    x"377D64EB",
    x"377D4540",
    x"377D2599",
    x"377D05F7",
    x"377CE658",
    x"377CC6BD",
    x"377CA726",
    x"377C8793",
    x"377C6804",
    x"377C4879",
    x"377C28F2",
    x"377C096F",
    x"377BE9F0",
    x"377BCA74",
    x"377BAAFD",
    x"377B8B8A",
    x"377B6C1A",
    x"377B4CAF",
    x"377B2D47",
    x"377B0DE3",
    x"377AEE84",
    x"377ACF28",
    x"377AAFD0",
    x"377A907C",
    x"377A712C",
    x"377A51DF",
    x"377A3297",
    x"377A1353",
    x"3779F412",
    x"3779D4D6",
    x"3779B59D",
    x"37799668",
    x"37797738",
    x"3779580B",
    x"377938E2",
    x"377919BC",
    x"3778FA9B",
    x"3778DB7E",
    x"3778BC64",
    x"37789D4F",
    x"37787E3D",
    x"37785F2F",
    x"37784025",
    x"3778211F",
    x"3778021D",
    x"3777E31E",
    x"3777C424",
    x"3777A52D",
    x"3777863B",
    x"3777674C",
    x"37774861",
    x"3777297A",
    x"37770A97",
    x"3776EBB7",
    x"3776CCDC",
    x"3776AE04",
    x"37768F30",
    x"37767060",
    x"37765194",
    x"377632CC",
    x"37761407",
    x"3775F547",
    x"3775D68A",
    x"3775B7D1",
    x"3775991C",
    x"37757A6B",
    x"37755BBD",
    x"37753D14",
    x"37751E6E",
    x"3774FFCC",
    x"3774E12E",
    x"3774C294",
    x"3774A3FE",
    x"3774856B",
    x"377466DC",
    x"37744851",
    x"377429CA",
    x"37740B47",
    x"3773ECC7",
    x"3773CE4C",
    x"3773AFD4",
    x"37739160",
    x"377372EF",
    x"37735483",
    x"3773361A",
    x"377317B5",
    x"3772F954",
    x"3772DAF7",
    x"3772BC9E",
    x"37729E48",
    x"37727FF6",
    x"377261A8",
    x"3772435E",
    x"37722517",
    x"377206D4",
    x"3771E895",
    x"3771CA5A",
    x"3771AC23",
    x"37718DEF",
    x"37716FBF",
    x"37715193",
    x"3771336B",
    x"37711546",
    x"3770F726",
    x"3770D909",
    x"3770BAEF",
    x"37709CDA",
    x"37707EC8",
    x"377060BA",
    x"377042B0",
    x"377024A9",
    x"377006A7",
    x"376FE8A8",
    x"376FCAAD",
    x"376FACB5",
    x"376F8EC1",
    x"376F70D1",
    x"376F52E5",
    x"376F34FD",
    x"376F1718",
    x"376EF937",
    x"376EDB5A",
    x"376EBD80",
    x"376E9FAA",
    x"376E81D8",
    x"376E640A",
    x"376E463F",
    x"376E2878",
    x"376E0AB5",
    x"376DECF6",
    x"376DCF3A",
    x"376DB182",
    x"376D93CD",
    x"376D761D",
    x"376D5870",
    x"376D3AC7",
    x"376D1D21",
    x"376CFF7F",
    x"376CE1E1",
    x"376CC447",
    x"376CA6B0",
    x"376C891D",
    x"376C6B8E",
    x"376C4E02",
    x"376C307B",
    x"376C12F6",
    x"376BF576",
    x"376BD7F9",
    x"376BBA80",
    x"376B9D0A",
    x"376B7F99",
    x"376B622A",
    x"376B44C0",
    x"376B2759",
    x"376B09F6",
    x"376AEC97",
    x"376ACF3B",
    x"376AB1E3",
    x"376A948F",
    x"376A773E",
    x"376A59F1",
    x"376A3CA7",
    x"376A1F62",
    x"376A021F",
    x"3769E4E1",
    x"3769C7A6",
    x"3769AA6F",
    x"37698D3C",
    x"3769700C",
    x"376952E0",
    x"376935B7",
    x"37691892",
    x"3768FB71",
    x"3768DE53",
    x"3768C139",
    x"3768A423",
    x"37688710",
    x"37686A01",
    x"37684CF6",
    x"37682FEE",
    x"376812EA",
    x"3767F5E9",
    x"3767D8EC",
    x"3767BBF3",
    x"37679EFD",
    x"3767820B",
    x"3767651D",
    x"37674832",
    x"37672B4B",
    x"37670E67",
    x"3766F187",
    x"3766D4AB",
    x"3766B7D2",
    x"37669AFD",
    x"37667E2B",
    x"3766615D",
    x"37664493",
    x"376627CC",
    x"37660B09",
    x"3765EE49",
    x"3765D18D",
    x"3765B4D5",
    x"37659820",
    x"37657B6F",
    x"37655EC1",
    x"37654217",
    x"37652571",
    x"376508CE",
    x"3764EC2F",
    x"3764CF93",
    x"3764B2FB",
    x"37649666",
    x"376479D5",
    x"37645D48",
    x"376440BE",
    x"37642438",
    x"376407B5",
    x"3763EB36",
    x"3763CEBA",
    x"3763B242",
    x"376395CD",
    x"3763795C",
    x"37635CEF",
    x"37634085",
    x"3763241F",
    x"376307BC",
    x"3762EB5D",
    x"3762CF01",
    x"3762B2A9",
    x"37629655",
    x"37627A04",
    x"37625DB6",
    x"3762416C",
    x"37622526",
    x"376208E3",
    x"3761ECA4",
    x"3761D068",
    x"3761B42F",
    x"376197FB",
    x"37617BC9",
    x"37615F9C",
    x"37614372",
    x"3761274B",
    x"37610B28",
    x"3760EF08",
    x"3760D2EC",
    x"3760B6D3",
    x"37609ABE",
    x"37607EAD",
    x"3760629F",
    x"37604694",
    x"37602A8D",
    x"37600E89",
    x"375FF289",
    x"375FD68D",
    x"375FBA94",
    x"375F9E9E",
    x"375F82AC",
    x"375F66BD",
    x"375F4AD2",
    x"375F2EEB",
    x"375F1307",
    x"375EF726",
    x"375EDB49",
    x"375EBF6F",
    x"375EA399",
    x"375E87C6",
    x"375E6BF7",
    x"375E502B",
    x"375E3463",
    x"375E189E",
    x"375DFCDD",
    x"375DE11F",
    x"375DC565",
    x"375DA9AE",
    x"375D8DFA",
    x"375D724A",
    x"375D569E",
    x"375D3AF4",
    x"375D1F4F",
    x"375D03AD",
    x"375CE80E",
    x"375CCC73",
    x"375CB0DB",
    x"375C9546",
    x"375C79B5",
    x"375C5E28",
    x"375C429E",
    x"375C2717",
    x"375C0B94",
    x"375BF014",
    x"375BD498",
    x"375BB91F",
    x"375B9DAA",
    x"375B8238",
    x"375B66C9",
    x"375B4B5E",
    x"375B2FF6",
    x"375B1492",
    x"375AF931",
    x"375ADDD4",
    x"375AC27A",
    x"375AA723",
    x"375A8BD0",
    x"375A7080",
    x"375A5534",
    x"375A39EB",
    x"375A1EA5",
    x"375A0363",
    x"3759E825",
    x"3759CCE9",
    x"3759B1B1",
    x"3759967D",
    x"37597B4C",
    x"3759601E",
    x"375944F4",
    x"375929CD",
    x"37590EA9",
    x"3758F389",
    x"3758D86C",
    x"3758BD53",
    x"3758A23D",
    x"3758872A",
    x"37586C1B",
    x"3758510F",
    x"37583607",
    x"37581B02",
    x"37580000",
    x"3757E502",
    x"3757CA07",
    x"3757AF0F",
    x"3757941B",
    x"3757792A",
    x"37575E3D",
    x"37574353",
    x"3757286C",
    x"37570D89",
    x"3756F2A9",
    x"3756D7CC",
    x"3756BCF3",
    x"3756A21D",
    x"3756874A",
    x"37566C7B",
    x"375651AF",
    x"375636E7",
    x"37561C21",
    x"37560160",
    x"3755E6A1",
    x"3755CBE6",
    x"3755B12E",
    x"3755967A",
    x"37557BC8",
    x"3755611B",
    x"37554670",
    x"37552BC9",
    x"37551125",
    x"3754F685",
    x"3754DBE8",
    x"3754C14E",
    x"3754A6B7",
    x"37548C24",
    x"37547194",
    x"37545708",
    x"37543C7F",
    x"375421F9",
    x"37540776",
    x"3753ECF7",
    x"3753D27B",
    x"3753B802",
    x"37539D8D",
    x"3753831B",
    x"375368AC",
    x"37534E41",
    x"375333D8",
    x"37531974",
    x"3752FF12",
    x"3752E4B4",
    x"3752CA59",
    x"3752B001",
    x"375295AD",
    x"37527B5C",
    x"3752610E",
    x"375246C4",
    x"37522C7C",
    x"37521238",
    x"3751F7F8",
    x"3751DDBA",
    x"3751C380",
    x"3751A94A",
    x"37518F16",
    x"375174E6",
    x"37515AB9",
    x"3751408F",
    x"37512669",
    x"37510C46",
    x"3750F226",
    x"3750D809",
    x"3750BDF0",
    x"3750A3D9",
    x"375089C7",
    x"37506FB7",
    x"375055AB",
    x"37503BA2",
    x"3750219C",
    x"37500799",
    x"374FED9A",
    x"374FD39E",
    x"374FB9A5",
    x"374F9FAF",
    x"374F85BD",
    x"374F6BCE",
    x"374F51E2",
    x"374F37FA",
    x"374F1E14",
    x"374F0432",
    x"374EEA53",
    x"374ED077",
    x"374EB69F",
    x"374E9CCA",
    x"374E82F8",
    x"374E6929",
    x"374E4F5D",
    x"374E3595",
    x"374E1BD0",
    x"374E020E",
    x"374DE850",
    x"374DCE94",
    x"374DB4DC",
    x"374D9B27",
    x"374D8175",
    x"374D67C7",
    x"374D4E1B",
    x"374D3473",
    x"374D1ACE",
    x"374D012C",
    x"374CE78E",
    x"374CCDF2",
    x"374CB45A",
    x"374C9AC5",
    x"374C8134",
    x"374C67A5",
    x"374C4E1A",
    x"374C3492",
    x"374C1B0D",
    x"374C018B",
    x"374BE80C",
    x"374BCE91",
    x"374BB519",
    x"374B9BA3",
    x"374B8232",
    x"374B68C3",
    x"374B4F57",
    x"374B35EF",
    x"374B1C8A",
    x"374B0328",
    x"374AE9C9",
    x"374AD06E",
    x"374AB715",
    x"374A9DC0",
    x"374A846E",
    x"374A6B1F",
    x"374A51D3",
    x"374A388A",
    x"374A1F45",
    x"374A0602",
    x"3749ECC3",
    x"3749D387",
    x"3749BA4E",
    x"3749A119",
    x"374987E6",
    x"37496EB7",
    x"3749558A",
    x"37493C61",
    x"3749233B",
    x"37490A18",
    x"3748F0F9",
    x"3748D7DC",
    x"3748BEC3",
    x"3748A5AC",
    x"37488C99",
    x"37487389",
    x"37485A7C",
    x"37484173",
    x"3748286C",
    x"37480F69",
    x"3747F668",
    x"3747DD6B",
    x"3747C471",
    x"3747AB7A",
    x"37479286",
    x"37477995",
    x"374760A8",
    x"374747BD",
    x"37472ED6",
    x"374715F1",
    x"3746FD10",
    x"3746E432",
    x"3746CB57",
    x"3746B27F",
    x"374699AB",
    x"374680D9",
    x"3746680A",
    x"37464F3F",
    x"37463677",
    x"37461DB1",
    x"374604EF",
    x"3745EC30",
    x"3745D374",
    x"3745BABB",
    x"3745A205",
    x"37458953",
    x"374570A3",
    x"374557F6",
    x"37453F4D",
    x"374526A7",
    x"37450E03",
    x"3744F563",
    x"3744DCC6",
    x"3744C42C",
    x"3744AB95",
    x"37449301",
    x"37447A70",
    x"374461E2",
    x"37444958",
    x"374430D0",
    x"3744184C",
    x"3743FFCA",
    x"3743E74C",
    x"3743CED0",
    x"3743B658",
    x"37439DE3",
    x"37438570",
    x"37436D01",
    x"37435495",
    x"37433C2C",
    x"374323C6",
    x"37430B63",
    x"3742F303",
    x"3742DAA6",
    x"3742C24D",
    x"3742A9F6",
    x"374291A2",
    x"37427951",
    x"37426104",
    x"374248B9",
    x"37423072",
    x"3742182D",
    x"3741FFEC",
    x"3741E7AD",
    x"3741CF72",
    x"3741B739",
    x"37419F04",
    x"374186D1",
    x"37416EA2",
    x"37415676",
    x"37413E4D",
    x"37412626",
    x"37410E03",
    x"3740F5E3",
    x"3740DDC6",
    x"3740C5AB",
    x"3740AD94",
    x"37409580",
    x"37407D6F",
    x"37406561",
    x"37404D55",
    x"3740354D",
    x"37401D48",
    x"37400546",
    x"373FED47",
    x"373FD54B",
    x"373FBD51",
    x"373FA55B",
    x"373F8D68",
    x"373F7578",
    x"373F5D8B",
    x"373F45A1",
    x"373F2DB9",
    x"373F15D5",
    x"373EFDF4",
    x"373EE616",
    x"373ECE3A",
    x"373EB662",
    x"373E9E8D",
    x"373E86BA",
    x"373E6EEB",
    x"373E571F",
    x"373E3F55",
    x"373E278F",
    x"373E0FCB",
    x"373DF80B",
    x"373DE04D",
    x"373DC893",
    x"373DB0DB",
    x"373D9927",
    x"373D8175",
    x"373D69C6",
    x"373D521A",
    x"373D3A72",
    x"373D22CC",
    x"373D0B29",
    x"373CF389",
    x"373CDBEC",
    x"373CC452",
    x"373CACBB",
    x"373C9527",
    x"373C7D96",
    x"373C6608",
    x"373C4E7C",
    x"373C36F4",
    x"373C1F6E",
    x"373C07EC",
    x"373BF06D",
    x"373BD8F0",
    x"373BC176",
    x"373BAA00",
    x"373B928C",
    x"373B7B1B",
    x"373B63AD",
    x"373B4C42",
    x"373B34DA",
    x"373B1D75",
    x"373B0613",
    x"373AEEB3",
    x"373AD757",
    x"373ABFFD",
    x"373AA8A7",
    x"373A9153",
    x"373A7A03",
    x"373A62B5",
    x"373A4B6A",
    x"373A3422",
    x"373A1CDD",
    x"373A059B",
    x"3739EE5B",
    x"3739D71F",
    x"3739BFE6",
    x"3739A8AF",
    x"3739917C",
    x"37397A4B",
    x"3739631D",
    x"37394BF2",
    x"373934CA",
    x"37391DA5",
    x"37390683",
    x"3738EF63",
    x"3738D847",
    x"3738C12D",
    x"3738AA16",
    x"37389303",
    x"37387BF2",
    x"373864E4",
    x"37384DD8",
    x"373836D0",
    x"37381FCB",
    x"373808C8",
    x"3737F1C9",
    x"3737DACC",
    x"3737C3D2",
    x"3737ACDB",
    x"373795E7",
    x"37377EF5",
    x"37376807",
    x"3737511B",
    x"37373A33",
    x"3737234D",
    x"37370C6A",
    x"3736F58A",
    x"3736DEAC",
    x"3736C7D2",
    x"3736B0FA",
    x"37369A26",
    x"37368354",
    x"37366C85",
    x"373655B9",
    x"37363EEF",
    x"37362829",
    x"37361165",
    x"3735FAA5",
    x"3735E3E7",
    x"3735CD2C",
    x"3735B673",
    x"37359FBE",
    x"3735890C",
    x"3735725C",
    x"37355BAF",
    x"37354505",
    x"37352E5E",
    x"373517B9",
    x"37350118",
    x"3734EA79",
    x"3734D3DD",
    x"3734BD44",
    x"3734A6AE",
    x"3734901A",
    x"3734798A",
    x"373462FC",
    x"37344C71",
    x"373435E9",
    x"37341F64",
    x"373408E1",
    x"3733F261",
    x"3733DBE4",
    x"3733C56A",
    x"3733AEF3",
    x"3733987F",
    x"3733820D",
    x"37336B9E",
    x"37335532",
    x"37333EC9",
    x"37332862",
    x"373311FF",
    x"3732FB9E",
    x"3732E540",
    x"3732CEE5",
    x"3732B88C",
    x"3732A236",
    x"37328BE4",
    x"37327593",
    x"37325F46",
    x"373248FC",
    x"373232B4",
    x"37321C6F",
    x"3732062D",
    x"3731EFED",
    x"3731D9B1",
    x"3731C377",
    x"3731AD40",
    x"3731970C",
    x"373180DA",
    x"37316AAB",
    x"37315480",
    x"37313E56",
    x"37312830",
    x"3731120C",
    x"3730FBEB",
    x"3730E5CD",
    x"3730CFB2",
    x"3730B999",
    x"3730A384",
    x"37308D71",
    x"37307760",
    x"37306153",
    x"37304B48",
    x"37303540",
    x"37301F3B",
    x"37300938",
    x"372FF338",
    x"372FDD3B",
    x"372FC741",
    x"372FB149",
    x"372F9B55",
    x"372F8563",
    x"372F6F73",
    x"372F5987",
    x"372F439D",
    x"372F2DB6",
    x"372F17D1",
    x"372F01F0",
    x"372EEC11",
    x"372ED635",
    x"372EC05B",
    x"372EAA85",
    x"372E94B1",
    x"372E7EE0",
    x"372E6911",
    x"372E5345",
    x"372E3D7C",
    x"372E27B6",
    x"372E11F2",
    x"372DFC31",
    x"372DE673",
    x"372DD0B8",
    x"372DBAFF",
    x"372DA549",
    x"372D8F96",
    x"372D79E5",
    x"372D6437",
    x"372D4E8C",
    x"372D38E4",
    x"372D233E",
    x"372D0D9B",
    x"372CF7FB",
    x"372CE25D",
    x"372CCCC2",
    x"372CB72A",
    x"372CA194",
    x"372C8C01",
    x"372C7671",
    x"372C60E4",
    x"372C4B59",
    x"372C35D1",
    x"372C204B",
    x"372C0AC9",
    x"372BF549",
    x"372BDFCB",
    x"372BCA51",
    x"372BB4D9",
    x"372B9F64",
    x"372B89F1",
    x"372B7481",
    x"372B5F14",
    x"372B49A9",
    x"372B3441",
    x"372B1EDC",
    x"372B097A",
    x"372AF41A",
    x"372ADEBD",
    x"372AC962",
    x"372AB40A",
    x"372A9EB5",
    x"372A8963",
    x"372A7413",
    x"372A5EC6",
    x"372A497B",
    x"372A3433",
    x"372A1EEE",
    x"372A09AC",
    x"3729F46C",
    x"3729DF2E",
    x"3729C9F4",
    x"3729B4BC",
    x"37299F87",
    x"37298A54",
    x"37297524",
    x"37295FF7",
    x"37294ACC",
    x"372935A4",
    x"3729207F",
    x"37290B5C",
    x"3728F63C",
    x"3728E11E",
    x"3728CC04",
    x"3728B6EB",
    x"3728A1D6",
    x"37288CC3",
    x"372877B3",
    x"372862A5",
    x"37284D9A",
    x"37283892",
    x"3728238C",
    x"37280E89",
    x"3727F988",
    x"3727E48A",
    x"3727CF8F",
    x"3727BA96",
    x"3727A5A0",
    x"372790AD",
    x"37277BBC",
    x"372766CE",
    x"372751E3",
    x"37273CFA",
    x"37272813",
    x"37271330",
    x"3726FE4F",
    x"3726E970",
    x"3726D494",
    x"3726BFBB",
    x"3726AAE4",
    x"37269610",
    x"3726813F",
    x"37266C70",
    x"372657A4",
    x"372642DA",
    x"37262E13",
    x"3726194E",
    x"3726048D",
    x"3725EFCD",
    x"3725DB11",
    x"3725C657",
    x"3725B19F",
    x"37259CEA",
    x"37258838",
    x"37257388",
    x"37255EDB",
    x"37254A30",
    x"37253588",
    x"372520E3",
    x"37250C40",
    x"3724F7A0",
    x"3724E302",
    x"3724CE67",
    x"3724B9CF",
    x"3724A539",
    x"372490A5",
    x"37247C15",
    x"37246786",
    x"372452FB",
    x"37243E72",
    x"372429EB",
    x"37241567",
    x"372400E6",
    x"3723EC67",
    x"3723D7EB",
    x"3723C371",
    x"3723AEFA",
    x"37239A85",
    x"37238613",
    x"372371A4",
    x"37235D37",
    x"372348CC",
    x"37233465",
    x"37231FFF",
    x"37230B9D",
    x"3722F73C",
    x"3722E2DF",
    x"3722CE84",
    x"3722BA2B",
    x"3722A5D5",
    x"37229182",
    x"37227D31",
    x"372268E2",
    x"37225496",
    x"3722404D",
    x"37222C06",
    x"372217C2",
    x"37220380",
    x"3721EF41",
    x"3721DB05",
    x"3721C6CB",
    x"3721B293",
    x"37219E5E",
    x"37218A2B",
    x"372175FB",
    x"372161CE",
    x"37214DA3",
    x"3721397A",
    x"37212555",
    x"37211131",
    x"3720FD10",
    x"3720E8F2",
    x"3720D4D6",
    x"3720C0BD",
    x"3720ACA6",
    x"37209891",
    x"37208480",
    x"37207070",
    x"37205C64",
    x"37204859",
    x"37203451",
    x"3720204C",
    x"37200C49",
    x"371FF849",
    x"371FE44B",
    x"371FD050",
    x"371FBC57",
    x"371FA861",
    x"371F946D",
    x"371F807C",
    x"371F6C8D",
    x"371F58A1",
    x"371F44B7",
    x"371F30D0",
    x"371F1CEB",
    x"371F0908",
    x"371EF528",
    x"371EE14B",
    x"371ECD70",
    x"371EB998",
    x"371EA5C2",
    x"371E91EE",
    x"371E7E1D",
    x"371E6A4F",
    x"371E5683",
    x"371E42B9",
    x"371E2EF2",
    x"371E1B2D",
    x"371E076B",
    x"371DF3AB",
    x"371DDFEE",
    x"371DCC33",
    x"371DB87B",
    x"371DA4C5",
    x"371D9112",
    x"371D7D61",
    x"371D69B3",
    x"371D5607",
    x"371D425D",
    x"371D2EB6",
    x"371D1B11",
    x"371D076F",
    x"371CF3D0",
    x"371CE032",
    x"371CCC98",
    x"371CB8FF",
    x"371CA569",
    x"371C91D6",
    x"371C7E45",
    x"371C6AB6",
    x"371C572A",
    x"371C43A1",
    x"371C3019",
    x"371C1C94",
    x"371C0912",
    x"371BF592",
    x"371BE215",
    x"371BCE9A",
    x"371BBB21",
    x"371BA7AB",
    x"371B9437",
    x"371B80C6",
    x"371B6D57",
    x"371B59EB",
    x"371B4680",
    x"371B3319",
    x"371B1FB4",
    x"371B0C51",
    x"371AF8F1",
    x"371AE593",
    x"371AD237",
    x"371ABEDE",
    x"371AAB88",
    x"371A9833",
    x"371A84E1",
    x"371A7192",
    x"371A5E45",
    x"371A4AFB",
    x"371A37B2",
    x"371A246D",
    x"371A1129",
    x"3719FDE8",
    x"3719EAAA",
    x"3719D76E",
    x"3719C434",
    x"3719B0FD",
    x"37199DC8",
    x"37198A95",
    x"37197765",
    x"37196437",
    x"3719510C",
    x"37193DE3",
    x"37192ABC",
    x"37191798",
    x"37190477",
    x"3718F157",
    x"3718DE3A",
    x"3718CB20",
    x"3718B807",
    x"3718A4F2",
    x"371891DE",
    x"37187ECD",
    x"37186BBF",
    x"371858B2",
    x"371845A8",
    x"371832A1",
    x"37181F9C",
    x"37180C99",
    x"3717F999",
    x"3717E69B",
    x"3717D39F",
    x"3717C0A6",
    x"3717ADAF",
    x"37179ABA",
    x"371787C8",
    x"371774D8",
    x"371761EB",
    x"37174F00",
    x"37173C17",
    x"37172931",
    x"3717164D",
    x"3717036B",
    x"3716F08C",
    x"3716DDAF",
    x"3716CAD5",
    x"3716B7FC",
    x"3716A527",
    x"37169253",
    x"37167F82",
    x"37166CB3",
    x"371659E7",
    x"3716471D",
    x"37163455",
    x"37162190",
    x"37160ECD",
    x"3715FC0C",
    x"3715E94E",
    x"3715D692",
    x"3715C3D8",
    x"3715B121",
    x"37159E6C",
    x"37158BB9",
    x"37157909",
    x"3715665B",
    x"371553AF",
    x"37154106",
    x"37152E5F",
    x"37151BBA",
    x"37150918",
    x"3714F678",
    x"3714E3DA",
    x"3714D13F",
    x"3714BEA6",
    x"3714AC0F",
    x"3714997B",
    x"371486E9",
    x"37147459",
    x"371461CC",
    x"37144F41",
    x"37143CB8",
    x"37142A32",
    x"371417AE",
    x"3714052C",
    x"3713F2AC",
    x"3713E02F",
    x"3713CDB4",
    x"3713BB3C",
    x"3713A8C5",
    x"37139651",
    x"371383E0",
    x"37137170",
    x"37135F03",
    x"37134C99",
    x"37133A30",
    x"371327CA",
    x"37131566",
    x"37130305",
    x"3712F0A6",
    x"3712DE49",
    x"3712CBEE",
    x"3712B996",
    x"3712A740",
    x"371294EC",
    x"3712829A",
    x"3712704B",
    x"37125DFE",
    x"37124BB4",
    x"3712396B",
    x"37122725",
    x"371214E2",
    x"371202A0",
    x"3711F061",
    x"3711DE24",
    x"3711CBE9",
    x"3711B9B1",
    x"3711A77B",
    x"37119547",
    x"37118316",
    x"371170E6",
    x"37115EB9",
    x"37114C8F",
    x"37113A66",
    x"37112840",
    x"3711161C",
    x"371103FB",
    x"3710F1DB",
    x"3710DFBE",
    x"3710CDA3",
    x"3710BB8B",
    x"3710A974",
    x"37109760",
    x"3710854F",
    x"3710733F",
    x"37106132",
    x"37104F27",
    x"37103D1E",
    x"37102B17",
    x"37101913",
    x"37100711",
    x"370FF511",
    x"370FE314",
    x"370FD119",
    x"370FBF20",
    x"370FAD29",
    x"370F9B34",
    x"370F8942",
    x"370F7752",
    x"370F6564",
    x"370F5379",
    x"370F418F",
    x"370F2FA8",
    x"370F1DC3",
    x"370F0BE1",
    x"370EFA00",
    x"370EE822",
    x"370ED646",
    x"370EC46D",
    x"370EB295",
    x"370EA0C0",
    x"370E8EED",
    x"370E7D1C",
    x"370E6B4E",
    x"370E5982",
    x"370E47B8",
    x"370E35F0",
    x"370E242A",
    x"370E1267",
    x"370E00A5",
    x"370DEEE6",
    x"370DDD2A",
    x"370DCB6F",
    x"370DB9B7",
    x"370DA801",
    x"370D964D",
    x"370D849B",
    x"370D72EC",
    x"370D613E",
    x"370D4F93",
    x"370D3DEB",
    x"370D2C44",
    x"370D1A9F",
    x"370D08FD",
    x"370CF75D",
    x"370CE5BF",
    x"370CD424",
    x"370CC28A",
    x"370CB0F3",
    x"370C9F5E",
    x"370C8DCB",
    x"370C7C3B",
    x"370C6AAC",
    x"370C5920",
    x"370C4796",
    x"370C360E",
    x"370C2488",
    x"370C1305",
    x"370C0184",
    x"370BF005",
    x"370BDE88",
    x"370BCD0D",
    x"370BBB94",
    x"370BAA1E",
    x"370B98AA",
    x"370B8738",
    x"370B75C8",
    x"370B645A",
    x"370B52EF",
    x"370B4186",
    x"370B301F",
    x"370B1EBA",
    x"370B0D57",
    x"370AFBF6",
    x"370AEA98",
    x"370AD93C",
    x"370AC7E2",
    x"370AB68A",
    x"370AA534",
    x"370A93E0",
    x"370A828F",
    x"370A7140",
    x"370A5FF3",
    x"370A4EA8",
    x"370A3D5F",
    x"370A2C18",
    x"370A1AD4",
    x"370A0992",
    x"3709F852",
    x"3709E714",
    x"3709D5D8",
    x"3709C49E",
    x"3709B367",
    x"3709A231",
    x"370990FE",
    x"37097FCD",
    x"37096E9E",
    x"37095D71",
    x"37094C47",
    x"37093B1E",
    x"370929F8",
    x"370918D4",
    x"370907B2",
    x"3708F692",
    x"3708E574",
    x"3708D459",
    x"3708C33F",
    x"3708B228",
    x"3708A113",
    x"37089000",
    x"37087EEF",
    x"37086DE0",
    x"37085CD3",
    x"37084BC9",
    x"37083AC0",
    x"370829BA",
    x"370818B6",
    x"370807B4",
    x"3707F6B4",
    x"3707E5B6",
    x"3707D4BA",
    x"3707C3C1",
    x"3707B2C9",
    x"3707A1D4",
    x"370790E1",
    x"37077FF0",
    x"37076F01",
    x"37075E14",
    x"37074D2A",
    x"37073C41",
    x"37072B5A",
    x"37071A76",
    x"37070994",
    x"3706F8B4",
    x"3706E7D6",
    x"3706D6FA",
    x"3706C620",
    x"3706B548",
    x"3706A473",
    x"3706939F",
    x"370682CE",
    x"370671FE",
    x"37066131",
    x"37065066",
    x"37063F9D",
    x"37062ED6",
    x"37061E11",
    x"37060D4F",
    x"3705FC8E",
    x"3705EBD0",
    x"3705DB13",
    x"3705CA59",
    x"3705B9A0",
    x"3705A8EA",
    x"37059836",
    x"37058784",
    x"370576D4",
    x"37056627",
    x"3705557B",
    x"370544D1",
    x"3705342A",
    x"37052384",
    x"370512E1",
    x"3705023F",
    x"3704F1A0",
    x"3704E103",
    x"3704D068",
    x"3704BFCF",
    x"3704AF38",
    x"37049EA3",
    x"37048E10",
    x"37047D80",
    x"37046CF1",
    x"37045C64",
    x"37044BDA",
    x"37043B51",
    x"37042ACB",
    x"37041A47",
    x"370409C4",
    x"3703F944",
    x"3703E8C6",
    x"3703D84A",
    x"3703C7D0",
    x"3703B758",
    x"3703A6E2",
    x"3703966E",
    x"370385FD",
    x"3703758D",
    x"3703651F",
    x"370354B4",
    x"3703444A",
    x"370333E3",
    x"3703237D",
    x"3703131A",
    x"370302B8",
    x"3702F259",
    x"3702E1FC",
    x"3702D1A1",
    x"3702C147",
    x"3702B0F0",
    x"3702A09B",
    x"37029048",
    x"37027FF7",
    x"37026FA8",
    x"37025F5B",
    x"37024F10",
    x"37023EC7",
    x"37022E81",
    x"37021E3C",
    x"37020DF9",
    x"3701FDB8",
    x"3701ED7A",
    x"3701DD3D",
    x"3701CD02",
    x"3701BCCA",
    x"3701AC93",
    x"37019C5E",
    x"37018C2C",
    x"37017BFB",
    x"37016BCD",
    x"37015BA0",
    x"37014B76",
    x"37013B4E",
    x"37012B27",
    x"37011B03",
    x"37010AE0",
    x"3700FAC0",
    x"3700EAA2",
    x"3700DA85",
    x"3700CA6B",
    x"3700BA53",
    x"3700AA3D",
    x"37009A28",
    x"37008A16",
    x"37007A06",
    x"370069F7",
    x"370059EB",
    x"370049E1",
    x"370039D9",
    x"370029D3",
    x"370019CE",
    x"370009CC",
    x"36FFF398",
    x"36FFD39B",
    x"36FFB3A3",
    x"36FF93AE",
    x"36FF73BE",
    x"36FF53D1",
    x"36FF33E9",
    x"36FF1404",
    x"36FEF424",
    x"36FED447",
    x"36FEB46F",
    x"36FE949A",
    x"36FE74CA",
    x"36FE54FD",
    x"36FE3535",
    x"36FE1570",
    x"36FDF5AF",
    x"36FDD5F2",
    x"36FDB63A",
    x"36FD9685",
    x"36FD76D4",
    x"36FD5727",
    x"36FD377E",
    x"36FD17D9",
    x"36FCF838",
    x"36FCD89B",
    x"36FCB902",
    x"36FC996D",
    x"36FC79DC",
    x"36FC5A4F",
    x"36FC3AC5",
    x"36FC1B40",
    x"36FBFBBE",
    x"36FBDC41",
    x"36FBBCC7",
    x"36FB9D52",
    x"36FB7DE0",
    x"36FB5E72",
    x"36FB3F08",
    x"36FB1FA2",
    x"36FB0040",
    x"36FAE0E2",
    x"36FAC188",
    x"36FAA232",
    x"36FA82E0",
    x"36FA6391",
    x"36FA4447",
    x"36FA2500",
    x"36FA05BE",
    x"36F9E67F",
    x"36F9C744",
    x"36F9A80D",
    x"36F988DA",
    x"36F969AB",
    x"36F94A7F",
    x"36F92B58",
    x"36F90C35",
    x"36F8ED15",
    x"36F8CDF9",
    x"36F8AEE2",
    x"36F88FCE",
    x"36F870BE",
    x"36F851B1",
    x"36F832A9",
    x"36F813A5",
    x"36F7F4A4",
    x"36F7D5A8",
    x"36F7B6AF",
    x"36F797BA",
    x"36F778C9",
    x"36F759DC",
    x"36F73AF2",
    x"36F71C0D",
    x"36F6FD2B",
    x"36F6DE4E",
    x"36F6BF74",
    x"36F6A09E",
    x"36F681CC",
    x"36F662FD",
    x"36F64433",
    x"36F6256C",
    x"36F606AA",
    x"36F5E7EB",
    x"36F5C930",
    x"36F5AA78",
    x"36F58BC5",
    x"36F56D15",
    x"36F54E6A",
    x"36F52FC2",
    x"36F5111E",
    x"36F4F27E",
    x"36F4D3E1",
    x"36F4B549",
    x"36F496B4",
    x"36F47823",
    x"36F45996",
    x"36F43B0D",
    x"36F41C87",
    x"36F3FE05",
    x"36F3DF88",
    x"36F3C10E",
    x"36F3A297",
    x"36F38425",
    x"36F365B6",
    x"36F3474B",
    x"36F328E4",
    x"36F30A81",
    x"36F2EC22",
    x"36F2CDC6",
    x"36F2AF6E",
    x"36F2911A",
    x"36F272CA",
    x"36F2547E",
    x"36F23635",
    x"36F217F0",
    x"36F1F9AF",
    x"36F1DB72",
    x"36F1BD38",
    x"36F19F02",
    x"36F180D0",
    x"36F162A2",
    x"36F14478",
    x"36F12651",
    x"36F1082E",
    x"36F0EA0F",
    x"36F0CBF4",
    x"36F0ADDC",
    x"36F08FC8",
    x"36F071B8",
    x"36F053AC",
    x"36F035A3",
    x"36F0179E",
    x"36EFF99D",
    x"36EFDBA0",
    x"36EFBDA6",
    x"36EF9FB1",
    x"36EF81BE",
    x"36EF63D0",
    x"36EF45E5",
    x"36EF27FF",
    x"36EF0A1B",
    x"36EEEC3C",
    x"36EECE60",
    x"36EEB088",
    x"36EE92B4",
    x"36EE74E4",
    x"36EE5717",
    x"36EE394E",
    x"36EE1B89",
    x"36EDFDC7",
    x"36EDE009",
    x"36EDC24F",
    x"36EDA499",
    x"36ED86E6",
    x"36ED6937",
    x"36ED4B8C",
    x"36ED2DE4",
    x"36ED1040",
    x"36ECF2A0",
    x"36ECD504",
    x"36ECB76B",
    x"36EC99D6",
    x"36EC7C44",
    x"36EC5EB7",
    x"36EC412D",
    x"36EC23A6",
    x"36EC0624",
    x"36EBE8A5",
    x"36EBCB2A",
    x"36EBADB2",
    x"36EB903E",
    x"36EB72CE",
    x"36EB5561",
    x"36EB37F9",
    x"36EB1A93",
    x"36EAFD32",
    x"36EADFD4",
    x"36EAC27A",
    x"36EAA524",
    x"36EA87D1",
    x"36EA6A82",
    x"36EA4D36",
    x"36EA2FEE",
    x"36EA12AA",
    x"36E9F56A",
    x"36E9D82D",
    x"36E9BAF4",
    x"36E99DBE",
    x"36E9808C",
    x"36E9635E",
    x"36E94633",
    x"36E9290C",
    x"36E90BE9",
    x"36E8EEC9",
    x"36E8D1AD",
    x"36E8B495",
    x"36E89780",
    x"36E87A6F",
    x"36E85D62",
    x"36E84058",
    x"36E82351",
    x"36E8064F",
    x"36E7E950",
    x"36E7CC55",
    x"36E7AF5D",
    x"36E79269",
    x"36E77578",
    x"36E7588B",
    x"36E73BA2",
    x"36E71EBC",
    x"36E701DA",
    x"36E6E4FC",
    x"36E6C821",
    x"36E6AB4A",
    x"36E68E76",
    x"36E671A6",
    x"36E654DA",
    x"36E63811",
    x"36E61B4C",
    x"36E5FE8A",
    x"36E5E1CC",
    x"36E5C512",
    x"36E5A85B",
    x"36E58BA8",
    x"36E56EF8",
    x"36E5524C",
    x"36E535A3",
    x"36E518FF",
    x"36E4FC5D",
    x"36E4DFBF",
    x"36E4C325",
    x"36E4A68F",
    x"36E489FC",
    x"36E46D6C",
    x"36E450E0",
    x"36E43458",
    x"36E417D3",
    x"36E3FB52",
    x"36E3DED4",
    x"36E3C25A",
    x"36E3A5E4",
    x"36E38971",
    x"36E36D01",
    x"36E35096",
    x"36E3342D",
    x"36E317C9",
    x"36E2FB67",
    x"36E2DF0A",
    x"36E2C2B0",
    x"36E2A659",
    x"36E28A06",
    x"36E26DB7",
    x"36E2516B",
    x"36E23522",
    x"36E218DD",
    x"36E1FC9C",
    x"36E1E05E",
    x"36E1C424",
    x"36E1A7ED",
    x"36E18BBA",
    x"36E16F8A",
    x"36E1535E",
    x"36E13735",
    x"36E11B10",
    x"36E0FEEF",
    x"36E0E2D0",
    x"36E0C6B6",
    x"36E0AA9F",
    x"36E08E8B",
    x"36E0727B",
    x"36E0566F",
    x"36E03A66",
    x"36E01E60",
    x"36E0025E",
    x"36DFE65F",
    x"36DFCA64",
    x"36DFAE6D",
    x"36DF9279",
    x"36DF7688",
    x"36DF5A9B",
    x"36DF3EB2",
    x"36DF22CB",
    x"36DF06E9",
    x"36DEEB0A",
    x"36DECF2E",
    x"36DEB356",
    x"36DE9781",
    x"36DE7BB0",
    x"36DE5FE2",
    x"36DE4418",
    x"36DE2851",
    x"36DE0C8E",
    x"36DDF0CE",
    x"36DDD512",
    x"36DDB959",
    x"36DD9DA3",
    x"36DD81F1",
    x"36DD6643",
    x"36DD4A98",
    x"36DD2EF0",
    x"36DD134C",
    x"36DCF7AB",
    x"36DCDC0E",
    x"36DCC074",
    x"36DCA4DE",
    x"36DC894B",
    x"36DC6DBC",
    x"36DC5230",
    x"36DC36A7",
    x"36DC1B22",
    x"36DBFFA0",
    x"36DBE422",
    x"36DBC8A7",
    x"36DBAD30",
    x"36DB91BC",
    x"36DB764C",
    x"36DB5ADF",
    x"36DB3F75",
    x"36DB240F",
    x"36DB08AC",
    x"36DAED4D",
    x"36DAD1F1",
    x"36DAB698",
    x"36DA9B43",
    x"36DA7FF1",
    x"36DA64A3",
    x"36DA4958",
    x"36DA2E11",
    x"36DA12CD",
    x"36D9F78C",
    x"36D9DC4F",
    x"36D9C115",
    x"36D9A5DE",
    x"36D98AAB",
    x"36D96F7C",
    x"36D9544F",
    x"36D93927",
    x"36D91E01",
    x"36D902DF",
    x"36D8E7C0",
    x"36D8CCA5",
    x"36D8B18D",
    x"36D89679",
    x"36D87B68",
    x"36D8605A",
    x"36D84550",
    x"36D82A49",
    x"36D80F45",
    x"36D7F445",
    x"36D7D948",
    x"36D7BE4E",
    x"36D7A358",
    x"36D78866",
    x"36D76D76",
    x"36D7528A",
    x"36D737A2",
    x"36D71CBC",
    x"36D701DA",
    x"36D6E6FC",
    x"36D6CC21",
    x"36D6B149",
    x"36D69674",
    x"36D67BA3",
    x"36D660D5",
    x"36D6460B",
    x"36D62B44",
    x"36D61080",
    x"36D5F5C0",
    x"36D5DB03",
    x"36D5C049",
    x"36D5A593",
    x"36D58AE0",
    x"36D57030",
    x"36D55584",
    x"36D53ADB",
    x"36D52035",
    x"36D50593",
    x"36D4EAF4",
    x"36D4D058",
    x"36D4B5BF",
    x"36D49B2A",
    x"36D48099",
    x"36D4660A",
    x"36D44B7F",
    x"36D430F7",
    x"36D41673",
    x"36D3FBF2",
    x"36D3E174",
    x"36D3C6F9",
    x"36D3AC82",
    x"36D3920E",
    x"36D3779E",
    x"36D35D30",
    x"36D342C6",
    x"36D32860",
    x"36D30DFC",
    x"36D2F39C",
    x"36D2D93F",
    x"36D2BEE6",
    x"36D2A490",
    x"36D28A3D",
    x"36D26FED",
    x"36D255A1",
    x"36D23B58",
    x"36D22112",
    x"36D206CF",
    x"36D1EC90",
    x"36D1D254",
    x"36D1B81C",
    x"36D19DE6",
    x"36D183B4",
    x"36D16985",
    x"36D14F5A",
    x"36D13531",
    x"36D11B0C",
    x"36D100EB",
    x"36D0E6CC",
    x"36D0CCB1",
    x"36D0B299",
    x"36D09884",
    x"36D07E73",
    x"36D06465",
    x"36D04A5A",
    x"36D03052",
    x"36D0164E",
    x"36CFFC4D",
    x"36CFE24F",
    x"36CFC854",
    x"36CFAE5D",
    x"36CF9468",
    x"36CF7A78",
    x"36CF608A",
    x"36CF469F",
    x"36CF2CB8",
    x"36CF12D4",
    x"36CEF8F3",
    x"36CEDF16",
    x"36CEC53C",
    x"36CEAB65",
    x"36CE9191",
    x"36CE77C0",
    x"36CE5DF3",
    x"36CE4429",
    x"36CE2A62",
    x"36CE109E",
    x"36CDF6DE",
    x"36CDDD20",
    x"36CDC366",
    x"36CDA9B0",
    x"36CD8FFC",
    x"36CD764C",
    x"36CD5C9E",
    x"36CD42F4",
    x"36CD294E",
    x"36CD0FAA",
    x"36CCF60A",
    x"36CCDC6D",
    x"36CCC2D3",
    x"36CCA93C",
    x"36CC8FA8",
    x"36CC7618",
    x"36CC5C8B",
    x"36CC4301",
    x"36CC297A",
    x"36CC0FF6",
    x"36CBF676",
    x"36CBDCF9",
    x"36CBC37F",
    x"36CBAA08",
    x"36CB9094",
    x"36CB7724",
    x"36CB5DB7",
    x"36CB444C",
    x"36CB2AE5",
    x"36CB1182",
    x"36CAF821",
    x"36CADEC4",
    x"36CAC569",
    x"36CAAC12",
    x"36CA92BE",
    x"36CA796E",
    x"36CA6020",
    x"36CA46D6",
    x"36CA2D8E",
    x"36CA144A",
    x"36C9FB09",
    x"36C9E1CB",
    x"36C9C891",
    x"36C9AF59",
    x"36C99625",
    x"36C97CF4",
    x"36C963C6",
    x"36C94A9B",
    x"36C93173",
    x"36C9184E",
    x"36C8FF2D",
    x"36C8E60F",
    x"36C8CCF3",
    x"36C8B3DB",
    x"36C89AC7",
    x"36C881B5",
    x"36C868A6",
    x"36C84F9B",
    x"36C83692",
    x"36C81D8D",
    x"36C8048B",
    x"36C7EB8C",
    x"36C7D290",
    x"36C7B997",
    x"36C7A0A2",
    x"36C787AF",
    x"36C76EC0",
    x"36C755D3",
    x"36C73CEA",
    x"36C72404",
    x"36C70B21",
    x"36C6F241",
    x"36C6D965",
    x"36C6C08B",
    x"36C6A7B4",
    x"36C68EE1",
    x"36C67611",
    x"36C65D43",
    x"36C64479",
    x"36C62BB2",
    x"36C612EE",
    x"36C5FA2E",
    x"36C5E170",
    x"36C5C8B5",
    x"36C5AFFE",
    x"36C59749",
    x"36C57E98",
    x"36C565EA",
    x"36C54D3E",
    x"36C53496",
    x"36C51BF1",
    x"36C5034F",
    x"36C4EAB0",
    x"36C4D215",
    x"36C4B97C",
    x"36C4A0E6",
    x"36C48854",
    x"36C46FC4",
    x"36C45738",
    x"36C43EAE",
    x"36C42628",
    x"36C40DA5",
    x"36C3F525",
    x"36C3DCA8",
    x"36C3C42E",
    x"36C3ABB7",
    x"36C39343",
    x"36C37AD2",
    x"36C36264",
    x"36C349F9",
    x"36C33191",
    x"36C3192D",
    x"36C300CB",
    x"36C2E86D",
    x"36C2D011",
    x"36C2B7B9",
    x"36C29F63",
    x"36C28711",
    x"36C26EC1",
    x"36C25675",
    x"36C23E2C",
    x"36C225E5",
    x"36C20DA2",
    x"36C1F562",
    x"36C1DD25",
    x"36C1C4EB",
    x"36C1ACB4",
    x"36C19480",
    x"36C17C4F",
    x"36C16420",
    x"36C14BF5",
    x"36C133CD",
    x"36C11BA9",
    x"36C10387",
    x"36C0EB68",
    x"36C0D34C",
    x"36C0BB33",
    x"36C0A31D",
    x"36C08B0A",
    x"36C072FA",
    x"36C05AED",
    x"36C042E3",
    x"36C02ADD",
    x"36C012D9",
    x"36BFFAD8",
    x"36BFE2DA",
    x"36BFCADF",
    x"36BFB2E7",
    x"36BF9AF2",
    x"36BF8301",
    x"36BF6B12",
    x"36BF5326",
    x"36BF3B3D",
    x"36BF2357",
    x"36BF0B74",
    x"36BEF394",
    x"36BEDBB7",
    x"36BEC3DD",
    x"36BEAC06",
    x"36BE9432",
    x"36BE7C61",
    x"36BE6493",
    x"36BE4CC8",
    x"36BE3500",
    x"36BE1D3B",
    x"36BE0579",
    x"36BDEDB9",
    x"36BDD5FD",
    x"36BDBE44",
    x"36BDA68E",
    x"36BD8EDA",
    x"36BD772A",
    x"36BD5F7C",
    x"36BD47D2",
    x"36BD302A",
    x"36BD1886",
    x"36BD00E4",
    x"36BCE946",
    x"36BCD1AA",
    x"36BCBA11",
    x"36BCA27C",
    x"36BC8AE9",
    x"36BC7359",
    x"36BC5BCC",
    x"36BC4442",
    x"36BC2CBB",
    x"36BC1537",
    x"36BBFDB5",
    x"36BBE637",
    x"36BBCEBC",
    x"36BBB744",
    x"36BB9FCE",
    x"36BB885C",
    x"36BB70EC",
    x"36BB597F",
    x"36BB4216",
    x"36BB2AAF",
    x"36BB134B",
    x"36BAFBEA",
    x"36BAE48C",
    x"36BACD31",
    x"36BAB5D9",
    x"36BA9E83",
    x"36BA8731",
    x"36BA6FE2",
    x"36BA5895",
    x"36BA414B",
    x"36BA2A05",
    x"36BA12C1",
    x"36B9FB80",
    x"36B9E442",
    x"36B9CD07",
    x"36B9B5CF",
    x"36B99E9A",
    x"36B98767",
    x"36B97038",
    x"36B9590B",
    x"36B941E1",
    x"36B92ABB",
    x"36B91397",
    x"36B8FC76",
    x"36B8E558",
    x"36B8CE3C",
    x"36B8B724",
    x"36B8A00F",
    x"36B888FC",
    x"36B871EC",
    x"36B85AE0",
    x"36B843D6",
    x"36B82CCF",
    x"36B815CA",
    x"36B7FEC9",
    x"36B7E7CB",
    x"36B7D0CF",
    x"36B7B9D7",
    x"36B7A2E1",
    x"36B78BEE",
    x"36B774FE",
    x"36B75E11",
    x"36B74726",
    x"36B7303F",
    x"36B7195A",
    x"36B70278",
    x"36B6EB9A",
    x"36B6D4BE",
    x"36B6BDE4",
    x"36B6A70E",
    x"36B6903B",
    x"36B6796A",
    x"36B6629C",
    x"36B64BD1",
    x"36B63509",
    x"36B61E44",
    x"36B60782",
    x"36B5F0C2",
    x"36B5DA06",
    x"36B5C34C",
    x"36B5AC95",
    x"36B595E1",
    x"36B57F2F",
    x"36B56881",
    x"36B551D5",
    x"36B53B2C",
    x"36B52486",
    x"36B50DE3",
    x"36B4F743",
    x"36B4E0A5",
    x"36B4CA0B",
    x"36B4B373",
    x"36B49CDE",
    x"36B4864C",
    x"36B46FBC",
    x"36B45930",
    x"36B442A6",
    x"36B42C1F",
    x"36B4159B",
    x"36B3FF1A",
    x"36B3E89B",
    x"36B3D220",
    x"36B3BBA7",
    x"36B3A531",
    x"36B38EBD",
    x"36B3784D",
    x"36B361DF",
    x"36B34B74",
    x"36B3350C",
    x"36B31EA7",
    x"36B30845",
    x"36B2F1E5",
    x"36B2DB88",
    x"36B2C52E",
    x"36B2AED7",
    x"36B29883",
    x"36B28231",
    x"36B26BE2",
    x"36B25596",
    x"36B23F4D",
    x"36B22906",
    x"36B212C2",
    x"36B1FC81",
    x"36B1E643",
    x"36B1D008",
    x"36B1B9CF",
    x"36B1A399",
    x"36B18D66",
    x"36B17736",
    x"36B16109",
    x"36B14ADE",
    x"36B134B6",
    x"36B11E91",
    x"36B1086E",
    x"36B0F24E",
    x"36B0DC32",
    x"36B0C617",
    x"36B0B000",
    x"36B099EB",
    x"36B083DA",
    x"36B06DCA",
    x"36B057BE",
    x"36B041B5",
    x"36B02BAE",
    x"36B015AA",
    x"36AFFFA8",
    x"36AFE9AA",
    x"36AFD3AE",
    x"36AFBDB5",
    x"36AFA7BE",
    x"36AF91CB",
    x"36AF7BDA",
    x"36AF65EC",
    x"36AF5000",
    x"36AF3A18",
    x"36AF2432",
    x"36AF0E4F",
    x"36AEF86E",
    x"36AEE291",
    x"36AECCB6",
    x"36AEB6DE",
    x"36AEA108",
    x"36AE8B35",
    x"36AE7565",
    x"36AE5F98",
    x"36AE49CD",
    x"36AE3405",
    x"36AE1E40",
    x"36AE087E",
    x"36ADF2BE",
    x"36ADDD01",
    x"36ADC747",
    x"36ADB18F",
    x"36AD9BDB",
    x"36AD8628",
    x"36AD7079",
    x"36AD5ACC",
    x"36AD4522",
    x"36AD2F7B",
    x"36AD19D6",
    x"36AD0435",
    x"36ACEE95",
    x"36ACD8F9",
    x"36ACC35F",
    x"36ACADC8",
    x"36AC9834",
    x"36AC82A2",
    x"36AC6D13",
    x"36AC5787",
    x"36AC41FD",
    x"36AC2C76",
    x"36AC16F2",
    x"36AC0171",
    x"36ABEBF2",
    x"36ABD676",
    x"36ABC0FC",
    x"36ABAB85",
    x"36AB9611",
    x"36AB80A0",
    x"36AB6B31",
    x"36AB55C5",
    x"36AB405C",
    x"36AB2AF5",
    x"36AB1591",
    x"36AB0030",
    x"36AAEAD1",
    x"36AAD575",
    x"36AAC01B",
    x"36AAAAC5",
    x"36AA9571",
    x"36AA801F",
    x"36AA6AD1",
    x"36AA5585",
    x"36AA403B",
    x"36AA2AF5",
    x"36AA15B1",
    x"36AA006F",
    x"36A9EB30",
    x"36A9D5F4",
    x"36A9C0BB",
    x"36A9AB84",
    x"36A99650",
    x"36A9811F",
    x"36A96BF0",
    x"36A956C4",
    x"36A9419A",
    x"36A92C73",
    x"36A9174F",
    x"36A9022D",
    x"36A8ED0E",
    x"36A8D7F2",
    x"36A8C2D9",
    x"36A8ADC1",
    x"36A898AD",
    x"36A8839B",
    x"36A86E8C",
    x"36A85980",
    x"36A84476",
    x"36A82F6F",
    x"36A81A6A",
    x"36A80568",
    x"36A7F069",
    x"36A7DB6C",
    x"36A7C672",
    x"36A7B17A",
    x"36A79C85",
    x"36A78793",
    x"36A772A3",
    x"36A75DB6",
    x"36A748CC",
    x"36A733E4",
    x"36A71EFF",
    x"36A70A1C",
    x"36A6F53D",
    x"36A6E05F",
    x"36A6CB84",
    x"36A6B6AC",
    x"36A6A1D7",
    x"36A68D04",
    x"36A67834",
    x"36A66366",
    x"36A64E9B",
    x"36A639D2",
    x"36A6250C",
    x"36A61049",
    x"36A5FB88",
    x"36A5E6CA",
    x"36A5D20E",
    x"36A5BD55",
    x"36A5A89F",
    x"36A593EB",
    x"36A57F3A",
    x"36A56A8C",
    x"36A555DF",
    x"36A54136",
    x"36A52C8F",
    x"36A517EB",
    x"36A50349",
    x"36A4EEAA",
    x"36A4DA0E",
    x"36A4C574",
    x"36A4B0DC",
    x"36A49C47",
    x"36A487B5",
    x"36A47325",
    x"36A45E98",
    x"36A44A0E",
    x"36A43586",
    x"36A42100",
    x"36A40C7E",
    x"36A3F7FD",
    x"36A3E380",
    x"36A3CF04",
    x"36A3BA8C",
    x"36A3A616",
    x"36A391A2",
    x"36A37D31",
    x"36A368C3",
    x"36A35457",
    x"36A33FEE",
    x"36A32B87",
    x"36A31723",
    x"36A302C1",
    x"36A2EE62",
    x"36A2DA06",
    x"36A2C5AC",
    x"36A2B154",
    x"36A29CFF",
    x"36A288AD",
    x"36A2745D",
    x"36A26010",
    x"36A24BC5",
    x"36A2377D",
    x"36A22337",
    x"36A20EF4",
    x"36A1FAB4",
    x"36A1E676",
    x"36A1D23A",
    x"36A1BE01",
    x"36A1A9CB",
    x"36A19597",
    x"36A18165",
    x"36A16D36",
    x"36A1590A",
    x"36A144E0",
    x"36A130B9",
    x"36A11C94",
    x"36A10872",
    x"36A0F452",
    x"36A0E034",
    x"36A0CC1A",
    x"36A0B801",
    x"36A0A3EC",
    x"36A08FD8",
    x"36A07BC8",
    x"36A067B9",
    x"36A053AE",
    x"36A03FA5",
    x"36A02B9E",
    x"36A0179A",
    x"36A00398",
    x"369FEF99",
    x"369FDB9C",
    x"369FC7A2",
    x"369FB3AA",
    x"369F9FB5",
    x"369F8BC2",
    x"369F77D2",
    x"369F63E4",
    x"369F4FF9",
    x"369F3C10",
    x"369F282A",
    x"369F1446",
    x"369F0065",
    x"369EEC86",
    x"369ED8AA",
    x"369EC4D0",
    x"369EB0F9",
    x"369E9D24",
    x"369E8951",
    x"369E7581",
    x"369E61B4",
    x"369E4DE9",
    x"369E3A20",
    x"369E265A",
    x"369E1297",
    x"369DFED6",
    x"369DEB17",
    x"369DD75B",
    x"369DC3A1",
    x"369DAFEA",
    x"369D9C35",
    x"369D8883",
    x"369D74D3",
    x"369D6126",
    x"369D4D7B",
    x"369D39D2",
    x"369D262C",
    x"369D1289",
    x"369CFEE8",
    x"369CEB49",
    x"369CD7AD",
    x"369CC413",
    x"369CB07C",
    x"369C9CE7",
    x"369C8955",
    x"369C75C5",
    x"369C6237",
    x"369C4EAC",
    x"369C3B24",
    x"369C279D",
    x"369C141A",
    x"369C0098",
    x"369BED1A",
    x"369BD99D",
    x"369BC623",
    x"369BB2AC",
    x"369B9F37",
    x"369B8BC4",
    x"369B7854",
    x"369B64E6",
    x"369B517A",
    x"369B3E11",
    x"369B2AAB",
    x"369B1747",
    x"369B03E5",
    x"369AF086",
    x"369ADD29",
    x"369AC9CE",
    x"369AB676",
    x"369AA321",
    x"369A8FCE",
    x"369A7C7D",
    x"369A692F",
    x"369A55E3",
    x"369A4299",
    x"369A2F52",
    x"369A1C0D",
    x"369A08CB",
    x"3699F58B",
    x"3699E24E",
    x"3699CF12",
    x"3699BBDA",
    x"3699A8A4",
    x"36999570",
    x"3699823E",
    x"36996F0F",
    x"36995BE2",
    x"369948B8",
    x"36993590",
    x"3699226B",
    x"36990F48",
    x"3698FC27",
    x"3698E909",
    x"3698D5ED",
    x"3698C2D3",
    x"3698AFBC",
    x"36989CA7",
    x"36988995",
    x"36987685",
    x"36986377",
    x"3698506C",
    x"36983D63",
    x"36982A5D",
    x"36981758",
    x"36980457",
    x"3697F157",
    x"3697DE5A",
    x"3697CB60",
    x"3697B868",
    x"3697A572",
    x"3697927E",
    x"36977F8D",
    x"36976C9E",
    x"369759B2",
    x"369746C8",
    x"369733E0",
    x"369720FB",
    x"36970E18",
    x"3696FB37",
    x"3696E859",
    x"3696D57D",
    x"3696C2A4",
    x"3696AFCD",
    x"36969CF8",
    x"36968A25",
    x"36967755",
    x"36966488",
    x"369651BC",
    x"36963EF3",
    x"36962C2C",
    x"36961968",
    x"369606A6",
    x"3695F3E6",
    x"3695E129",
    x"3695CE6E",
    x"3695BBB5",
    x"3695A8FF",
    x"3695964B",
    x"3695839A",
    x"369570EA",
    x"36955E3D",
    x"36954B93",
    x"369538EA",
    x"36952645",
    x"369513A1",
    x"36950100",
    x"3694EE61",
    x"3694DBC4",
    x"3694C92A",
    x"3694B692",
    x"3694A3FC",
    x"36949169",
    x"36947ED8",
    x"36946C49",
    x"369459BD",
    x"36944733",
    x"369434AB",
    x"36942225",
    x"36940FA2",
    x"3693FD22",
    x"3693EAA3",
    x"3693D827",
    x"3693C5AD",
    x"3693B335",
    x"3693A0C0",
    x"36938E4D",
    x"36937BDD",
    x"3693696E",
    x"36935702",
    x"36934499",
    x"36933231",
    x"36931FCC",
    x"36930D69",
    x"3692FB09",
    x"3692E8AA",
    x"3692D64E",
    x"3692C3F5",
    x"3692B19D",
    x"36929F48",
    x"36928CF6",
    x"36927AA5",
    x"36926857",
    x"3692560B",
    x"369243C1",
    x"3692317A",
    x"36921F35",
    x"36920CF2",
    x"3691FAB2",
    x"3691E874",
    x"3691D638",
    x"3691C3FE",
    x"3691B1C7",
    x"36919F92",
    x"36918D5F",
    x"36917B2E",
    x"36916900",
    x"369156D4",
    x"369144AA",
    x"36913283",
    x"3691205E",
    x"36910E3B",
    x"3690FC1A",
    x"3690E9FC",
    x"3690D7E0",
    x"3690C5C6",
    x"3690B3AE",
    x"3690A199",
    x"36908F86",
    x"36907D75",
    x"36906B66",
    x"3690595A",
    x"36904750",
    x"36903548",
    x"36902343",
    x"36901140",
    x"368FFF3E",
    x"368FED40",
    x"368FDB43",
    x"368FC949",
    x"368FB751",
    x"368FA55B",
    x"368F9368",
    x"368F8176",
    x"368F6F87",
    x"368F5D9A",
    x"368F4BB0",
    x"368F39C7",
    x"368F27E1",
    x"368F15FD",
    x"368F041C",
    x"368EF23C",
    x"368EE05F",
    x"368ECE84",
    x"368EBCAC",
    x"368EAAD5",
    x"368E9901",
    x"368E872F",
    x"368E755F",
    x"368E6392",
    x"368E51C6",
    x"368E3FFD",
    x"368E2E36",
    x"368E1C72",
    x"368E0AAF",
    x"368DF8EF",
    x"368DE731",
    x"368DD575",
    x"368DC3BC",
    x"368DB204",
    x"368DA04F",
    x"368D8E9C",
    x"368D7CEB",
    x"368D6B3D",
    x"368D5991",
    x"368D47E6",
    x"368D363F",
    x"368D2499",
    x"368D12F5",
    x"368D0154",
    x"368CEFB5",
    x"368CDE18",
    x"368CCC7E",
    x"368CBAE5",
    x"368CA94F",
    x"368C97BB",
    x"368C8629",
    x"368C7499",
    x"368C630C",
    x"368C5180",
    x"368C3FF7",
    x"368C2E70",
    x"368C1CEC",
    x"368C0B69",
    x"368BF9E9",
    x"368BE86B",
    x"368BD6EF",
    x"368BC575",
    x"368BB3FD",
    x"368BA288",
    x"368B9115",
    x"368B7FA4",
    x"368B6E35",
    x"368B5CC8",
    x"368B4B5E",
    x"368B39F5",
    x"368B288F",
    x"368B172B",
    x"368B05C9",
    x"368AF46A",
    x"368AE30C",
    x"368AD1B1",
    x"368AC058",
    x"368AAF01",
    x"368A9DAC",
    x"368A8C5A",
    x"368A7B09",
    x"368A69BB",
    x"368A586F",
    x"368A4725",
    x"368A35DD",
    x"368A2497",
    x"368A1354",
    x"368A0212",
    x"3689F0D3",
    x"3689DF96",
    x"3689CE5B",
    x"3689BD23",
    x"3689ABEC",
    x"36899AB8",
    x"36898985",
    x"36897855",
    x"36896727",
    x"368955FB",
    x"368944D2",
    x"368933AA",
    x"36892285",
    x"36891162",
    x"36890040",
    x"3688EF22",
    x"3688DE05",
    x"3688CCEA",
    x"3688BBD1",
    x"3688AABB",
    x"368899A7",
    x"36888895",
    x"36887785",
    x"36886677",
    x"3688556B",
    x"36884461",
    x"3688335A",
    x"36882255",
    x"36881151",
    x"36880050",
    x"3687EF51",
    x"3687DE54",
    x"3687CD5A",
    x"3687BC61",
    x"3687AB6B",
    x"36879A76",
    x"36878984",
    x"36877894",
    x"368767A6",
    x"368756BA",
    x"368745D0",
    x"368734E8",
    x"36872403",
    x"3687131F",
    x"3687023E",
    x"3686F15F",
    x"3686E082",
    x"3686CFA7",
    x"3686BECE",
    x"3686ADF7",
    x"36869D22",
    x"36868C50",
    x"36867B7F",
    x"36866AB1",
    x"368659E5",
    x"3686491A",
    x"36863852",
    x"3686278C",
    x"368616C8",
    x"36860607",
    x"3685F547",
    x"3685E489",
    x"3685D3CE",
    x"3685C314",
    x"3685B25D",
    x"3685A1A8",
    x"368590F5",
    x"36858044",
    x"36856F95",
    x"36855EE8",
    x"36854E3D",
    x"36853D94",
    x"36852CED",
    x"36851C49",
    x"36850BA6",
    x"3684FB06",
    x"3684EA68",
    x"3684D9CB",
    x"3684C931",
    x"3684B899",
    x"3684A803",
    x"3684976F",
    x"368486DD",
    x"3684764D",
    x"368465C0",
    x"36845534",
    x"368444AA",
    x"36843423",
    x"3684239D",
    x"3684131A",
    x"36840298",
    x"3683F219",
    x"3683E19C",
    x"3683D121",
    x"3683C0A8",
    x"3683B031",
    x"36839FBC",
    x"36838F49",
    x"36837ED8",
    x"36836E69",
    x"36835DFC",
    x"36834D91",
    x"36833D29",
    x"36832CC2",
    x"36831C5E",
    x"36830BFB",
    x"3682FB9B",
    x"3682EB3C",
    x"3682DAE0",
    x"3682CA85",
    x"3682BA2D",
    x"3682A9D7",
    x"36829983",
    x"36828931",
    x"368278E0",
    x"36826892",
    x"36825846",
    x"368247FC",
    x"368237B4",
    x"3682276E",
    x"3682172A",
    x"368206E9",
    x"3681F6A9",
    x"3681E66B",
    x"3681D62F",
    x"3681C5F5",
    x"3681B5BE",
    x"3681A588",
    x"36819554",
    x"36818523",
    x"368174F3",
    x"368164C5",
    x"3681549A",
    x"36814470",
    x"36813449",
    x"36812423",
    x"36811400",
    x"368103DE",
    x"3680F3BF",
    x"3680E3A1",
    x"3680D386",
    x"3680C36C",
    x"3680B355",
    x"3680A33F",
    x"3680932C",
    x"3680831B",
    x"3680730B",
    x"368062FE",
    x"368052F3",
    x"368042E9",
    x"368032E2",
    x"368022DC",
    x"368012D9",
    x"368002D8",
    x"367FE5B1",
    x"367FC5B6",
    x"367FA5BF",
    x"367F85CD",
    x"367F65DE",
    x"367F45F3",
    x"367F260C",
    x"367F062A",
    x"367EE64B",
    x"367EC670",
    x"367EA699",
    x"367E86C6",
    x"367E66F8",
    x"367E472D",
    x"367E2766",
    x"367E07A3",
    x"367DE7E4",
    x"367DC829",
    x"367DA872",
    x"367D88BF",
    x"367D6910",
    x"367D4964",
    x"367D29BD",
    x"367D0A1A",
    x"367CEA7B",
    x"367CCADF",
    x"367CAB48",
    x"367C8BB5",
    x"367C6C25",
    x"367C4C9A",
    x"367C2D12",
    x"367C0D8E",
    x"367BEE0F",
    x"367BCE93",
    x"367BAF1B",
    x"367B8FA7",
    x"367B7037",
    x"367B50CB",
    x"367B3163",
    x"367B11FF",
    x"367AF29E",
    x"367AD342",
    x"367AB3EA",
    x"367A9495",
    x"367A7544",
    x"367A55F8",
    x"367A36AF",
    x"367A176A",
    x"3679F829",
    x"3679D8EC",
    x"3679B9B3",
    x"36799A7E",
    x"36797B4C",
    x"36795C1F",
    x"36793CF5",
    x"36791DCF",
    x"3678FEAE",
    x"3678DF90",
    x"3678C076",
    x"3678A160",
    x"3678824D",
    x"3678633F",
    x"36784435",
    x"3678252E",
    x"3678062B",
    x"3677E72C",
    x"3677C832",
    x"3677A93A",
    x"36778A47",
    x"36776B58",
    x"36774C6C",
    x"36772D85",
    x"36770EA1",
    x"3676EFC1",
    x"3676D0E5",
    x"3676B20D",
    x"36769339",
    x"36767468",
    x"3676559B",
    x"367636D3",
    x"3676180E",
    x"3675F94D",
    x"3675DA8F",
    x"3675BBD6",
    x"36759D20",
    x"36757E6F",
    x"36755FC1",
    x"36754117",
    x"36752271",
    x"367503CE",
    x"3674E530",
    x"3674C695",
    x"3674A7FE",
    x"3674896B",
    x"36746ADC",
    x"36744C50",
    x"36742DC9",
    x"36740F45",
    x"3673F0C5",
    x"3673D249",
    x"3673B3D0",
    x"3673955C",
    x"367376EB",
    x"3673587E",
    x"36733A15",
    x"36731BAF",
    x"3672FD4E",
    x"3672DEF0",
    x"3672C096",
    x"3672A240",
    x"367283ED",
    x"3672659F",
    x"36724754",
    x"3672290D",
    x"36720ACA",
    x"3671EC8A",
    x"3671CE4F",
    x"3671B017",
    x"367191E3",
    x"367173B2",
    x"36715586",
    x"3671375D",
    x"36711938",
    x"3670FB17",
    x"3670DCF9",
    x"3670BEDF",
    x"3670A0C9",
    x"367082B7",
    x"367064A9",
    x"3670469E",
    x"36702897",
    x"36700A94",
    x"366FEC94",
    x"366FCE99",
    x"366FB0A1",
    x"366F92AD",
    x"366F74BC",
    x"366F56CF",
    x"366F38E6",
    x"366F1B01",
    x"366EFD20",
    x"366EDF42",
    x"366EC168",
    x"366EA392",
    x"366E85BF",
    x"366E67F0",
    x"366E4A25",
    x"366E2C5E",
    x"366E0E9A",
    x"366DF0DA",
    x"366DD31E",
    x"366DB565",
    x"366D97B0",
    x"366D79FF",
    x"366D5C52",
    x"366D3EA8",
    x"366D2102",
    x"366D0360",
    x"366CE5C1",
    x"366CC826",
    x"366CAA8F",
    x"366C8CFC",
    x"366C6F6C",
    x"366C51E0",
    x"366C3458",
    x"366C16D3",
    x"366BF952",
    x"366BDBD4",
    x"366BBE5B",
    x"366BA0E5",
    x"366B8373",
    x"366B6604",
    x"366B4899",
    x"366B2B32",
    x"366B0DCE",
    x"366AF06E",
    x"366AD312",
    x"366AB5BA",
    x"366A9865",
    x"366A7B14",
    x"366A5DC6",
    x"366A407C",
    x"366A2336",
    x"366A05F3",
    x"3669E8B4",
    x"3669CB79",
    x"3669AE42",
    x"3669910E",
    x"366973DD",
    x"366956B1",
    x"36693988",
    x"36691C62",
    x"3668FF41",
    x"3668E222",
    x"3668C508",
    x"3668A7F1",
    x"36688ADE",
    x"36686DCE",
    x"366850C3",
    x"366833BA",
    x"366816B6",
    x"3667F9B5",
    x"3667DCB7",
    x"3667BFBD",
    x"3667A2C7",
    x"366785D5",
    x"366768E6",
    x"36674BFA",
    x"36672F13",
    x"3667122F",
    x"3666F54E",
    x"3666D871",
    x"3666BB98",
    x"36669EC2",
    x"366681F0",
    x"36666522",
    x"36664857",
    x"36662B90",
    x"36660ECC",
    x"3665F20C",
    x"3665D550",
    x"3665B897",
    x"36659BE2",
    x"36657F30",
    x"36656282",
    x"366545D7",
    x"36652930",
    x"36650C8D",
    x"3664EFED",
    x"3664D351",
    x"3664B6B8",
    x"36649A23",
    x"36647D92",
    x"36646104",
    x"3664447A",
    x"366427F3",
    x"36640B70",
    x"3663EEF0",
    x"3663D274",
    x"3663B5FB",
    x"36639986",
    x"36637D15",
    x"366360A7",
    x"3663443D",
    x"366327D6",
    x"36630B73",
    x"3662EF13",
    x"3662D2B7",
    x"3662B65F",
    x"36629A09",
    x"36627DB8",
    x"3662616A",
    x"36624520",
    x"366228D9",
    x"36620C95",
    x"3661F056",
    x"3661D419",
    x"3661B7E1",
    x"36619BAB",
    x"36617F7A",
    x"3661634C",
    x"36614721",
    x"36612AFA",
    x"36610ED6",
    x"3660F2B6",
    x"3660D699",
    x"3660BA80",
    x"36609E6B",
    x"36608259",
    x"3660664A",
    x"36604A3F",
    x"36602E38",
    x"36601234",
    x"365FF633",
    x"365FDA36",
    x"365FBE3D",
    x"365FA247",
    x"365F8654",
    x"365F6A65",
    x"365F4E79",
    x"365F3291",
    x"365F16AD",
    x"365EFACC",
    x"365EDEEE",
    x"365EC314",
    x"365EA73D",
    x"365E8B6A",
    x"365E6F9A",
    x"365E53CE",
    x"365E3805",
    x"365E1C40",
    x"365E007E",
    x"365DE4C0",
    x"365DC905",
    x"365DAD4E",
    x"365D919A",
    x"365D75E9",
    x"365D5A3C",
    x"365D3E93",
    x"365D22ED",
    x"365D074A",
    x"365CEBAB",
    x"365CD00F",
    x"365CB477",
    x"365C98E2",
    x"365C7D51",
    x"365C61C3",
    x"365C4638",
    x"365C2AB1",
    x"365C0F2E",
    x"365BF3AD",
    x"365BD831",
    x"365BBCB7",
    x"365BA141",
    x"365B85CF",
    x"365B6A60",
    x"365B4EF4",
    x"365B338C",
    x"365B1828",
    x"365AFCC6",
    x"365AE168",
    x"365AC60E",
    x"365AAAB7",
    x"365A8F63",
    x"365A7413",
    x"365A58C6",
    x"365A3D7D",
    x"365A2237",
    x"365A06F4",
    x"3659EBB5",
    x"3659D079",
    x"3659B541",
    x"36599A0C",
    x"36597EDA",
    x"365963AC",
    x"36594882",
    x"36592D5A",
    x"36591236",
    x"3658F716",
    x"3658DBF8",
    x"3658C0DF",
    x"3658A5C8",
    x"36588AB5",
    x"36586FA6",
    x"36585499",
    x"36583990",
    x"36581E8B",
    x"36580389",
    x"3657E88A",
    x"3657CD8F",
    x"3657B297",
    x"365797A2",
    x"36577CB1",
    x"365761C3",
    x"365746D8",
    x"36572BF1",
    x"3657110D",
    x"3656F62D",
    x"3656DB50",
    x"3656C076",
    x"3656A5A0",
    x"36568ACD",
    x"36566FFD",
    x"36565531",
    x"36563A68",
    x"36561FA2",
    x"365604E0",
    x"3655EA21",
    x"3655CF65",
    x"3655B4AD",
    x"365599F8",
    x"36557F46",
    x"36556498",
    x"365549ED",
    x"36552F46",
    x"365514A1",
    x"3654FA01",
    x"3654DF63",
    x"3654C4C9",
    x"3654AA32",
    x"36548F9E",
    x"3654750E",
    x"36545A81",
    x"36543FF7",
    x"36542571",
    x"36540AEE",
    x"3653F06E",
    x"3653D5F2",
    x"3653BB79",
    x"3653A103",
    x"36538690",
    x"36536C21",
    x"365351B5",
    x"3653374D",
    x"36531CE8",
    x"36530286",
    x"3652E827",
    x"3652CDCC",
    x"3652B373",
    x"3652991F",
    x"36527ECD",
    x"3652647F",
    x"36524A34",
    x"36522FEC",
    x"365215A8",
    x"3651FB67",
    x"3651E129",
    x"3651C6EF",
    x"3651ACB8",
    x"36519284",
    x"36517853",
    x"36515E25",
    x"365143FB",
    x"365129D4",
    x"36510FB1",
    x"3650F591",
    x"3650DB73",
    x"3650C15A",
    x"3650A743",
    x"36508D30",
    x"36507320",
    x"36505913",
    x"36503F0A",
    x"36502503",
    x"36500B00",
    x"364FF101",
    x"364FD704",
    x"364FBD0B",
    x"364FA315",
    x"364F8922",
    x"364F6F33",
    x"364F5546",
    x"364F3B5D",
    x"364F2177",
    x"364F0795",
    x"364EEDB6",
    x"364ED3D9",
    x"364EBA01",
    x"364EA02B",
    x"364E8659",
    x"364E6C89",
    x"364E52BD",
    x"364E38F5",
    x"364E1F2F",
    x"364E056D",
    x"364DEBAE",
    x"364DD1F2",
    x"364DB839",
    x"364D9E84",
    x"364D84D2",
    x"364D6B23",
    x"364D5177",
    x"364D37CE",
    x"364D1E29",
    x"364D0487",
    x"364CEAE8",
    x"364CD14C",
    x"364CB7B3",
    x"364C9E1E",
    x"364C848C",
    x"364C6AFD",
    x"364C5171",
    x"364C37E9",
    x"364C1E63",
    x"364C04E1",
    x"364BEB62",
    x"364BD1E6",
    x"364BB86E",
    x"364B9EF8",
    x"364B8586",
    x"364B6C17",
    x"364B52AB",
    x"364B3942",
    x"364B1FDC",
    x"364B067A",
    x"364AED1B",
    x"364AD3BF",
    x"364ABA66",
    x"364AA110",
    x"364A87BE",
    x"364A6E6E",
    x"364A5522",
    x"364A3BD9",
    x"364A2293",
    x"364A0950",
    x"3649F011",
    x"3649D6D4",
    x"3649BD9B",
    x"3649A465",
    x"36498B32",
    x"36497202",
    x"364958D5",
    x"36493FAC",
    x"36492685",
    x"36490D62",
    x"3648F442",
    x"3648DB25",
    x"3648C20B",
    x"3648A8F5",
    x"36488FE1",
    x"364876D1",
    x"36485DC3",
    x"364844B9",
    x"36482BB2",
    x"364812AE",
    x"3647F9AE",
    x"3647E0B0",
    x"3647C7B5",
    x"3647AEBE",
    x"364795CA",
    x"36477CD9",
    x"364763EA",
    x"36474B00",
    x"36473218",
    x"36471933",
    x"36470051",
    x"3646E773",
    x"3646CE98",
    x"3646B5BF",
    x"36469CEA",
    x"36468418",
    x"36466B49",
    x"3646527D",
    x"364639B4",
    x"364620EF",
    x"3646082C",
    x"3645EF6D",
    x"3645D6B0",
    x"3645BDF7",
    x"3645A541",
    x"36458C8E",
    x"364573DE",
    x"36455B31",
    x"36454287",
    x"364529E0",
    x"3645113D",
    x"3644F89C",
    x"3644DFFE",
    x"3644C764",
    x"3644AECD",
    x"36449638",
    x"36447DA7",
    x"36446519",
    x"36444C8E",
    x"36443406",
    x"36441B81",
    x"364402FF",
    x"3643EA80",
    x"3643D204",
    x"3643B98B",
    x"3643A116",
    x"364388A3",
    x"36437034",
    x"364357C7",
    x"36433F5E",
    x"364326F7",
    x"36430E94",
    x"3642F634",
    x"3642DDD6",
    x"3642C57C",
    x"3642AD25",
    x"364294D1",
    x"36427C80",
    x"36426432",
    x"36424BE7",
    x"3642339F",
    x"36421B5A",
    x"36420318",
    x"3641EAD9",
    x"3641D29D",
    x"3641BA64",
    x"3641A22F",
    x"364189FC",
    x"364171CC",
    x"3641599F",
    x"36414176",
    x"3641294F",
    x"3641112B",
    x"3640F90B",
    x"3640E0ED",
    x"3640C8D3",
    x"3640B0BB",
    x"364098A6",
    x"36408095",
    x"36406886",
    x"3640507B",
    x"36403872",
    x"3640206D",
    x"3640086A",
    x"363FF06A",
    x"363FD86E",
    x"363FC074",
    x"363FA87E",
    x"363F908A",
    x"363F789A",
    x"363F60AC",
    x"363F48C1",
    x"363F30DA",
    x"363F18F5",
    x"363F0114",
    x"363EE935",
    x"363ED159",
    x"363EB981",
    x"363EA1AB",
    x"363E89D8",
    x"363E7208",
    x"363E5A3C",
    x"363E4272",
    x"363E2AAB",
    x"363E12E7",
    x"363DFB26",
    x"363DE368",
    x"363DCBAD",
    x"363DB3F6",
    x"363D9C41",
    x"363D848E",
    x"363D6CDF",
    x"363D5533",
    x"363D3D8A",
    x"363D25E4",
    x"363D0E41",
    x"363CF6A0",
    x"363CDF03",
    x"363CC769",
    x"363CAFD1",
    x"363C983D",
    x"363C80AB",
    x"363C691C",
    x"363C5191",
    x"363C3A08",
    x"363C2282",
    x"363C0AFF",
    x"363BF37F",
    x"363BDC03",
    x"363BC488",
    x"363BAD11",
    x"363B959D",
    x"363B7E2C",
    x"363B66BE",
    x"363B4F52",
    x"363B37EA",
    x"363B2084",
    x"363B0922",
    x"363AF1C2",
    x"363ADA65",
    x"363AC30B",
    x"363AABB5",
    x"363A9461",
    x"363A7D0F",
    x"363A65C1",
    x"363A4E76",
    x"363A372E",
    x"363A1FE8",
    x"363A08A6",
    x"3639F166",
    x"3639DA29",
    x"3639C2EF",
    x"3639ABB9",
    x"36399485",
    x"36397D53",
    x"36396625",
    x"36394EFA",
    x"363937D1",
    x"363920AC",
    x"36390989",
    x"3638F26A",
    x"3638DB4D",
    x"3638C433",
    x"3638AD1C",
    x"36389607",
    x"36387EF6",
    x"363867E8",
    x"363850DC",
    x"363839D3",
    x"363822CE",
    x"36380BCB",
    x"3637F4CB",
    x"3637DDCE",
    x"3637C6D3",
    x"3637AFDC",
    x"363798E7",
    x"363781F6",
    x"36376B07",
    x"3637541B",
    x"36373D32",
    x"3637264C",
    x"36370F68",
    x"3636F888",
    x"3636E1AA",
    x"3636CACF",
    x"3636B3F7",
    x"36369D22",
    x"36368650",
    x"36366F81",
    x"363658B4",
    x"363641EB",
    x"36362B24",
    x"36361460",
    x"3635FD9F",
    x"3635E6E0",
    x"3635D025",
    x"3635B96C",
    x"3635A2B7",
    x"36358C04",
    x"36357554",
    x"36355EA6",
    x"363547FC",
    x"36353154",
    x"36351AB0",
    x"3635040E",
    x"3634ED6F",
    x"3634D6D2",
    x"3634C039",
    x"3634A9A2",
    x"3634930E",
    x"36347C7E",
    x"363465EF",
    x"36344F64",
    x"363438DC",
    x"36342256",
    x"36340BD3",
    x"3633F553",
    x"3633DED6",
    x"3633C85B",
    x"3633B1E4",
    x"36339B6F",
    x"363384FD",
    x"36336E8D",
    x"36335821",
    x"363341B7",
    x"36332B51",
    x"363314ED",
    x"3632FE8B",
    x"3632E82D",
    x"3632D1D1",
    x"3632BB78",
    x"3632A522",
    x"36328ECF",
    x"3632787F",
    x"36326231",
    x"36324BE6",
    x"3632359E",
    x"36321F59",
    x"36320916",
    x"3631F2D7",
    x"3631DC9A",
    x"3631C65F",
    x"3631B028",
    x"363199F3",
    x"363183C1",
    x"36316D92",
    x"36315766",
    x"3631413D",
    x"36312B16",
    x"363114F2",
    x"3630FED1",
    x"3630E8B2",
    x"3630D296",
    x"3630BC7D",
    x"3630A667",
    x"36309054",
    x"36307A43",
    x"36306435",
    x"36304E2A",
    x"36303822",
    x"3630221C",
    x"36300C19",
    x"362FF619",
    x"362FE01C",
    x"362FCA21",
    x"362FB429",
    x"362F9E34",
    x"362F8842",
    x"362F7252",
    x"362F5C65",
    x"362F467B",
    x"362F3093",
    x"362F1AAF",
    x"362F04CD",
    x"362EEEED",
    x"362ED911",
    x"362EC337",
    x"362EAD60",
    x"362E978C",
    x"362E81BA",
    x"362E6BEB",
    x"362E561F",
    x"362E4056",
    x"362E2A8F",
    x"362E14CB",
    x"362DFF0A",
    x"362DE94B",
    x"362DD390",
    x"362DBDD7",
    x"362DA820",
    x"362D926D",
    x"362D7CBC",
    x"362D670D",
    x"362D5162",
    x"362D3BB9",
    x"362D2613",
    x"362D1070",
    x"362CFACF",
    x"362CE531",
    x"362CCF96",
    x"362CB9FD",
    x"362CA467",
    x"362C8ED4",
    x"362C7943",
    x"362C63B5",
    x"362C4E2A",
    x"362C38A2",
    x"362C231C",
    x"362C0D99",
    x"362BF819",
    x"362BE29B",
    x"362BCD20",
    x"362BB7A8",
    x"362BA232",
    x"362B8CBF",
    x"362B774F",
    x"362B61E1",
    x"362B4C77",
    x"362B370E",
    x"362B21A9",
    x"362B0C46",
    x"362AF6E6",
    x"362AE188",
    x"362ACC2D",
    x"362AB6D5",
    x"362AA180",
    x"362A8C2D",
    x"362A76DD",
    x"362A618F",
    x"362A4C44",
    x"362A36FC",
    x"362A21B6",
    x"362A0C74",
    x"3629F733",
    x"3629E1F6",
    x"3629CCBB",
    x"3629B783",
    x"3629A24D",
    x"36298D1A",
    x"362977EA",
    x"362962BC",
    x"36294D91",
    x"36293869",
    x"36292343",
    x"36290E20",
    x"3628F8FF",
    x"3628E3E2",
    x"3628CEC6",
    x"3628B9AE",
    x"3628A498",
    x"36288F85",
    x"36287A74",
    x"36286566",
    x"3628505B",
    x"36283B52",
    x"3628264C",
    x"36281148",
    x"3627FC48",
    x"3627E749",
    x"3627D24E",
    x"3627BD55",
    x"3627A85E",
    x"3627936B",
    x"36277E7A",
    x"3627698B",
    x"3627549F",
    x"36273FB6",
    x"36272ACF",
    x"362715EB",
    x"3627010A",
    x"3626EC2B",
    x"3626D74F",
    x"3626C275",
    x"3626AD9E",
    x"362698CA",
    x"362683F8",
    x"36266F29",
    x"36265A5C",
    x"36264592",
    x"362630CB",
    x"36261C06",
    x"36260744",
    x"3625F284",
    x"3625DDC7",
    x"3625C90D",
    x"3625B455",
    x"36259FA0",
    x"36258AED",
    x"3625763D",
    x"3625618F",
    x"36254CE5",
    x"3625383C",
    x"36252396",
    x"36250EF3",
    x"3624FA53",
    x"3624E5B5",
    x"3624D119",
    x"3624BC80",
    x"3624A7EA",
    x"36249356",
    x"36247EC5",
    x"36246A37",
    x"362455AB",
    x"36244121",
    x"36242C9A",
    x"36241816",
    x"36240394",
    x"3623EF15",
    x"3623DA99",
    x"3623C61F",
    x"3623B1A7",
    x"36239D32",
    x"362388C0",
    x"36237450",
    x"36235FE3",
    x"36234B78",
    x"36233710",
    x"362322AA",
    x"36230E47",
    x"3622F9E7",
    x"3622E589",
    x"3622D12D",
    x"3622BCD4",
    x"3622A87E",
    x"3622942A",
    x"36227FD9",
    x"36226B8A",
    x"3622573E",
    x"362242F5",
    x"36222EAD",
    x"36221A69",
    x"36220627",
    x"3621F1E7",
    x"3621DDAA",
    x"3621C970",
    x"3621B538",
    x"3621A103",
    x"36218CD0",
    x"3621789F",
    x"36216472",
    x"36215046",
    x"36213C1E",
    x"362127F7",
    x"362113D4",
    x"3620FFB2",
    x"3620EB94",
    x"3620D777",
    x"3620C35E",
    x"3620AF47",
    x"36209B32",
    x"36208720",
    x"36207310",
    x"36205F03",
    x"36204AF8",
    x"362036F0",
    x"362022EB",
    x"36200EE8",
    x"361FFAE7",
    x"361FE6E9",
    x"361FD2ED",
    x"361FBEF4",
    x"361FAAFE",
    x"361F9709",
    x"361F8318",
    x"361F6F29",
    x"361F5B3C",
    x"361F4752",
    x"361F336A",
    x"361F1F85",
    x"361F0BA2",
    x"361EF7C2",
    x"361EE3E4",
    x"361ED009",
    x"361EBC30",
    x"361EA85A",
    x"361E9486",
    x"361E80B5",
    x"361E6CE6",
    x"361E591A",
    x"361E4550",
    x"361E3188",
    x"361E1DC3",
    x"361E0A01",
    x"361DF641",
    x"361DE283",
    x"361DCEC8",
    x"361DBB10",
    x"361DA759",
    x"361D93A6",
    x"361D7FF5",
    x"361D6C46",
    x"361D589A",
    x"361D44F0",
    x"361D3148",
    x"361D1DA3",
    x"361D0A01",
    x"361CF661",
    x"361CE2C3",
    x"361CCF28",
    x"361CBB8F",
    x"361CA7F9",
    x"361C9465",
    x"361C80D4",
    x"361C6D45",
    x"361C59B9",
    x"361C462F",
    x"361C32A7",
    x"361C1F22",
    x"361C0BA0",
    x"361BF81F",
    x"361BE4A1",
    x"361BD126",
    x"361BBDAD",
    x"361BAA37",
    x"361B96C3",
    x"361B8351",
    x"361B6FE2",
    x"361B5C75",
    x"361B490B",
    x"361B35A3",
    x"361B223D",
    x"361B0EDA",
    x"361AFB7A",
    x"361AE81B",
    x"361AD4C0",
    x"361AC166",
    x"361AAE0F",
    x"361A9ABB",
    x"361A8769",
    x"361A7419",
    x"361A60CB",
    x"361A4D81",
    x"361A3A38",
    x"361A26F2",
    x"361A13AE",
    x"361A006D",
    x"3619ED2E",
    x"3619D9F2",
    x"3619C6B8",
    x"3619B380",
    x"3619A04B",
    x"36198D18",
    x"361979E8",
    x"361966BA",
    x"3619538E",
    x"36194065",
    x"36192D3E",
    x"36191A19",
    x"361906F7",
    x"3618F3D8",
    x"3618E0BA",
    x"3618CD9F",
    x"3618BA87",
    x"3618A771",
    x"3618945D",
    x"3618814C",
    x"36186E3D",
    x"36185B30",
    x"36184826",
    x"3618351E",
    x"36182219",
    x"36180F16",
    x"3617FC15",
    x"3617E917",
    x"3617D61B",
    x"3617C321",
    x"3617B02A",
    x"36179D35",
    x"36178A43",
    x"36177752",
    x"36176465",
    x"36175179",
    x"36173E90",
    x"36172BAA",
    x"361718C5",
    x"361705E4",
    x"3616F304",
    x"3616E027",
    x"3616CD4C",
    x"3616BA73",
    x"3616A79D",
    x"361694CA",
    x"361681F8",
    x"36166F29",
    x"36165C5C",
    x"36164992",
    x"361636CA",
    x"36162404",
    x"36161141",
    x"3615FE80",
    x"3615EBC1",
    x"3615D905",
    x"3615C64B",
    x"3615B393",
    x"3615A0DE",
    x"36158E2B",
    x"36157B7B",
    x"361568CC",
    x"36155620",
    x"36154377",
    x"361530D0",
    x"36151E2B",
    x"36150B88",
    x"3614F8E8",
    x"3614E64A",
    x"3614D3AE",
    x"3614C115",
    x"3614AE7E",
    x"36149BE9",
    x"36148957",
    x"361476C7",
    x"36146439",
    x"361451AE",
    x"36143F25",
    x"36142C9E",
    x"36141A1A",
    x"36140798",
    x"3613F518",
    x"3613E29A",
    x"3613D01F",
    x"3613BDA6",
    x"3613AB30",
    x"361398BB",
    x"36138649",
    x"361373DA",
    x"3613616D",
    x"36134F02",
    x"36133C99",
    x"36132A32",
    x"361317CE",
    x"3613056C",
    x"3612F30D",
    x"3612E0B0",
    x"3612CE55",
    x"3612BBFC",
    x"3612A9A6",
    x"36129752",
    x"36128500",
    x"361272B0",
    x"36126063",
    x"36124E18",
    x"36123BD0",
    x"36122989",
    x"36121745",
    x"36120504",
    x"3611F2C4",
    x"3611E087",
    x"3611CE4C",
    x"3611BC13",
    x"3611A9DD",
    x"361197A9",
    x"36118577",
    x"36117347",
    x"3611611A",
    x"36114EEF",
    x"36113CC6",
    x"36112AA0",
    x"3611187C",
    x"3611065A",
    x"3610F43A",
    x"3610E21D",
    x"3610D002",
    x"3610BDE9",
    x"3610ABD2",
    x"361099BE",
    x"361087AC",
    x"3610759C",
    x"3610638E",
    x"36105183",
    x"36103F7A",
    x"36102D73",
    x"36101B6F",
    x"3610096C",
    x"360FF76C",
    x"360FE56E",
    x"360FD373",
    x"360FC17A",
    x"360FAF83",
    x"360F9D8E",
    x"360F8B9B",
    x"360F79AB",
    x"360F67BD",
    x"360F55D1",
    x"360F43E7",
    x"360F3200",
    x"360F201B",
    x"360F0E38",
    x"360EFC57",
    x"360EEA79",
    x"360ED89D",
    x"360EC6C3",
    x"360EB4EB",
    x"360EA315",
    x"360E9142",
    x"360E7F71",
    x"360E6DA2",
    x"360E5BD6",
    x"360E4A0B",
    x"360E3843",
    x"360E267D",
    x"360E14BA",
    x"360E02F8",
    x"360DF139",
    x"360DDF7C",
    x"360DCDC1",
    x"360DBC08",
    x"360DAA52",
    x"360D989E",
    x"360D86EC",
    x"360D753C",
    x"360D638E",
    x"360D51E3",
    x"360D403A",
    x"360D2E93",
    x"360D1CEE",
    x"360D0B4C",
    x"360CF9AB",
    x"360CE80D",
    x"360CD671",
    x"360CC4D8",
    x"360CB340",
    x"360CA1AB",
    x"360C9018",
    x"360C7E87",
    x"360C6CF8",
    x"360C5B6C",
    x"360C49E1",
    x"360C3859",
    x"360C26D3",
    x"360C1550",
    x"360C03CE",
    x"360BF24F",
    x"360BE0D1",
    x"360BCF56",
    x"360BBDDE",
    x"360BAC67",
    x"360B9AF2",
    x"360B8980",
    x"360B7810",
    x"360B66A2",
    x"360B5536",
    x"360B43CD",
    x"360B3265",
    x"360B2100",
    x"360B0F9D",
    x"360AFE3C",
    x"360AECDE",
    x"360ADB81",
    x"360ACA27",
    x"360AB8CF",
    x"360AA779",
    x"360A9625",
    x"360A84D3",
    x"360A7384",
    x"360A6236",
    x"360A50EB",
    x"360A3FA2",
    x"360A2E5B",
    x"360A1D16",
    x"360A0BD4",
    x"3609FA93",
    x"3609E955",
    x"3609D819",
    x"3609C6DF",
    x"3609B5A7",
    x"3609A472",
    x"3609933E",
    x"3609820D",
    x"360970DE",
    x"36095FB1",
    x"36094E86",
    x"36093D5D",
    x"36092C36",
    x"36091B12",
    x"360909F0",
    x"3608F8CF",
    x"3608E7B1",
    x"3608D696",
    x"3608C57C",
    x"3608B464",
    x"3608A34F",
    x"3608923B",
    x"3608812A",
    x"3608701B",
    x"36085F0E",
    x"36084E03",
    x"36083CFB",
    x"36082BF4",
    x"36081AF0",
    x"360809ED",
    x"3607F8ED",
    x"3607E7EF",
    x"3607D6F3",
    x"3607C5F9",
    x"3607B502",
    x"3607A40C",
    x"36079319",
    x"36078227",
    x"36077138",
    x"3607604B",
    x"36074F60",
    x"36073E77",
    x"36072D90",
    x"36071CAC",
    x"36070BC9",
    x"3606FAE9",
    x"3606EA0B",
    x"3606D92E",
    x"3606C854",
    x"3606B77C",
    x"3606A6A6",
    x"360695D3",
    x"36068501",
    x"36067431",
    x"36066364",
    x"36065299",
    x"360641CF",
    x"36063108",
    x"36062043",
    x"36060F80",
    x"3605FEBF",
    x"3605EE00",
    x"3605DD44",
    x"3605CC89",
    x"3605BBD0",
    x"3605AB1A",
    x"36059A66",
    x"360589B3",
    x"36057903",
    x"36056855",
    x"360557A9",
    x"360546FF",
    x"36053657",
    x"360525B2",
    x"3605150E",
    x"3605046C",
    x"3604F3CD",
    x"3604E32F",
    x"3604D294",
    x"3604C1FB",
    x"3604B164",
    x"3604A0CE",
    x"3604903B",
    x"36047FAA",
    x"36046F1B",
    x"36045E8F",
    x"36044E04",
    x"36043D7B",
    x"36042CF4",
    x"36041C70",
    x"36040BED",
    x"3603FB6D",
    x"3603EAEF",
    x"3603DA72",
    x"3603C9F8",
    x"3603B980",
    x"3603A90A",
    x"36039895",
    x"36038823",
    x"360377B3",
    x"36036745",
    x"360356DA",
    x"36034670",
    x"36033608",
    x"360325A2",
    x"3603153F",
    x"360304DD",
    x"3602F47D",
    x"3602E420",
    x"3602D3C4",
    x"3602C36B",
    x"3602B313",
    x"3602A2BE",
    x"3602926B",
    x"36028219",
    x"360271CA",
    x"3602617D",
    x"36025132",
    x"360240E9",
    x"360230A2",
    x"3602205D",
    x"3602101A",
    x"3601FFD9",
    x"3601EF9A",
    x"3601DF5D",
    x"3601CF22",
    x"3601BEE9",
    x"3601AEB2",
    x"36019E7D",
    x"36018E4A",
    x"36017E1A",
    x"36016DEB",
    x"36015DBE",
    x"36014D93",
    x"36013D6B",
    x"36012D44",
    x"36011D1F",
    x"36010CFD",
    x"3600FCDC",
    x"3600ECBE",
    x"3600DCA1",
    x"3600CC86",
    x"3600BC6E",
    x"3600AC57",
    x"36009C43",
    x"36008C30",
    x"36007C20",
    x"36006C11",
    x"36005C05",
    x"36004BFA",
    x"36003BF2",
    x"36002BEB",
    x"36001BE7",
    x"36000BE4",
    x"35FFF7C8",
    x"35FFD7CB",
    x"35FFB7D2",
    x"35FF97DD",
    x"35FF77EC",
    x"35FF57FF",
    x"35FF3816",
    x"35FF1831",
    x"35FEF850",
    x"35FED873",
    x"35FEB899",
    x"35FE98C4",
    x"35FE78F3",
    x"35FE5926",
    x"35FE395D",
    x"35FE1998",
    x"35FDF9D7",
    x"35FDDA19",
    x"35FDBA60",
    x"35FD9AAB",
    x"35FD7AF9",
    x"35FD5B4C",
    x"35FD3BA3",
    x"35FD1BFD",
    x"35FCFC5C",
    x"35FCDCBE",
    x"35FCBD24",
    x"35FC9D8F",
    x"35FC7DFD",
    x"35FC5E6F",
    x"35FC3EE5",
    x"35FC1F5F",
    x"35FBFFDE",
    x"35FBE060",
    x"35FBC0E5",
    x"35FBA16F",
    x"35FB81FD",
    x"35FB628F",
    x"35FB4324",
    x"35FB23BE",
    x"35FB045B",
    x"35FAE4FD",
    x"35FAC5A2",
    x"35FAA64C",
    x"35FA86F9",
    x"35FA67AA",
    x"35FA485F",
    x"35FA2918",
    x"35FA09D4",
    x"35F9EA95",
    x"35F9CB5A",
    x"35F9AC22",
    x"35F98CEF",
    x"35F96DBF",
    x"35F94E93",
    x"35F92F6B",
    x"35F91048",
    x"35F8F127",
    x"35F8D20B",
    x"35F8B2F3",
    x"35F893DE",
    x"35F874CE",
    x"35F855C1",
    x"35F836B9",
    x"35F817B4",
    x"35F7F8B3",
    x"35F7D9B5",
    x"35F7BABC",
    x"35F79BC7",
    x"35F77CD5",
    x"35F75DE8",
    x"35F73EFE",
    x"35F72018",
    x"35F70136",
    x"35F6E257",
    x"35F6C37D",
    x"35F6A4A7",
    x"35F685D4",
    x"35F66705",
    x"35F6483A",
    x"35F62973",
    x"35F60AB0",
    x"35F5EBF0",
    x"35F5CD35",
    x"35F5AE7D",
    x"35F58FC9",
    x"35F57119",
    x"35F5526D",
    x"35F533C5",
    x"35F51520",
    x"35F4F67F",
    x"35F4D7E2",
    x"35F4B949",
    x"35F49AB4",
    x"35F47C23",
    x"35F45D95",
    x"35F43F0B",
    x"35F42085",
    x"35F40203",
    x"35F3E385",
    x"35F3C50A",
    x"35F3A694",
    x"35F38821",
    x"35F369B1",
    x"35F34B46",
    x"35F32CDF",
    x"35F30E7B",
    x"35F2F01B",
    x"35F2D1BF",
    x"35F2B367",
    x"35F29512",
    x"35F276C1",
    x"35F25874",
    x"35F23A2B",
    x"35F21BE6",
    x"35F1FDA4",
    x"35F1DF66",
    x"35F1C12C",
    x"35F1A2F6",
    x"35F184C4",
    x"35F16695",
    x"35F1486A",
    x"35F12A43",
    x"35F10C1F",
    x"35F0EE00",
    x"35F0CFE4",
    x"35F0B1CC",
    x"35F093B7",
    x"35F075A7",
    x"35F0579A",
    x"35F03991",
    x"35F01B8C",
    x"35EFFD8A",
    x"35EFDF8C",
    x"35EFC192",
    x"35EFA39C",
    x"35EF85A9",
    x"35EF67BA",
    x"35EF49CF",
    x"35EF2BE8",
    x"35EF0E04",
    x"35EEF025",
    x"35EED248",
    x"35EEB470",
    x"35EE969B",
    x"35EE78CA",
    x"35EE5AFD",
    x"35EE3D34",
    x"35EE1F6E",
    x"35EE01AC",
    x"35EDE3ED",
    x"35EDC633",
    x"35EDA87C",
    x"35ED8AC9",
    x"35ED6D19",
    x"35ED4F6D",
    x"35ED31C5",
    x"35ED1421",
    x"35ECF680",
    x"35ECD8E3",
    x"35ECBB4A",
    x"35EC9DB4",
    x"35EC8023",
    x"35EC6294",
    x"35EC450A",
    x"35EC2783",
    x"35EC0A00",
    x"35EBEC81",
    x"35EBCF05",
    x"35EBB18D",
    x"35EB9419",
    x"35EB76A8",
    x"35EB593B",
    x"35EB3BD2",
    x"35EB1E6C",
    x"35EB010A",
    x"35EAE3AC",
    x"35EAC651",
    x"35EAA8FA",
    x"35EA8BA7",
    x"35EA6E57",
    x"35EA510B",
    x"35EA33C3",
    x"35EA167E",
    x"35E9F93D",
    x"35E9DC00",
    x"35E9BEC6",
    x"35E9A190",
    x"35E9845E",
    x"35E9672F",
    x"35E94A04",
    x"35E92CDD",
    x"35E90FB9",
    x"35E8F299",
    x"35E8D57C",
    x"35E8B863",
    x"35E89B4E",
    x"35E87E3D",
    x"35E8612F",
    x"35E84424",
    x"35E8271E",
    x"35E80A1A",
    x"35E7ED1B",
    x"35E7D01F",
    x"35E7B327",
    x"35E79632",
    x"35E77941",
    x"35E75C54",
    x"35E73F6A",
    x"35E72284",
    x"35E705A2",
    x"35E6E8C3",
    x"35E6CBE8",
    x"35E6AF10",
    x"35E6923C",
    x"35E6756B",
    x"35E6589E",
    x"35E63BD5",
    x"35E61F0F",
    x"35E6024D",
    x"35E5E58F",
    x"35E5C8D4",
    x"35E5AC1D",
    x"35E58F69",
    x"35E572B9",
    x"35E5560C",
    x"35E53963",
    x"35E51CBE",
    x"35E5001C",
    x"35E4E37E",
    x"35E4C6E3",
    x"35E4AA4C",
    x"35E48DB9",
    x"35E47129",
    x"35E4549C",
    x"35E43814",
    x"35E41B8E",
    x"35E3FF0D",
    x"35E3E28F",
    x"35E3C614",
    x"35E3A99D",
    x"35E38D2A",
    x"35E370BA",
    x"35E3544D",
    x"35E337E5",
    x"35E31B7F",
    x"35E2FF1E",
    x"35E2E2C0",
    x"35E2C665",
    x"35E2AA0E",
    x"35E28DBB",
    x"35E2716B",
    x"35E2551E",
    x"35E238D5",
    x"35E21C90",
    x"35E2004E",
    x"35E1E410",
    x"35E1C7D5",
    x"35E1AB9E",
    x"35E18F6A",
    x"35E1733A",
    x"35E1570E",
    x"35E13AE4",
    x"35E11EBF",
    x"35E1029D",
    x"35E0E67E",
    x"35E0CA63",
    x"35E0AE4C",
    x"35E09237",
    x"35E07627",
    x"35E05A1A",
    x"35E03E10",
    x"35E0220A",
    x"35E00608",
    x"35DFEA09",
    x"35DFCE0D",
    x"35DFB215",
    x"35DF9621",
    x"35DF7A30",
    x"35DF5E42",
    x"35DF4258",
    x"35DF2672",
    x"35DF0A8F",
    x"35DEEEAF",
    x"35DED2D3",
    x"35DEB6FA",
    x"35DE9B25",
    x"35DE7F54",
    x"35DE6385",
    x"35DE47BB",
    x"35DE2BF4",
    x"35DE1030",
    x"35DDF46F",
    x"35DDD8B3",
    x"35DDBCF9",
    x"35DDA143",
    x"35DD8591",
    x"35DD69E2",
    x"35DD4E37",
    x"35DD328E",
    x"35DD16EA",
    x"35DCFB49",
    x"35DCDFAB",
    x"35DCC411",
    x"35DCA87A",
    x"35DC8CE7",
    x"35DC7157",
    x"35DC55CA",
    x"35DC3A41",
    x"35DC1EBC",
    x"35DC033A",
    x"35DBE7BB",
    x"35DBCC40",
    x"35DBB0C8",
    x"35DB9554",
    x"35DB79E3",
    x"35DB5E75",
    x"35DB430B",
    x"35DB27A4",
    x"35DB0C41",
    x"35DAF0E1",
    x"35DAD585",
    x"35DABA2C",
    x"35DA9ED6",
    x"35DA8384",
    x"35DA6835",
    x"35DA4CEA",
    x"35DA31A2",
    x"35DA165E",
    x"35D9FB1D",
    x"35D9DFDF",
    x"35D9C4A5",
    x"35D9A96E",
    x"35D98E3A",
    x"35D9730A",
    x"35D957DE",
    x"35D93CB4",
    x"35D9218E",
    x"35D9066C",
    x"35D8EB4D",
    x"35D8D031",
    x"35D8B519",
    x"35D89A04",
    x"35D87EF2",
    x"35D863E4",
    x"35D848D9",
    x"35D82DD2",
    x"35D812CE",
    x"35D7F7CD",
    x"35D7DCD0",
    x"35D7C1D6",
    x"35D7A6DF",
    x"35D78BEC",
    x"35D770FC",
    x"35D75610",
    x"35D73B27",
    x"35D72041",
    x"35D7055F",
    x"35D6EA80",
    x"35D6CFA4",
    x"35D6B4CC",
    x"35D699F7",
    x"35D67F25",
    x"35D66457",
    x"35D6498C",
    x"35D62EC5",
    x"35D61401",
    x"35D5F940",
    x"35D5DE82",
    x"35D5C3C8",
    x"35D5A911",
    x"35D58E5E",
    x"35D573AE",
    x"35D55901",
    x"35D53E58",
    x"35D523B1",
    x"35D5090F",
    x"35D4EE6F",
    x"35D4D3D3",
    x"35D4B93A",
    x"35D49EA5",
    x"35D48413",
    x"35D46984",
    x"35D44EF8",
    x"35D43470",
    x"35D419EB",
    x"35D3FF69",
    x"35D3E4EB",
    x"35D3CA70",
    x"35D3AFF9",
    x"35D39584",
    x"35D37B13",
    x"35D360A5",
    x"35D3463B",
    x"35D32BD4",
    x"35D31170",
    x"35D2F710",
    x"35D2DCB2",
    x"35D2C258",
    x"35D2A802",
    x"35D28DAE",
    x"35D2735E",
    x"35D25912",
    x"35D23EC8",
    x"35D22482",
    x"35D20A3F",
    x"35D1EFFF",
    x"35D1D5C3",
    x"35D1BB8A",
    x"35D1A154",
    x"35D18721",
    x"35D16CF2",
    x"35D152C6",
    x"35D1389E",
    x"35D11E78",
    x"35D10456",
    x"35D0EA37",
    x"35D0D01B",
    x"35D0B603",
    x"35D09BEE",
    x"35D081DC",
    x"35D067CD",
    x"35D04DC2",
    x"35D033BA",
    x"35D019B5",
    x"35CFFFB4",
    x"35CFE5B5",
    x"35CFCBBA",
    x"35CFB1C2",
    x"35CF97CE",
    x"35CF7DDC",
    x"35CF63EE",
    x"35CF4A03",
    x"35CF301C",
    x"35CF1637",
    x"35CEFC56",
    x"35CEE278",
    x"35CEC89E",
    x"35CEAEC6",
    x"35CE94F2",
    x"35CE7B21",
    x"35CE6153",
    x"35CE4788",
    x"35CE2DC1",
    x"35CE13FD",
    x"35CDFA3C",
    x"35CDE07E",
    x"35CDC6C4",
    x"35CDAD0D",
    x"35CD9359",
    x"35CD79A8",
    x"35CD5FFA",
    x"35CD4650",
    x"35CD2CA9",
    x"35CD1305",
    x"35CCF964",
    x"35CCDFC6",
    x"35CCC62C",
    x"35CCAC95",
    x"35CC9301",
    x"35CC7970",
    x"35CC5FE3",
    x"35CC4658",
    x"35CC2CD1",
    x"35CC134D",
    x"35CBF9CC",
    x"35CBE04F",
    x"35CBC6D4",
    x"35CBAD5D",
    x"35CB93E9",
    x"35CB7A78",
    x"35CB610A",
    x"35CB47A0",
    x"35CB2E38",
    x"35CB14D4",
    x"35CAFB73",
    x"35CAE215",
    x"35CAC8BA",
    x"35CAAF63",
    x"35CA960F",
    x"35CA7CBD",
    x"35CA636F",
    x"35CA4A25",
    x"35CA30DD",
    x"35CA1798",
    x"35C9FE57",
    x"35C9E519",
    x"35C9CBDE",
    x"35C9B2A6",
    x"35C99971",
    x"35C9803F",
    x"35C96711",
    x"35C94DE6",
    x"35C934BE",
    x"35C91B99",
    x"35C90277",
    x"35C8E958",
    x"35C8D03C",
    x"35C8B724",
    x"35C89E0F",
    x"35C884FC",
    x"35C86BED",
    x"35C852E1",
    x"35C839D9",
    x"35C820D3",
    x"35C807D0",
    x"35C7EED1",
    x"35C7D5D5",
    x"35C7BCDB",
    x"35C7A3E5",
    x"35C78AF2",
    x"35C77203",
    x"35C75916",
    x"35C7402C",
    x"35C72746",
    x"35C70E63",
    x"35C6F582",
    x"35C6DCA5",
    x"35C6C3CB",
    x"35C6AAF4",
    x"35C69220",
    x"35C67950",
    x"35C66082",
    x"35C647B8",
    x"35C62EF0",
    x"35C6162C",
    x"35C5FD6B",
    x"35C5E4AD",
    x"35C5CBF1",
    x"35C5B33A",
    x"35C59A85",
    x"35C581D3",
    x"35C56924",
    x"35C55079",
    x"35C537D0",
    x"35C51F2B",
    x"35C50688",
    x"35C4EDE9",
    x"35C4D54D",
    x"35C4BCB4",
    x"35C4A41E",
    x"35C48B8B",
    x"35C472FB",
    x"35C45A6E",
    x"35C441E4",
    x"35C4295D",
    x"35C410DA",
    x"35C3F859",
    x"35C3DFDC",
    x"35C3C761",
    x"35C3AEEA",
    x"35C39676",
    x"35C37E04",
    x"35C36596",
    x"35C34D2B",
    x"35C334C3",
    x"35C31C5E",
    x"35C303FC",
    x"35C2EB9D",
    x"35C2D341",
    x"35C2BAE8",
    x"35C2A292",
    x"35C28A3F",
    x"35C271EF",
    x"35C259A3",
    x"35C24159",
    x"35C22912",
    x"35C210CF",
    x"35C1F88E",
    x"35C1E051",
    x"35C1C816",
    x"35C1AFDF",
    x"35C197AA",
    x"35C17F79",
    x"35C1674A",
    x"35C14F1F",
    x"35C136F7",
    x"35C11ED1",
    x"35C106AF",
    x"35C0EE8F",
    x"35C0D673",
    x"35C0BE5A",
    x"35C0A644",
    x"35C08E30",
    x"35C07620",
    x"35C05E13",
    x"35C04609",
    x"35C02E01",
    x"35C015FD",
    x"35BFFDFC",
    x"35BFE5FE",
    x"35BFCE02",
    x"35BFB60A",
    x"35BF9E15",
    x"35BF8622",
    x"35BF6E33",
    x"35BF5647",
    x"35BF3E5E",
    x"35BF2677",
    x"35BF0E94",
    x"35BEF6B4",
    x"35BEDED6",
    x"35BEC6FC",
    x"35BEAF25",
    x"35BE9750",
    x"35BE7F7F",
    x"35BE67B0",
    x"35BE4FE5",
    x"35BE381C",
    x"35BE2057",
    x"35BE0894",
    x"35BDF0D5",
    x"35BDD918",
    x"35BDC15E",
    x"35BDA9A8",
    x"35BD91F4",
    x"35BD7A43",
    x"35BD6295",
    x"35BD4AEB",
    x"35BD3343",
    x"35BD1B9E",
    x"35BD03FC",
    x"35BCEC5D",
    x"35BCD4C1",
    x"35BCBD28",
    x"35BCA591",
    x"35BC8DFE",
    x"35BC766E",
    x"35BC5EE1",
    x"35BC4756",
    x"35BC2FCF",
    x"35BC184A",
    x"35BC00C9",
    x"35BBE94A",
    x"35BBD1CE",
    x"35BBBA56",
    x"35BBA2E0",
    x"35BB8B6D",
    x"35BB73FD",
    x"35BB5C90",
    x"35BB4526",
    x"35BB2DBF",
    x"35BB165A",
    x"35BAFEF9",
    x"35BAE79B",
    x"35BAD03F",
    x"35BAB8E7",
    x"35BAA191",
    x"35BA8A3E",
    x"35BA72EE",
    x"35BA5BA1",
    x"35BA4457",
    x"35BA2D10",
    x"35BA15CC",
    x"35B9FE8B",
    x"35B9E74D",
    x"35B9D011",
    x"35B9B8D8",
    x"35B9A1A3",
    x"35B98A70",
    x"35B97340",
    x"35B95C13",
    x"35B944E9",
    x"35B92DC2",
    x"35B9169E",
    x"35B8FF7C",
    x"35B8E85E",
    x"35B8D142",
    x"35B8BA2A",
    x"35B8A314",
    x"35B88C01",
    x"35B874F1",
    x"35B85DE4",
    x"35B846D9",
    x"35B82FD2",
    x"35B818CD",
    x"35B801CC",
    x"35B7EACD",
    x"35B7D3D1",
    x"35B7BCD8",
    x"35B7A5E2",
    x"35B78EEE",
    x"35B777FE",
    x"35B76110",
    x"35B74A26",
    x"35B7333E",
    x"35B71C59",
    x"35B70577",
    x"35B6EE98",
    x"35B6D7BB",
    x"35B6C0E2",
    x"35B6AA0B",
    x"35B69337",
    x"35B67C66",
    x"35B66598",
    x"35B64ECD",
    x"35B63804",
    x"35B6213F",
    x"35B60A7C",
    x"35B5F3BC",
    x"35B5DCFF",
    x"35B5C645",
    x"35B5AF8E",
    x"35B598D9",
    x"35B58227",
    x"35B56B78",
    x"35B554CC",
    x"35B53E23",
    x"35B5277D",
    x"35B510D9",
    x"35B4FA39",
    x"35B4E39B",
    x"35B4CD00",
    x"35B4B668",
    x"35B49FD2",
    x"35B48940",
    x"35B472B0",
    x"35B45C23",
    x"35B44599",
    x"35B42F12",
    x"35B4188D",
    x"35B4020B",
    x"35B3EB8D",
    x"35B3D511",
    x"35B3BE97",
    x"35B3A821",
    x"35B391AD",
    x"35B37B3C",
    x"35B364CE",
    x"35B34E63",
    x"35B337FB",
    x"35B32195",
    x"35B30B32",
    x"35B2F4D2",
    x"35B2DE75",
    x"35B2C81B",
    x"35B2B1C3",
    x"35B29B6E",
    x"35B2851C",
    x"35B26ECD",
    x"35B25881",
    x"35B24237",
    x"35B22BF0",
    x"35B215AC",
    x"35B1FF6B",
    x"35B1E92C",
    x"35B1D2F0",
    x"35B1BCB7",
    x"35B1A681",
    x"35B1904E",
    x"35B17A1D",
    x"35B163EF",
    x"35B14DC4",
    x"35B1379C",
    x"35B12176",
    x"35B10B53",
    x"35B0F533",
    x"35B0DF16",
    x"35B0C8FC",
    x"35B0B2E4",
    x"35B09CCF",
    x"35B086BD",
    x"35B070AD",
    x"35B05AA1",
    x"35B04497",
    x"35B02E8F",
    x"35B0188B",
    x"35B00289",
    x"35AFEC8A",
    x"35AFD68E",
    x"35AFC095",
    x"35AFAA9E",
    x"35AF94AA",
    x"35AF7EB9",
    x"35AF68CA",
    x"35AF52DF",
    x"35AF3CF6",
    x"35AF270F",
    x"35AF112C",
    x"35AEFB4B",
    x"35AEE56D",
    x"35AECF92",
    x"35AEB9B9",
    x"35AEA3E3",
    x"35AE8E10",
    x"35AE7840",
    x"35AE6272",
    x"35AE4CA7",
    x"35AE36DF",
    x"35AE2119",
    x"35AE0B57",
    x"35ADF597",
    x"35ADDFD9",
    x"35ADCA1F",
    x"35ADB467",
    x"35AD9EB2",
    x"35AD88FF",
    x"35AD734F",
    x"35AD5DA2",
    x"35AD47F8",
    x"35AD3250",
    x"35AD1CAB",
    x"35AD0709",
    x"35ACF16A",
    x"35ACDBCD",
    x"35ACC633",
    x"35ACB09B",
    x"35AC9B06",
    x"35AC8574",
    x"35AC6FE5",
    x"35AC5A58",
    x"35AC44CE",
    x"35AC2F47",
    x"35AC19C3",
    x"35AC0441",
    x"35ABEEC2",
    x"35ABD945",
    x"35ABC3CB",
    x"35ABAE54",
    x"35AB98E0",
    x"35AB836E",
    x"35AB6DFF",
    x"35AB5892",
    x"35AB4329",
    x"35AB2DC2",
    x"35AB185D",
    x"35AB02FC",
    x"35AAED9D",
    x"35AAD840",
    x"35AAC2E6",
    x"35AAAD8F",
    x"35AA983B",
    x"35AA82E9",
    x"35AA6D9A",
    x"35AA584E",
    x"35AA4304",
    x"35AA2DBD",
    x"35AA1879",
    x"35AA0337",
    x"35A9EDF8",
    x"35A9D8BC",
    x"35A9C382",
    x"35A9AE4B",
    x"35A99916",
    x"35A983E4",
    x"35A96EB5",
    x"35A95989",
    x"35A9445F",
    x"35A92F38",
    x"35A91A13",
    x"35A904F1",
    x"35A8EFD2",
    x"35A8DAB5",
    x"35A8C59B",
    x"35A8B084",
    x"35A89B6F",
    x"35A8865D",
    x"35A8714D",
    x"35A85C41",
    x"35A84736",
    x"35A8322F",
    x"35A81D2A",
    x"35A80828",
    x"35A7F328",
    x"35A7DE2B",
    x"35A7C930",
    x"35A7B438",
    x"35A79F43",
    x"35A78A51",
    x"35A77561",
    x"35A76073",
    x"35A74B89",
    x"35A736A0",
    x"35A721BB",
    x"35A70CD8",
    x"35A6F7F8",
    x"35A6E31A",
    x"35A6CE3F",
    x"35A6B966",
    x"35A6A491",
    x"35A68FBD",
    x"35A67AED",
    x"35A6661F",
    x"35A65153",
    x"35A63C8A",
    x"35A627C4",
    x"35A61300",
    x"35A5FE3F",
    x"35A5E981",
    x"35A5D4C5",
    x"35A5C00B",
    x"35A5AB55",
    x"35A596A1",
    x"35A581EF",
    x"35A56D40",
    x"35A55894",
    x"35A543EA",
    x"35A52F43",
    x"35A51A9E",
    x"35A505FC",
    x"35A4F15D",
    x"35A4DCC0",
    x"35A4C826",
    x"35A4B38E",
    x"35A49EF9",
    x"35A48A66",
    x"35A475D6",
    x"35A46149",
    x"35A44CBE",
    x"35A43835",
    x"35A423B0",
    x"35A40F2C",
    x"35A3FAAC",
    x"35A3E62E",
    x"35A3D1B2",
    x"35A3BD39",
    x"35A3A8C3",
    x"35A3944F",
    x"35A37FDE",
    x"35A36B6F",
    x"35A35703",
    x"35A34299",
    x"35A32E32",
    x"35A319CE",
    x"35A3056C",
    x"35A2F10D",
    x"35A2DCB0",
    x"35A2C855",
    x"35A2B3FE",
    x"35A29FA8",
    x"35A28B56",
    x"35A27706",
    x"35A262B8",
    x"35A24E6D",
    x"35A23A24",
    x"35A225DE",
    x"35A2119B",
    x"35A1FD5A",
    x"35A1E91C",
    x"35A1D4E0",
    x"35A1C0A6",
    x"35A1AC70",
    x"35A1983B",
    x"35A18409",
    x"35A16FDA",
    x"35A15BAE",
    x"35A14783",
    x"35A1335C",
    x"35A11F36",
    x"35A10B14",
    x"35A0F6F4",
    x"35A0E2D6",
    x"35A0CEBB",
    x"35A0BAA2",
    x"35A0A68C",
    x"35A09279",
    x"35A07E68",
    x"35A06A59",
    x"35A0564D",
    x"35A04244",
    x"35A02E3D",
    x"35A01A38",
    x"35A00636",
    x"359FF236",
    x"359FDE39",
    x"359FCA3F",
    x"359FB647",
    x"359FA251",
    x"359F8E5E",
    x"359F7A6E",
    x"359F6680",
    x"359F5294",
    x"359F3EAB",
    x"359F2AC4",
    x"359F16E0",
    x"359F02FF",
    x"359EEF20",
    x"359EDB43",
    x"359EC769",
    x"359EB391",
    x"359E9FBC",
    x"359E8BE9",
    x"359E7819",
    x"359E644B",
    x"359E5080",
    x"359E3CB7",
    x"359E28F1",
    x"359E152D",
    x"359E016B",
    x"359DEDAC",
    x"359DD9F0",
    x"359DC636",
    x"359DB27E",
    x"359D9EC9",
    x"359D8B17",
    x"359D7767",
    x"359D63B9",
    x"359D500E",
    x"359D3C65",
    x"359D28BF",
    x"359D151B",
    x"359D0179",
    x"359CEDDA",
    x"359CDA3E",
    x"359CC6A4",
    x"359CB30C",
    x"359C9F77",
    x"359C8BE4",
    x"359C7854",
    x"359C64C6",
    x"359C513B",
    x"359C3DB2",
    x"359C2A2B",
    x"359C16A7",
    x"359C0326",
    x"359BEFA7",
    x"359BDC2A",
    x"359BC8AF",
    x"359BB538",
    x"359BA1C2",
    x"359B8E4F",
    x"359B7ADF",
    x"359B6770",
    x"359B5405",
    x"359B409B",
    x"359B2D35",
    x"359B19D0",
    x"359B066E",
    x"359AF30F",
    x"359ADFB1",
    x"359ACC57",
    x"359AB8FE",
    x"359AA5A8",
    x"359A9255",
    x"359A7F04",
    x"359A6BB5",
    x"359A5869",
    x"359A451F",
    x"359A31D8",
    x"359A1E93",
    x"359A0B50",
    x"3599F810",
    x"3599E4D2",
    x"3599D197",
    x"3599BE5E",
    x"3599AB27",
    x"359997F3",
    x"359984C1",
    x"35997192",
    x"35995E65",
    x"35994B3A",
    x"35993812",
    x"359924EC",
    x"359911C9",
    x"3598FEA7",
    x"3598EB89",
    x"3598D86D",
    x"3598C553",
    x"3598B23B",
    x"35989F26",
    x"35988C13",
    x"35987903",
    x"359865F5",
    x"359852EA",
    x"35983FE1",
    x"35982CDA",
    x"359819D5",
    x"359806D3",
    x"3597F3D4",
    x"3597E0D6",
    x"3597CDDB",
    x"3597BAE3",
    x"3597A7ED",
    x"359794F9",
    x"35978207",
    x"35976F18",
    x"35975C2C",
    x"35974941",
    x"35973659",
    x"35972374",
    x"35971090",
    x"3596FDB0",
    x"3596EAD1",
    x"3596D7F5",
    x"3596C51B",
    x"3596B244",
    x"35969F6E",
    x"35968C9C",
    x"359679CB",
    x"359666FD",
    x"35965432",
    x"35964168",
    x"35962EA1",
    x"35961BDD",
    x"3596091A",
    x"3595F65A",
    x"3595E39D",
    x"3595D0E1",
    x"3595BE28",
    x"3595AB72",
    x"359598BE",
    x"3595860C",
    x"3595735C",
    x"359560AF",
    x"35954E04",
    x"35953B5B",
    x"359528B5",
    x"35951611",
    x"35950370",
    x"3594F0D0",
    x"3594DE33",
    x"3594CB99",
    x"3594B900",
    x"3594A66A",
    x"359493D7",
    x"35948146",
    x"35946EB7",
    x"35945C2A",
    x"3594499F",
    x"35943717",
    x"35942492",
    x"3594120E",
    x"3593FF8D",
    x"3593ED0E",
    x"3593DA92",
    x"3593C818",
    x"3593B5A0",
    x"3593A32A",
    x"359390B7",
    x"35937E46",
    x"35936BD8",
    x"3593596B",
    x"35934701",
    x"35933499",
    x"35932234",
    x"35930FD1",
    x"3592FD70",
    x"3592EB12",
    x"3592D8B5",
    x"3592C65B",
    x"3592B404",
    x"3592A1AE",
    x"35928F5B",
    x"35927D0B",
    x"35926ABC",
    x"35925870",
    x"35924626",
    x"359233DE",
    x"35922199",
    x"35920F56",
    x"3591FD15",
    x"3591EAD7",
    x"3591D89A",
    x"3591C660",
    x"3591B429",
    x"3591A1F3",
    x"35918FC0",
    x"35917D90",
    x"35916B61",
    x"35915935",
    x"3591470B",
    x"359134E3",
    x"359122BD",
    x"3591109A",
    x"3590FE79",
    x"3590EC5B",
    x"3590DA3E",
    x"3590C824",
    x"3590B60C",
    x"3590A3F7",
    x"359091E3",
    x"35907FD2",
    x"35906DC3",
    x"35905BB7",
    x"359049AC",
    x"359037A4",
    x"3590259E",
    x"3590139B",
    x"35900199",
    x"358FEF9A",
    x"358FDD9E",
    x"358FCBA3",
    x"358FB9AB",
    x"358FA7B5",
    x"358F95C1",
    x"358F83CF",
    x"358F71E0",
    x"358F5FF3",
    x"358F4E08",
    x"358F3C1F",
    x"358F2A39",
    x"358F1855",
    x"358F0673",
    x"358EF493",
    x"358EE2B6",
    x"358ED0DA",
    x"358EBF01",
    x"358EAD2B",
    x"358E9B56",
    x"358E8984",
    x"358E77B4",
    x"358E65E6",
    x"358E541A",
    x"358E4251",
    x"358E308A",
    x"358E1EC5",
    x"358E0D02",
    x"358DFB41",
    x"358DE983",
    x"358DD7C7",
    x"358DC60D",
    x"358DB455",
    x"358DA2A0",
    x"358D90ED",
    x"358D7F3C",
    x"358D6D8D",
    x"358D5BE0",
    x"358D4A36",
    x"358D388E",
    x"358D26E8",
    x"358D1544",
    x"358D03A3",
    x"358CF203",
    x"358CE066",
    x"358CCECB",
    x"358CBD32",
    x"358CAB9C",
    x"358C9A08",
    x"358C8875",
    x"358C76E5",
    x"358C6558",
    x"358C53CC",
    x"358C4243",
    x"358C30BB",
    x"358C1F36",
    x"358C0DB4",
    x"358BFC33",
    x"358BEAB5",
    x"358BD938",
    x"358BC7BE",
    x"358BB646",
    x"358BA4D1",
    x"358B935D",
    x"358B81EC",
    x"358B707D",
    x"358B5F10",
    x"358B4DA5",
    x"358B3C3C",
    x"358B2AD6",
    x"358B1972",
    x"358B0810",
    x"358AF6B0",
    x"358AE552",
    x"358AD3F6",
    x"358AC29D",
    x"358AB146",
    x"358A9FF1",
    x"358A8E9E",
    x"358A7D4D",
    x"358A6BFE",
    x"358A5AB2",
    x"358A4968",
    x"358A3820",
    x"358A26DA",
    x"358A1596",
    x"358A0454",
    x"3589F315",
    x"3589E1D7",
    x"3589D09C",
    x"3589BF63",
    x"3589AE2C",
    x"35899CF8",
    x"35898BC5",
    x"35897A95",
    x"35896967",
    x"3589583A",
    x"35894711",
    x"358935E9",
    x"358924C3",
    x"358913A0",
    x"3589027E",
    x"3588F15F",
    x"3588E042",
    x"3588CF27",
    x"3588BE0E",
    x"3588ACF7",
    x"35889BE3",
    x"35888AD0",
    x"358879C0",
    x"358868B2",
    x"358857A6",
    x"3588469C",
    x"35883594",
    x"3588248F",
    x"3588138B",
    x"3588028A",
    x"3587F18A",
    x"3587E08D",
    x"3587CF92",
    x"3587BE99",
    x"3587ADA3",
    x"35879CAE",
    x"35878BBC",
    x"35877ACB",
    x"358769DD",
    x"358758F1",
    x"35874807",
    x"3587371F",
    x"35872639",
    x"35871555",
    x"35870473",
    x"3586F394",
    x"3586E2B7",
    x"3586D1DB",
    x"3586C102",
    x"3586B02B",
    x"35869F56",
    x"35868E83",
    x"35867DB2",
    x"35866CE4",
    x"35865C17",
    x"35864B4D",
    x"35863A84",
    x"358629BE",
    x"358618FA",
    x"35860838",
    x"3585F778",
    x"3585E6BA",
    x"3585D5FE",
    x"3585C545",
    x"3585B48D",
    x"3585A3D7",
    x"35859324",
    x"35858273",
    x"358571C3",
    x"35856116",
    x"3585506B",
    x"35853FC2",
    x"35852F1B",
    x"35851E76",
    x"35850DD4",
    x"3584FD33",
    x"3584EC94",
    x"3584DBF8",
    x"3584CB5D",
    x"3584BAC5",
    x"3584AA2F",
    x"3584999A",
    x"35848908",
    x"35847878",
    x"358467EA",
    x"3584575E",
    x"358446D4",
    x"3584364C",
    x"358425C7",
    x"35841543",
    x"358404C1",
    x"3583F442",
    x"3583E3C4",
    x"3583D349",
    x"3583C2CF",
    x"3583B258",
    x"3583A1E3",
    x"35839170",
    x"358380FE",
    x"3583708F",
    x"35836022",
    x"35834FB7",
    x"35833F4E",
    x"35832EE7",
    x"35831E83",
    x"35830E20",
    x"3582FDBF",
    x"3582ED60",
    x"3582DD04",
    x"3582CCA9",
    x"3582BC51",
    x"3582ABFA",
    x"35829BA6",
    x"35828B53",
    x"35827B03",
    x"35826AB4",
    x"35825A68",
    x"35824A1E",
    x"358239D6",
    x"3582298F",
    x"3582194B",
    x"35820909",
    x"3581F8C9",
    x"3581E88B",
    x"3581D84F",
    x"3581C815",
    x"3581B7DD",
    x"3581A7A7",
    x"35819773",
    x"35818741",
    x"35817711",
    x"358166E3",
    x"358156B7",
    x"3581468D",
    x"35813666",
    x"35812640",
    x"3581161C",
    x"358105FA",
    x"3580F5DB",
    x"3580E5BD",
    x"3580D5A1",
    x"3580C587",
    x"3580B570",
    x"3580A55A",
    x"35809546",
    x"35808535",
    x"35807525",
    x"35806518",
    x"3580550C",
    x"35804502",
    x"358034FB",
    x"358024F5",
    x"358014F1",
    x"358004F0",
    x"357FE9E0",
    x"357FC9E5",
    x"357FA9EE",
    x"357F89FB",
    x"357F6A0B",
    x"357F4A20",
    x"357F2A39",
    x"357F0A56",
    x"357EEA76",
    x"357ECA9B",
    x"357EAAC4",
    x"357E8AF0",
    x"357E6B21",
    x"357E4B55",
    x"357E2B8E",
    x"357E0BCB",
    x"357DEC0B",
    x"357DCC50",
    x"357DAC98",
    x"357D8CE4",
    x"357D6D35",
    x"357D4D89",
    x"357D2DE1",
    x"357D0E3E",
    x"357CEE9E",
    x"357CCF02",
    x"357CAF6A",
    x"357C8FD6",
    x"357C7046",
    x"357C50BA",
    x"357C3132",
    x"357C11AE",
    x"357BF22D",
    x"357BD2B1",
    x"357BB339",
    x"357B93C4",
    x"357B7454",
    x"357B54E7",
    x"357B357F",
    x"357B161A",
    x"357AF6B9",
    x"357AD75C",
    x"357AB803",
    x"357A98AE",
    x"357A795D",
    x"357A5A10",
    x"357A3AC7",
    x"357A1B81",
    x"3579FC40",
    x"3579DD02",
    x"3579BDC8",
    x"35799E93",
    x"35797F61",
    x"35796033",
    x"35794109",
    x"357921E3",
    x"357902C0",
    x"3578E3A2",
    x"3578C487",
    x"3578A571",
    x"3578865E",
    x"3578674F",
    x"35784844",
    x"3578293D",
    x"35780A3A",
    x"3577EB3B",
    x"3577CC3F",
    x"3577AD47",
    x"35778E54",
    x"35776F64",
    x"35775078",
    x"35773190",
    x"357712AC",
    x"3576F3CB",
    x"3576D4EF",
    x"3576B616",
    x"35769741",
    x"35767870",
    x"357659A3",
    x"35763ADA",
    x"35761C14",
    x"3575FD53",
    x"3575DE95",
    x"3575BFDB",
    x"3575A125",
    x"35758273",
    x"357563C4",
    x"3575451A",
    x"35752673",
    x"357507D0",
    x"3574E931",
    x"3574CA96",
    x"3574ABFE",
    x"35748D6B",
    x"35746EDB",
    x"3574504F",
    x"357431C7",
    x"35741343",
    x"3573F4C2",
    x"3573D646",
    x"3573B7CD",
    x"35739958",
    x"35737AE6",
    x"35735C79",
    x"35733E0F",
    x"35731FA9",
    x"35730147",
    x"3572E2E9",
    x"3572C48F",
    x"3572A638",
    x"357287E5",
    x"35726996",
    x"35724B4B",
    x"35722D03",
    x"35720EBF",
    x"3571F07F",
    x"3571D243",
    x"3571B40B",
    x"357195D6",
    x"357177A5",
    x"35715978",
    x"35713B4F",
    x"35711D29",
    x"3570FF08",
    x"3570E0EA",
    x"3570C2CF",
    x"3570A4B9",
    x"357086A6",
    x"35706897",
    x"35704A8C",
    x"35702C85",
    x"35700E81",
    x"356FF081",
    x"356FD285",
    x"356FB48C",
    x"356F9698",
    x"356F78A7",
    x"356F5ABA",
    x"356F3CD0",
    x"356F1EEA",
    x"356F0108",
    x"356EE32A",
    x"356EC550",
    x"356EA779",
    x"356E89A6",
    x"356E6BD6",
    x"356E4E0B",
    x"356E3043",
    x"356E127F",
    x"356DF4BE",
    x"356DD702",
    x"356DB948",
    x"356D9B93",
    x"356D7DE2",
    x"356D6034",
    x"356D428A",
    x"356D24E3",
    x"356D0740",
    x"356CE9A1",
    x"356CCC06",
    x"356CAE6E",
    x"356C90DA",
    x"356C734A",
    x"356C55BD",
    x"356C3835",
    x"356C1AAF",
    x"356BFD2E",
    x"356BDFB0",
    x"356BC236",
    x"356BA4C0",
    x"356B874D",
    x"356B69DE",
    x"356B4C72",
    x"356B2F0B",
    x"356B11A7",
    x"356AF446",
    x"356AD6EA",
    x"356AB990",
    x"356A9C3B",
    x"356A7EE9",
    x"356A619B",
    x"356A4451",
    x"356A270A",
    x"356A09C7",
    x"3569EC88",
    x"3569CF4C",
    x"3569B214",
    x"356994E0",
    x"356977AF",
    x"35695A82",
    x"35693D58",
    x"35692032",
    x"35690310",
    x"3568E5F2",
    x"3568C8D7",
    x"3568ABBF",
    x"35688EAC",
    x"3568719C",
    x"3568548F",
    x"35683787",
    x"35681A81",
    x"3567FD80",
    x"3567E082",
    x"3567C388",
    x"3567A691",
    x"3567899E",
    x"35676CAF",
    x"35674FC3",
    x"356732DB",
    x"356715F6",
    x"3566F915",
    x"3566DC38",
    x"3566BF5E",
    x"3566A288",
    x"356685B6",
    x"356668E7",
    x"35664C1B",
    x"35662F54",
    x"35661290",
    x"3565F5CF",
    x"3565D912",
    x"3565BC59",
    x"35659FA3",
    x"356582F1",
    x"35656642",
    x"35654997",
    x"35652CF0",
    x"3565104C",
    x"3564F3AC",
    x"3564D70F",
    x"3564BA76",
    x"35649DE1",
    x"3564814F",
    x"356464C0",
    x"35644835",
    x"35642BAE",
    x"35640F2B",
    x"3563F2AA",
    x"3563D62E",
    x"3563B9B5",
    x"35639D3F",
    x"356380CE",
    x"3563645F",
    x"356347F4",
    x"35632B8D",
    x"35630F2A",
    x"3562F2C9",
    x"3562D66D",
    x"3562BA14",
    x"35629DBE",
    x"3562816C",
    x"3562651E",
    x"356248D3",
    x"35622C8C",
    x"35621048",
    x"3561F408",
    x"3561D7CB",
    x"3561BB92",
    x"35619F5C",
    x"3561832A",
    x"356166FB",
    x"35614AD0",
    x"35612EA9",
    x"35611285",
    x"3560F664",
    x"3560DA47",
    x"3560BE2D",
    x"3560A217",
    x"35608605",
    x"356069F6",
    x"35604DEA",
    x"356031E2",
    x"356015DE",
    x"355FF9DD",
    x"355FDDDF",
    x"355FC1E5",
    x"355FA5EF",
    x"355F89FC",
    x"355F6E0C",
    x"355F5220",
    x"355F3638",
    x"355F1A53",
    x"355EFE71",
    x"355EE293",
    x"355EC6B9",
    x"355EAAE2",
    x"355E8F0E",
    x"355E733E",
    x"355E5771",
    x"355E3BA8",
    x"355E1FE2",
    x"355E0420",
    x"355DE861",
    x"355DCCA6",
    x"355DB0EE",
    x"355D953A",
    x"355D7989",
    x"355D5DDB",
    x"355D4231",
    x"355D268B",
    x"355D0AE8",
    x"355CEF48",
    x"355CD3AC",
    x"355CB813",
    x"355C9C7E",
    x"355C80EC",
    x"355C655E",
    x"355C49D3",
    x"355C2E4B",
    x"355C12C7",
    x"355BF746",
    x"355BDBC9",
    x"355BC04F",
    x"355BA4D9",
    x"355B8966",
    x"355B6DF7",
    x"355B528B",
    x"355B3722",
    x"355B1BBD",
    x"355B005B",
    x"355AE4FD",
    x"355AC9A2",
    x"355AAE4A",
    x"355A92F6",
    x"355A77A6",
    x"355A5C59",
    x"355A410F",
    x"355A25C8",
    x"355A0A85",
    x"3559EF46",
    x"3559D409",
    x"3559B8D1",
    x"35599D9B",
    x"35598269",
    x"3559673B",
    x"35594C0F",
    x"355930E8",
    x"355915C3",
    x"3558FAA2",
    x"3558DF85",
    x"3558C46A",
    x"3558A953",
    x"35588E40",
    x"35587330",
    x"35585823",
    x"35583D1A",
    x"35582214",
    x"35580711",
    x"3557EC12",
    x"3557D116",
    x"3557B61E",
    x"35579B29",
    x"35578037",
    x"35576549",
    x"35574A5E",
    x"35572F76",
    x"35571492",
    x"3556F9B1",
    x"3556DED3",
    x"3556C3F9",
    x"3556A922",
    x"35568E4F",
    x"3556737F",
    x"355658B2",
    x"35563DE9",
    x"35562323",
    x"35560860",
    x"3555EDA1",
    x"3555D2E4",
    x"3555B82C",
    x"35559D76",
    x"355582C4",
    x"35556816",
    x"35554D6A",
    x"355532C2",
    x"3555181E",
    x"3554FD7C",
    x"3554E2DE",
    x"3554C844",
    x"3554ADAC",
    x"35549318",
    x"35547887",
    x"35545DFA",
    x"35544370",
    x"355428E9",
    x"35540E66",
    x"3553F3E6",
    x"3553D969",
    x"3553BEEF",
    x"3553A479",
    x"35538A06",
    x"35536F97",
    x"3553552A",
    x"35533AC1",
    x"3553205C",
    x"355305F9",
    x"3552EB9A",
    x"3552D13E",
    x"3552B6E6",
    x"35529C91",
    x"3552823F",
    x"355267F0",
    x"35524DA5",
    x"3552335D",
    x"35521918",
    x"3551FED6",
    x"3551E498",
    x"3551CA5D",
    x"3551B025",
    x"355195F1",
    x"35517BC0",
    x"35516192",
    x"35514768",
    x"35512D40",
    x"3551131C",
    x"3550F8FC",
    x"3550DEDE",
    x"3550C4C4",
    x"3550AAAD",
    x"35509099",
    x"35507689",
    x"35505C7C",
    x"35504272",
    x"3550286B",
    x"35500E67",
    x"354FF467",
    x"354FDA6A",
    x"354FC071",
    x"354FA67A",
    x"354F8C87",
    x"354F7297",
    x"354F58AA",
    x"354F3EC1",
    x"354F24DB",
    x"354F0AF8",
    x"354EF118",
    x"354ED73B",
    x"354EBD62",
    x"354EA38C",
    x"354E89B9",
    x"354E6FEA",
    x"354E561D",
    x"354E3C54",
    x"354E228E",
    x"354E08CC",
    x"354DEF0C",
    x"354DD550",
    x"354DBB97",
    x"354DA1E1",
    x"354D882E",
    x"354D6E7F",
    x"354D54D3",
    x"354D3B2A",
    x"354D2184",
    x"354D07E1",
    x"354CEE42",
    x"354CD4A6",
    x"354CBB0D",
    x"354CA177",
    x"354C87E4",
    x"354C6E55",
    x"354C54C9",
    x"354C3B40",
    x"354C21BA",
    x"354C0837",
    x"354BEEB8",
    x"354BD53C",
    x"354BBBC3",
    x"354BA24D",
    x"354B88DA",
    x"354B6F6A",
    x"354B55FE",
    x"354B3C95",
    x"354B232F",
    x"354B09CC",
    x"354AF06D",
    x"354AD710",
    x"354ABDB7",
    x"354AA461",
    x"354A8B0E",
    x"354A71BE",
    x"354A5871",
    x"354A3F28",
    x"354A25E1",
    x"354A0C9E",
    x"3549F35E",
    x"3549DA21",
    x"3549C0E8",
    x"3549A7B1",
    x"35498E7E",
    x"3549754E",
    x"35495C21",
    x"354942F7",
    x"354929D0",
    x"354910AC",
    x"3548F78C",
    x"3548DE6E",
    x"3548C554",
    x"3548AC3D",
    x"35489329",
    x"35487A18",
    x"3548610A",
    x"35484800",
    x"35482EF8",
    x"354815F4",
    x"3547FCF3",
    x"3547E3F5",
    x"3547CAFA",
    x"3547B202",
    x"3547990D",
    x"3547801C",
    x"3547672D",
    x"35474E42",
    x"3547355A",
    x"35471C75",
    x"35470393",
    x"3546EAB4",
    x"3546D1D8",
    x"3546B8FF",
    x"3546A02A",
    x"35468757",
    x"35466E88",
    x"354655BC",
    x"35463CF3",
    x"3546242C",
    x"35460B69",
    x"3545F2AA",
    x"3545D9ED",
    x"3545C133",
    x"3545A87D",
    x"35458FC9",
    x"35457719",
    x"35455E6B",
    x"354545C1",
    x"35452D1A",
    x"35451476",
    x"3544FBD5",
    x"3544E337",
    x"3544CA9C",
    x"3544B204",
    x"3544996F",
    x"354480DE",
    x"3544684F",
    x"35444FC4",
    x"3544373B",
    x"35441EB6",
    x"35440634",
    x"3543EDB4",
    x"3543D538",
    x"3543BCBF",
    x"3543A449",
    x"35438BD6",
    x"35437366",
    x"35435AF9",
    x"3543428F",
    x"35432A28",
    x"354311C5",
    x"3542F964",
    x"3542E106",
    x"3542C8AC",
    x"3542B054",
    x"35429800",
    x"35427FAE",
    x"35426760",
    x"35424F14",
    x"354236CC",
    x"35421E87",
    x"35420644",
    x"3541EE05",
    x"3541D5C9",
    x"3541BD90",
    x"3541A559",
    x"35418D26",
    x"354174F6",
    x"35415CC9",
    x"3541449F",
    x"35412C78",
    x"35411454",
    x"3540FC33",
    x"3540E415",
    x"3540CBFA",
    x"3540B3E2",
    x"35409BCD",
    x"354083BB",
    x"35406BAC",
    x"354053A0",
    x"35403B97",
    x"35402391",
    x"35400B8E",
    x"353FF38E",
    x"353FDB91",
    x"353FC397",
    x"353FABA0",
    x"353F93AC",
    x"353F7BBB",
    x"353F63CD",
    x"353F4BE2",
    x"353F33FA",
    x"353F1C15",
    x"353F0433",
    x"353EEC54",
    x"353ED478",
    x"353EBC9F",
    x"353EA4C9",
    x"353E8CF6",
    x"353E7526",
    x"353E5D59",
    x"353E458F",
    x"353E2DC7",
    x"353E1603",
    x"353DFE42",
    x"353DE684",
    x"353DCEC8",
    x"353DB710",
    x"353D9F5A",
    x"353D87A8",
    x"353D6FF9",
    x"353D584C",
    x"353D40A2",
    x"353D28FC",
    x"353D1158",
    x"353CF9B8",
    x"353CE21A",
    x"353CCA7F",
    x"353CB2E7",
    x"353C9B52",
    x"353C83C0",
    x"353C6C31",
    x"353C54A5",
    x"353C3D1C",
    x"353C2596",
    x"353C0E13",
    x"353BF693",
    x"353BDF15",
    x"353BC79B",
    x"353BB023",
    x"353B98AF",
    x"353B813D",
    x"353B69CE",
    x"353B5263",
    x"353B3AFA",
    x"353B2394",
    x"353B0C31",
    x"353AF4D1",
    x"353ADD74",
    x"353AC619",
    x"353AAEC2",
    x"353A976E",
    x"353A801C",
    x"353A68CE",
    x"353A5182",
    x"353A3A39",
    x"353A22F4",
    x"353A0BB1",
    x"3539F471",
    x"3539DD34",
    x"3539C5F9",
    x"3539AEC2",
    x"3539978E",
    x"3539805C",
    x"3539692E",
    x"35395202",
    x"35393AD9",
    x"353923B3",
    x"35390C90",
    x"3538F570",
    x"3538DE53",
    x"3538C738",
    x"3538B021",
    x"3538990C",
    x"353881FB",
    x"35386AEC",
    x"353853E0",
    x"35383CD7",
    x"353825D1",
    x"35380ECD",
    x"3537F7CD",
    x"3537E0D0",
    x"3537C9D5",
    x"3537B2DD",
    x"35379BE8",
    x"353784F6",
    x"35376E07",
    x"3537571B",
    x"35374031",
    x"3537294B",
    x"35371267",
    x"3536FB86",
    x"3536E4A8",
    x"3536CDCD",
    x"3536B6F4",
    x"3536A01F",
    x"3536894C",
    x"3536727D",
    x"35365BB0",
    x"353644E6",
    x"35362E1F",
    x"3536175A",
    x"35360099",
    x"3535E9DA",
    x"3535D31E",
    x"3535BC65",
    x"3535A5AF",
    x"35358EFC",
    x"3535784B",
    x"3535619E",
    x"35354AF3",
    x"3535344B",
    x"35351DA6",
    x"35350704",
    x"3534F064",
    x"3534D9C8",
    x"3534C32E",
    x"3534AC97",
    x"35349603",
    x"35347F71",
    x"353468E3",
    x"35345257",
    x"35343BCE",
    x"35342548",
    x"35340EC5",
    x"3533F844",
    x"3533E1C7",
    x"3533CB4C",
    x"3533B4D4",
    x"35339E5F",
    x"353387EC",
    x"3533717D",
    x"35335B10",
    x"353344A6",
    x"35332E3F",
    x"353317DA",
    x"35330179",
    x"3532EB1A",
    x"3532D4BE",
    x"3532BE65",
    x"3532A80E",
    x"353291BB",
    x"35327B6A",
    x"3532651C",
    x"35324ED1",
    x"35323888",
    x"35322243",
    x"35320C00",
    x"3531F5C0",
    x"3531DF82",
    x"3531C948",
    x"3531B310",
    x"35319CDB",
    x"353186A9",
    x"35317079",
    x"35315A4D",
    x"35314423",
    x"35312DFC",
    x"353117D7",
    x"353101B6",
    x"3530EB97",
    x"3530D57B",
    x"3530BF61",
    x"3530A94B",
    x"35309337",
    x"35307D26",
    x"35306718",
    x"3530510C",
    x"35303B04",
    x"353024FE",
    x"35300EFA",
    x"352FF8FA",
    x"352FE2FC",
    x"352FCD01",
    x"352FB709",
    x"352FA113",
    x"352F8B21",
    x"352F7531",
    x"352F5F43",
    x"352F4959",
    x"352F3371",
    x"352F1D8C",
    x"352F07AA",
    x"352EF1CA",
    x"352EDBED",
    x"352EC613",
    x"352EB03C",
    x"352E9A67",
    x"352E8495",
    x"352E6EC6",
    x"352E58F9",
    x"352E4330",
    x"352E2D68",
    x"352E17A4",
    x"352E01E3",
    x"352DEC24",
    x"352DD668",
    x"352DC0AE",
    x"352DAAF7",
    x"352D9543",
    x"352D7F92",
    x"352D69E3",
    x"352D5438",
    x"352D3E8E",
    x"352D28E8",
    x"352D1344",
    x"352CFDA3",
    x"352CE805",
    x"352CD269",
    x"352CBCD0",
    x"352CA73A",
    x"352C91A6",
    x"352C7C16",
    x"352C6687",
    x"352C50FC",
    x"352C3B73",
    x"352C25ED",
    x"352C106A",
    x"352BFAE9",
    x"352BE56B",
    x"352BCFF0",
    x"352BBA77",
    x"352BA501",
    x"352B8F8E",
    x"352B7A1D",
    x"352B64AF",
    x"352B4F44",
    x"352B39DB",
    x"352B2475",
    x"352B0F12",
    x"352AF9B2",
    x"352AE454",
    x"352ACEF9",
    x"352AB9A0",
    x"352AA44A",
    x"352A8EF7",
    x"352A79A6",
    x"352A6459",
    x"352A4F0D",
    x"352A39C5",
    x"352A247F",
    x"352A0F3C",
    x"3529F9FB",
    x"3529E4BD",
    x"3529CF82",
    x"3529BA49",
    x"3529A513",
    x"35298FE0",
    x"35297AAF",
    x"35296581",
    x"35295056",
    x"35293B2D",
    x"35292607",
    x"352910E4",
    x"3528FBC3",
    x"3528E6A5",
    x"3528D189",
    x"3528BC70",
    x"3528A75A",
    x"35289247",
    x"35287D36",
    x"35286827",
    x"3528531C",
    x"35283E13",
    x"3528290C",
    x"35281408",
    x"3527FF07",
    x"3527EA08",
    x"3527D50D",
    x"3527C013",
    x"3527AB1D",
    x"35279628",
    x"35278137",
    x"35276C48",
    x"3527575C",
    x"35274272",
    x"35272D8B",
    x"352718A7",
    x"352703C5",
    x"3526EEE6",
    x"3526DA09",
    x"3526C52F",
    x"3526B058",
    x"35269B83",
    x"352686B1",
    x"352671E2",
    x"35265D15",
    x"3526484A",
    x"35263383",
    x"35261EBE",
    x"352609FB",
    x"3525F53B",
    x"3525E07E",
    x"3525CBC3",
    x"3525B70B",
    x"3525A255",
    x"35258DA2",
    x"352578F2",
    x"35256444",
    x"35254F99",
    x"35253AF0",
    x"3525264A",
    x"352511A6",
    x"3524FD06",
    x"3524E867",
    x"3524D3CB",
    x"3524BF32",
    x"3524AA9C",
    x"35249608",
    x"35248176",
    x"35246CE7",
    x"3524585B",
    x"352443D1",
    x"35242F4A",
    x"35241AC5",
    x"35240643",
    x"3523F1C4",
    x"3523DD47",
    x"3523C8CC",
    x"3523B455",
    x"35239FDF",
    x"35238B6D",
    x"352376FD",
    x"3523628F",
    x"35234E24",
    x"352339BB",
    x"35232555",
    x"352310F2",
    x"3522FC91",
    x"3522E833",
    x"3522D3D7",
    x"3522BF7E",
    x"3522AB27",
    x"352296D3",
    x"35228282",
    x"35226E33",
    x"352259E6",
    x"3522459C",
    x"35223155",
    x"35221D10",
    x"352208CD",
    x"3521F48E",
    x"3521E050",
    x"3521CC15",
    x"3521B7DD",
    x"3521A3A7",
    x"35218F74",
    x"35217B44",
    x"35216715",
    x"352152EA",
    x"35213EC1",
    x"35212A9A",
    x"35211676",
    x"35210255",
    x"3520EE35",
    x"3520DA19",
    x"3520C5FF",
    x"3520B1E7",
    x"35209DD2",
    x"352089C0",
    x"352075B0",
    x"352061A3",
    x"35204D98",
    x"3520398F",
    x"35202589",
    x"35201186",
    x"351FFD85",
    x"351FE986",
    x"351FD58A",
    x"351FC191",
    x"351FAD9A",
    x"351F99A6",
    x"351F85B4",
    x"351F71C4",
    x"351F5DD7",
    x"351F49ED",
    x"351F3605",
    x"351F221F",
    x"351F0E3C",
    x"351EFA5C",
    x"351EE67E",
    x"351ED2A2",
    x"351EBEC9",
    x"351EAAF2",
    x"351E971E",
    x"351E834D",
    x"351E6F7D",
    x"351E5BB1",
    x"351E47E7",
    x"351E341F",
    x"351E2059",
    x"351E0C97",
    x"351DF8D6",
    x"351DE518",
    x"351DD15D",
    x"351DBDA4",
    x"351DA9EE",
    x"351D963A",
    x"351D8288",
    x"351D6ED9",
    x"351D5B2C",
    x"351D4782",
    x"351D33DA",
    x"351D2035",
    x"351D0C92",
    x"351CF8F2",
    x"351CE554",
    x"351CD1B9",
    x"351CBE20",
    x"351CAA89",
    x"351C96F5",
    x"351C8363",
    x"351C6FD4",
    x"351C5C48",
    x"351C48BD",
    x"351C3535",
    x"351C21B0",
    x"351C0E2D",
    x"351BFAAC",
    x"351BE72E",
    x"351BD3B3",
    x"351BC039",
    x"351BACC3",
    x"351B994E",
    x"351B85DC",
    x"351B726D",
    x"351B5F00",
    x"351B4B95",
    x"351B382D",
    x"351B24C7",
    x"351B1163",
    x"351AFE03",
    x"351AEAA4",
    x"351AD748",
    x"351AC3EE",
    x"351AB097",
    x"351A9D42",
    x"351A89F0",
    x"351A76A0",
    x"351A6352",
    x"351A5007",
    x"351A3CBE",
    x"351A2978",
    x"351A1634",
    x"351A02F2",
    x"3519EFB3",
    x"3519DC76",
    x"3519C93C",
    x"3519B604",
    x"3519A2CE",
    x"35198F9B",
    x"35197C6A",
    x"3519693C",
    x"35195610",
    x"351942E6",
    x"35192FBF",
    x"35191C9A",
    x"35190978",
    x"3518F658",
    x"3518E33B",
    x"3518D01F",
    x"3518BD06",
    x"3518A9F0",
    x"351896DC",
    x"351883CA",
    x"351870BB",
    x"35185DAE",
    x"35184AA4",
    x"3518379B",
    x"35182496",
    x"35181192",
    x"3517FE91",
    x"3517EB93",
    x"3517D896",
    x"3517C59D",
    x"3517B2A5",
    x"35179FB0",
    x"35178CBD",
    x"351779CD",
    x"351766DF",
    x"351753F3",
    x"3517410A",
    x"35172E23",
    x"35171B3E",
    x"3517085C",
    x"3516F57C",
    x"3516E29F",
    x"3516CFC3",
    x"3516BCEB",
    x"3516AA14",
    x"35169740",
    x"3516846E",
    x"3516719F",
    x"35165ED2",
    x"35164C07",
    x"3516393F",
    x"35162679",
    x"351613B5",
    x"351600F4",
    x"3515EE35",
    x"3515DB78",
    x"3515C8BE",
    x"3515B606",
    x"3515A351",
    x"3515909D",
    x"35157DED",
    x"35156B3E",
    x"35155892",
    x"351545E8",
    x"35153340",
    x"3515209B",
    x"35150DF8",
    x"3514FB58",
    x"3514E8B9",
    x"3514D61D",
    x"3514C384",
    x"3514B0EC",
    x"35149E58",
    x"35148BC5",
    x"35147935",
    x"351466A7",
    x"3514541B",
    x"35144192",
    x"35142F0B",
    x"35141C86",
    x"35140A03",
    x"3513F783",
    x"3513E506",
    x"3513D28A",
    x"3513C011",
    x"3513AD9A",
    x"35139B25",
    x"351388B3",
    x"35137643",
    x"351363D6",
    x"3513516A",
    x"35133F01",
    x"35132C9B",
    x"35131A36",
    x"351307D4",
    x"3512F574",
    x"3512E317",
    x"3512D0BB",
    x"3512BE62",
    x"3512AC0C",
    x"351299B7",
    x"35128765",
    x"35127516",
    x"351262C8",
    x"3512507D",
    x"35123E34",
    x"35122BED",
    x"351219A9",
    x"35120767",
    x"3511F527",
    x"3511E2EA",
    x"3511D0AE",
    x"3511BE76",
    x"3511AC3F",
    x"35119A0A",
    x"351187D8",
    x"351175A8",
    x"3511637B",
    x"35115150",
    x"35113F27",
    x"35112D00",
    x"35111ADB",
    x"351108B9",
    x"3510F699",
    x"3510E47B",
    x"3510D260",
    x"3510C047",
    x"3510AE30",
    x"35109C1B",
    x"35108A09",
    x"351077F9",
    x"351065EB",
    x"351053DF",
    x"351041D6",
    x"35102FCF",
    x"35101DCA",
    x"35100BC7",
    x"350FF9C7",
    x"350FE7C9",
    x"350FD5CD",
    x"350FC3D4",
    x"350FB1DC",
    x"350F9FE7",
    x"350F8DF4",
    x"350F7C04",
    x"350F6A15",
    x"350F5829",
    x"350F463F",
    x"350F3457",
    x"350F2272",
    x"350F108F",
    x"350EFEAE",
    x"350EECCF",
    x"350EDAF3",
    x"350EC918",
    x"350EB740",
    x"350EA56B",
    x"350E9397",
    x"350E81C6",
    x"350E6FF7",
    x"350E5E2A",
    x"350E4C5F",
    x"350E3A97",
    x"350E28D0",
    x"350E170C",
    x"350E054B",
    x"350DF38B",
    x"350DE1CE",
    x"350DD013",
    x"350DBE5A",
    x"350DACA3",
    x"350D9AEF",
    x"350D893C",
    x"350D778C",
    x"350D65DE",
    x"350D5433",
    x"350D4289",
    x"350D30E2",
    x"350D1F3D",
    x"350D0D9A",
    x"350CFBFA",
    x"350CEA5B",
    x"350CD8BF",
    x"350CC725",
    x"350CB58D",
    x"350CA3F8",
    x"350C9264",
    x"350C80D3",
    x"350C6F44",
    x"350C5DB7",
    x"350C4C2D",
    x"350C3AA4",
    x"350C291E",
    x"350C179A",
    x"350C0618",
    x"350BF499",
    x"350BE31B",
    x"350BD1A0",
    x"350BC027",
    x"350BAEB0",
    x"350B9D3B",
    x"350B8BC8",
    x"350B7A58",
    x"350B68EA",
    x"350B577E",
    x"350B4614",
    x"350B34AC",
    x"350B2347",
    x"350B11E4",
    x"350B0082",
    x"350AEF23",
    x"350ADDC7",
    x"350ACC6C",
    x"350ABB13",
    x"350AA9BD",
    x"350A9869",
    x"350A8717",
    x"350A75C7",
    x"350A647A",
    x"350A532E",
    x"350A41E5",
    x"350A309E",
    x"350A1F59",
    x"350A0E16",
    x"3509FCD5",
    x"3509EB97",
    x"3509DA5A",
    x"3509C920",
    x"3509B7E8",
    x"3509A6B2",
    x"3509957E",
    x"3509844D",
    x"3509731D",
    x"350961F0",
    x"350950C5",
    x"35093F9C",
    x"35092E75",
    x"35091D50",
    x"35090C2E",
    x"3508FB0D",
    x"3508E9EF",
    x"3508D8D3",
    x"3508C7B9",
    x"3508B6A1",
    x"3508A58B",
    x"35089477",
    x"35088366",
    x"35087256",
    x"35086149",
    x"3508503E",
    x"35083F35",
    x"35082E2E",
    x"35081D2A",
    x"35080C27",
    x"3507FB27",
    x"3507EA28",
    x"3507D92C",
    x"3507C832",
    x"3507B73A",
    x"3507A644",
    x"35079550",
    x"3507845F",
    x"3507736F",
    x"35076282",
    x"35075197",
    x"350740AE",
    x"35072FC6",
    x"35071EE2",
    x"35070DFF",
    x"3506FD1E",
    x"3506EC3F",
    x"3506DB63",
    x"3506CA89",
    x"3506B9B0",
    x"3506A8DA",
    x"35069806",
    x"35068734",
    x"35067664",
    x"35066597",
    x"350654CB",
    x"35064401",
    x"3506333A",
    x"35062275",
    x"350611B1",
    x"350600F0",
    x"3505F031",
    x"3505DF74",
    x"3505CEB9",
    x"3505BE00",
    x"3505AD4A",
    x"35059C95",
    x"35058BE3",
    x"35057B32",
    x"35056A84",
    x"350559D8",
    x"3505492D",
    x"35053885",
    x"350527DF",
    x"3505173B",
    x"35050699",
    x"3504F5FA",
    x"3504E55C",
    x"3504D4C0",
    x"3504C427",
    x"3504B38F",
    x"3504A2FA",
    x"35049266",
    x"350481D5",
    x"35047146",
    x"350460B9",
    x"3504502E",
    x"35043FA5",
    x"35042F1E",
    x"35041E99",
    x"35040E16",
    x"3503FD96",
    x"3503ED17",
    x"3503DC9A",
    x"3503CC20",
    x"3503BBA7",
    x"3503AB31",
    x"35039ABC",
    x"35038A4A",
    x"350379DA",
    x"3503696C",
    x"35035900",
    x"35034895",
    x"3503382D",
    x"350327C7",
    x"35031763",
    x"35030702",
    x"3502F6A2",
    x"3502E644",
    x"3502D5E8",
    x"3502C58E",
    x"3502B537",
    x"3502A4E1",
    x"3502948E",
    x"3502843C",
    x"350273EC",
    x"3502639F",
    x"35025354",
    x"3502430A",
    x"350232C3",
    x"3502227D",
    x"3502123A",
    x"350201F9",
    x"3501F1BA",
    x"3501E17C",
    x"3501D141",
    x"3501C108",
    x"3501B0D1",
    x"3501A09C",
    x"35019069",
    x"35018038",
    x"35017009",
    x"35015FDC",
    x"35014FB1",
    x"35013F88",
    x"35012F61",
    x"35011F3C",
    x"35010F19",
    x"3500FEF8",
    x"3500EED9",
    x"3500DEBD",
    x"3500CEA2",
    x"3500BE89",
    x"3500AE72",
    x"35009E5D",
    x"35008E4B",
    x"35007E3A",
    x"35006E2B",
    x"35005E1E",
    x"35004E13",
    x"35003E0B",
    x"35002E04",
    x"35001DFF",
    x"35000DFC",
    x"34FFFBF7",
    x"34FFDBFA",
    x"34FFBC00",
    x"34FF9C0B",
    x"34FF7C19",
    x"34FF5C2C",
    x"34FF3C42",
    x"34FF1C5D",
    x"34FEFC7B",
    x"34FEDC9E",
    x"34FEBCC4",
    x"34FE9CEE",
    x"34FE7D1D",
    x"34FE5D4F",
    x"34FE3D86",
    x"34FE1DC0",
    x"34FDFDFE",
    x"34FDDE40",
    x"34FDBE87",
    x"34FD9ED1",
    x"34FD7F1F",
    x"34FD5F71",
    x"34FD3FC7",
    x"34FD2021",
    x"34FD007F",
    x"34FCE0E1",
    x"34FCC147",
    x"34FCA1B0",
    x"34FC821E",
    x"34FC6290",
    x"34FC4306",
    x"34FC237F",
    x"34FC03FD",
    x"34FBE47E",
    x"34FBC504",
    x"34FBA58D",
    x"34FB861A",
    x"34FB66AB",
    x"34FB4741",
    x"34FB27DA",
    x"34FB0877",
    x"34FAE918",
    x"34FAC9BC",
    x"34FAAA65",
    x"34FA8B12",
    x"34FA6BC2",
    x"34FA4C77",
    x"34FA2D2F",
    x"34FA0DEB",
    x"34F9EEAC",
    x"34F9CF70",
    x"34F9B038",
    x"34F99104",
    x"34F971D4",
    x"34F952A7",
    x"34F9337F",
    x"34F9145A",
    x"34F8F53A",
    x"34F8D61D",
    x"34F8B704",
    x"34F897EF",
    x"34F878DE",
    x"34F859D1",
    x"34F83AC8",
    x"34F81BC2",
    x"34F7FCC1",
    x"34F7DDC3",
    x"34F7BEC9",
    x"34F79FD4",
    x"34F780E2",
    x"34F761F3",
    x"34F74309",
    x"34F72423",
    x"34F70540",
    x"34F6E661",
    x"34F6C786",
    x"34F6A8AF",
    x"34F689DC",
    x"34F66B0D",
    x"34F64C41",
    x"34F62D7A",
    x"34F60EB6",
    x"34F5EFF6",
    x"34F5D13A",
    x"34F5B282",
    x"34F593CD",
    x"34F5751D",
    x"34F55670",
    x"34F537C7",
    x"34F51922",
    x"34F4FA81",
    x"34F4DBE4",
    x"34F4BD4A",
    x"34F49EB4",
    x"34F48022",
    x"34F46194",
    x"34F4430A",
    x"34F42484",
    x"34F40601",
    x"34F3E782",
    x"34F3C907",
    x"34F3AA90",
    x"34F38C1C",
    x"34F36DAD",
    x"34F34F41",
    x"34F330D9",
    x"34F31275",
    x"34F2F414",
    x"34F2D5B8",
    x"34F2B75F",
    x"34F2990A",
    x"34F27AB9",
    x"34F25C6B",
    x"34F23E22",
    x"34F21FDC",
    x"34F2019A",
    x"34F1E35B",
    x"34F1C521",
    x"34F1A6EA",
    x"34F188B7",
    x"34F16A88",
    x"34F14C5C",
    x"34F12E35",
    x"34F11011",
    x"34F0F1F1",
    x"34F0D3D4",
    x"34F0B5BC",
    x"34F097A7",
    x"34F07996",
    x"34F05B88",
    x"34F03D7F",
    x"34F01F79",
    x"34F00177",
    x"34EFE379",
    x"34EFC57E",
    x"34EFA787",
    x"34EF8994",
    x"34EF6BA5",
    x"34EF4DB9",
    x"34EF2FD2",
    x"34EF11ED",
    x"34EEF40D",
    x"34EED630",
    x"34EEB858",
    x"34EE9A82",
    x"34EE7CB1",
    x"34EE5EE3",
    x"34EE4119",
    x"34EE2353",
    x"34EE0590",
    x"34EDE7D1",
    x"34EDCA16",
    x"34EDAC5F",
    x"34ED8EAB",
    x"34ED70FB",
    x"34ED534F",
    x"34ED35A6",
    x"34ED1802",
    x"34ECFA60",
    x"34ECDCC3",
    x"34ECBF29",
    x"34ECA193",
    x"34EC8401",
    x"34EC6672",
    x"34EC48E7",
    x"34EC2B60",
    x"34EC0DDC",
    x"34EBF05D",
    x"34EBD2E0",
    x"34EBB568",
    x"34EB97F3",
    x"34EB7A82",
    x"34EB5D14",
    x"34EB3FAB",
    x"34EB2244",
    x"34EB04E2",
    x"34EAE783",
    x"34EACA28",
    x"34EAACD1",
    x"34EA8F7D",
    x"34EA722D",
    x"34EA54E0",
    x"34EA3798",
    x"34EA1A52",
    x"34E9FD11",
    x"34E9DFD3",
    x"34E9C299",
    x"34E9A563",
    x"34E98830",
    x"34E96B00",
    x"34E94DD5",
    x"34E930AD",
    x"34E91389",
    x"34E8F668",
    x"34E8D94B",
    x"34E8BC32",
    x"34E89F1C",
    x"34E8820A",
    x"34E864FC",
    x"34E847F1",
    x"34E82AEA",
    x"34E80DE6",
    x"34E7F0E6",
    x"34E7D3EA",
    x"34E7B6F1",
    x"34E799FC",
    x"34E77D0B",
    x"34E7601D",
    x"34E74333",
    x"34E7264C",
    x"34E70969",
    x"34E6EC8A",
    x"34E6CFAE",
    x"34E6B2D6",
    x"34E69601",
    x"34E67930",
    x"34E65C63",
    x"34E63F99",
    x"34E622D3",
    x"34E60610",
    x"34E5E952",
    x"34E5CC96",
    x"34E5AFDE",
    x"34E5932A",
    x"34E5767A",
    x"34E559CD",
    x"34E53D23",
    x"34E5207D",
    x"34E503DB",
    x"34E4E73C",
    x"34E4CAA1",
    x"34E4AE0A",
    x"34E49176",
    x"34E474E5",
    x"34E45858",
    x"34E43BCF",
    x"34E41F4A",
    x"34E402C7",
    x"34E3E649",
    x"34E3C9CE",
    x"34E3AD56",
    x"34E390E2",
    x"34E37472",
    x"34E35805",
    x"34E33B9C",
    x"34E31F36",
    x"34E302D4",
    x"34E2E676",
    x"34E2CA1B",
    x"34E2ADC3",
    x"34E2916F",
    x"34E2751F",
    x"34E258D2",
    x"34E23C89",
    x"34E22043",
    x"34E20401",
    x"34E1E7C2",
    x"34E1CB87",
    x"34E1AF4F",
    x"34E1931B",
    x"34E176EA",
    x"34E15ABD",
    x"34E13E94",
    x"34E1226D",
    x"34E1064B",
    x"34E0EA2C",
    x"34E0CE10",
    x"34E0B1F8",
    x"34E095E4",
    x"34E079D3",
    x"34E05DC5",
    x"34E041BB",
    x"34E025B5",
    x"34E009B2",
    x"34DFEDB3",
    x"34DFD1B7",
    x"34DFB5BE",
    x"34DF99C9",
    x"34DF7DD8",
    x"34DF61EA",
    x"34DF45FF",
    x"34DF2A18",
    x"34DF0E35",
    x"34DEF255",
    x"34DED678",
    x"34DEBA9F",
    x"34DE9EC9",
    x"34DE82F7",
    x"34DE6729",
    x"34DE4B5E",
    x"34DE2F96",
    x"34DE13D2",
    x"34DDF811",
    x"34DDDC54",
    x"34DDC09A",
    x"34DDA4E3",
    x"34DD8931",
    x"34DD6D81",
    x"34DD51D5",
    x"34DD362D",
    x"34DD1A88",
    x"34DCFEE6",
    x"34DCE348",
    x"34DCC7AD",
    x"34DCAC16",
    x"34DC9082",
    x"34DC74F2",
    x"34DC5965",
    x"34DC3DDC",
    x"34DC2256",
    x"34DC06D3",
    x"34DBEB54",
    x"34DBCFD8",
    x"34DBB460",
    x"34DB98EB",
    x"34DB7D7A",
    x"34DB620C",
    x"34DB46A1",
    x"34DB2B3A",
    x"34DB0FD6",
    x"34DAF476",
    x"34DAD919",
    x"34DABDC0",
    x"34DAA26A",
    x"34DA8717",
    x"34DA6BC8",
    x"34DA507C",
    x"34DA3534",
    x"34DA19EF",
    x"34D9FEAD",
    x"34D9E36F",
    x"34D9C835",
    x"34D9ACFD",
    x"34D991C9",
    x"34D97699",
    x"34D95B6C",
    x"34D94042",
    x"34D9251C",
    x"34D909F9",
    x"34D8EED9",
    x"34D8D3BD",
    x"34D8B8A4",
    x"34D89D8F",
    x"34D8827D",
    x"34D8676E",
    x"34D84C63",
    x"34D8315B",
    x"34D81657",
    x"34D7FB55",
    x"34D7E058",
    x"34D7C55D",
    x"34D7AA66",
    x"34D78F73",
    x"34D77483",
    x"34D75996",
    x"34D73EAC",
    x"34D723C6",
    x"34D708E3",
    x"34D6EE04",
    x"34D6D328",
    x"34D6B84F",
    x"34D69D7A",
    x"34D682A8",
    x"34D667D9",
    x"34D64D0E",
    x"34D63246",
    x"34D61781",
    x"34D5FCC0",
    x"34D5E202",
    x"34D5C747",
    x"34D5AC90",
    x"34D591DC",
    x"34D5772C",
    x"34D55C7E",
    x"34D541D4",
    x"34D5272E",
    x"34D50C8B",
    x"34D4F1EB",
    x"34D4D74E",
    x"34D4BCB5",
    x"34D4A21F",
    x"34D4878C",
    x"34D46CFD",
    x"34D45271",
    x"34D437E8",
    x"34D41D63",
    x"34D402E1",
    x"34D3E862",
    x"34D3CDE7",
    x"34D3B36F",
    x"34D398FA",
    x"34D37E89",
    x"34D3641B",
    x"34D349B0",
    x"34D32F48",
    x"34D314E4",
    x"34D2FA83",
    x"34D2E025",
    x"34D2C5CB",
    x"34D2AB74",
    x"34D29120",
    x"34D276D0",
    x"34D25C82",
    x"34D24238",
    x"34D227F2",
    x"34D20DAE",
    x"34D1F36E",
    x"34D1D932",
    x"34D1BEF8",
    x"34D1A4C2",
    x"34D18A8F",
    x"34D1705F",
    x"34D15633",
    x"34D13C0A",
    x"34D121E4",
    x"34D107C1",
    x"34D0EDA2",
    x"34D0D386",
    x"34D0B96D",
    x"34D09F57",
    x"34D08545",
    x"34D06B36",
    x"34D0512A",
    x"34D03722",
    x"34D01D1D",
    x"34D0031A",
    x"34CFE91C",
    x"34CFCF20",
    x"34CFB528",
    x"34CF9B33",
    x"34CF8141",
    x"34CF6753",
    x"34CF4D67",
    x"34CF337F",
    x"34CF199A",
    x"34CEFFB9",
    x"34CEE5DB",
    x"34CECBFF",
    x"34CEB228",
    x"34CE9853",
    x"34CE7E81",
    x"34CE64B3",
    x"34CE4AE8",
    x"34CE3120",
    x"34CE175C",
    x"34CDFD9B",
    x"34CDE3DD",
    x"34CDCA22",
    x"34CDB06A",
    x"34CD96B6",
    x"34CD7D04",
    x"34CD6356",
    x"34CD49AC",
    x"34CD3004",
    x"34CD1660",
    x"34CCFCBE",
    x"34CCE320",
    x"34CCC986",
    x"34CCAFEE",
    x"34CC965A",
    x"34CC7CC8",
    x"34CC633A",
    x"34CC49B0",
    x"34CC3028",
    x"34CC16A4",
    x"34CBFD22",
    x"34CBE3A4",
    x"34CBCA29",
    x"34CBB0B2",
    x"34CB973D",
    x"34CB7DCC",
    x"34CB645E",
    x"34CB4AF3",
    x"34CB318B",
    x"34CB1826",
    x"34CAFEC5",
    x"34CAE567",
    x"34CACC0C",
    x"34CAB2B4",
    x"34CA995F",
    x"34CA800D",
    x"34CA66BF",
    x"34CA4D74",
    x"34CA342C",
    x"34CA1AE7",
    x"34CA01A5",
    x"34C9E866",
    x"34C9CF2B",
    x"34C9B5F2",
    x"34C99CBD",
    x"34C9838B",
    x"34C96A5C",
    x"34C95131",
    x"34C93808",
    x"34C91EE3",
    x"34C905C0",
    x"34C8ECA1",
    x"34C8D385",
    x"34C8BA6C",
    x"34C8A157",
    x"34C88844",
    x"34C86F35",
    x"34C85628",
    x"34C83D1F",
    x"34C82419",
    x"34C80B16",
    x"34C7F216",
    x"34C7D919",
    x"34C7C020",
    x"34C7A729",
    x"34C78E36",
    x"34C77546",
    x"34C75C59",
    x"34C7436F",
    x"34C72A88",
    x"34C711A4",
    x"34C6F8C3",
    x"34C6DFE6",
    x"34C6C70B",
    x"34C6AE34",
    x"34C69560",
    x"34C67C8F",
    x"34C663C1",
    x"34C64AF6",
    x"34C6322E",
    x"34C61969",
    x"34C600A8",
    x"34C5E7E9",
    x"34C5CF2E",
    x"34C5B675",
    x"34C59DC0",
    x"34C5850E",
    x"34C56C5F",
    x"34C553B3",
    x"34C53B0A",
    x"34C52264",
    x"34C509C1",
    x"34C4F122",
    x"34C4D885",
    x"34C4BFEC",
    x"34C4A755",
    x"34C48EC2",
    x"34C47631",
    x"34C45DA4",
    x"34C4451A",
    x"34C42C93",
    x"34C4140F",
    x"34C3FB8E",
    x"34C3E310",
    x"34C3CA95",
    x"34C3B21D",
    x"34C399A9",
    x"34C38137",
    x"34C368C8",
    x"34C3505D",
    x"34C337F4",
    x"34C31F8F",
    x"34C3072C",
    x"34C2EECD",
    x"34C2D671",
    x"34C2BE17",
    x"34C2A5C1",
    x"34C28D6E",
    x"34C2751E",
    x"34C25CD1",
    x"34C24486",
    x"34C22C3F",
    x"34C213FB",
    x"34C1FBBA",
    x"34C1E37C",
    x"34C1CB42",
    x"34C1B30A",
    x"34C19AD5",
    x"34C182A3",
    x"34C16A74",
    x"34C15248",
    x"34C13A20",
    x"34C121FA",
    x"34C109D7",
    x"34C0F1B7",
    x"34C0D99B",
    x"34C0C181",
    x"34C0A96A",
    x"34C09157",
    x"34C07946",
    x"34C06138",
    x"34C0492E",
    x"34C03126",
    x"34C01921",
    x"34C00120",
    x"34BFE921",
    x"34BFD125",
    x"34BFB92D",
    x"34BFA137",
    x"34BF8944",
    x"34BF7155",
    x"34BF5968",
    x"34BF417E",
    x"34BF2998",
    x"34BF11B4",
    x"34BEF9D3",
    x"34BEE1F6",
    x"34BECA1B",
    x"34BEB243",
    x"34BE9A6E",
    x"34BE829C",
    x"34BE6ACE",
    x"34BE5302",
    x"34BE3B39",
    x"34BE2373",
    x"34BE0BB0",
    x"34BDF3F0",
    x"34BDDC33",
    x"34BDC479",
    x"34BDACC2",
    x"34BD950E",
    x"34BD7D5D",
    x"34BD65AE",
    x"34BD4E03",
    x"34BD365B",
    x"34BD1EB6",
    x"34BD0713",
    x"34BCEF74",
    x"34BCD7D7",
    x"34BCC03E",
    x"34BCA8A7",
    x"34BC9114",
    x"34BC7983",
    x"34BC61F5",
    x"34BC4A6B",
    x"34BC32E3",
    x"34BC1B5E",
    x"34BC03DC",
    x"34BBEC5D",
    x"34BBD4E1",
    x"34BBBD68",
    x"34BBA5F1",
    x"34BB8E7E",
    x"34BB770E",
    x"34BB5FA0",
    x"34BB4836",
    x"34BB30CE",
    x"34BB196A",
    x"34BB0208",
    x"34BAEAA9",
    x"34BAD34D",
    x"34BABBF4",
    x"34BAA49E",
    x"34BA8D4B",
    x"34BA75FB",
    x"34BA5EAE",
    x"34BA4763",
    x"34BA301C",
    x"34BA18D7",
    x"34BA0196",
    x"34B9EA57",
    x"34B9D31B",
    x"34B9BBE2",
    x"34B9A4AC",
    x"34B98D79",
    x"34B97649",
    x"34B95F1B",
    x"34B947F1",
    x"34B930C9",
    x"34B919A5",
    x"34B90283",
    x"34B8EB64",
    x"34B8D448",
    x"34B8BD2F",
    x"34B8A619",
    x"34B88F06",
    x"34B877F5",
    x"34B860E8",
    x"34B849DD",
    x"34B832D5",
    x"34B81BD0",
    x"34B804CE",
    x"34B7EDCF",
    x"34B7D6D3",
    x"34B7BFD9",
    x"34B7A8E3",
    x"34B791EF",
    x"34B77AFE",
    x"34B76410",
    x"34B74D25",
    x"34B7363D",
    x"34B71F58",
    x"34B70875",
    x"34B6F196",
    x"34B6DAB9",
    x"34B6C3DF",
    x"34B6AD08",
    x"34B69634",
    x"34B67F62",
    x"34B66894",
    x"34B651C8",
    x"34B63AFF",
    x"34B62439",
    x"34B60D76",
    x"34B5F6B6",
    x"34B5DFF9",
    x"34B5C93E",
    x"34B5B286",
    x"34B59BD1",
    x"34B5851F",
    x"34B56E70",
    x"34B557C4",
    x"34B5411A",
    x"34B52A73",
    x"34B513D0",
    x"34B4FD2E",
    x"34B4E690",
    x"34B4CFF5",
    x"34B4B95C",
    x"34B4A2C7",
    x"34B48C34",
    x"34B475A3",
    x"34B45F16",
    x"34B4488C",
    x"34B43204",
    x"34B41B7F",
    x"34B404FD",
    x"34B3EE7E",
    x"34B3D802",
    x"34B3C188",
    x"34B3AB11",
    x"34B3949D",
    x"34B37E2C",
    x"34B367BE",
    x"34B35152",
    x"34B33AE9",
    x"34B32483",
    x"34B30E20",
    x"34B2F7C0",
    x"34B2E162",
    x"34B2CB07",
    x"34B2B4AF",
    x"34B29E5A",
    x"34B28808",
    x"34B271B8",
    x"34B25B6B",
    x"34B24521",
    x"34B22EDA",
    x"34B21896",
    x"34B20254",
    x"34B1EC15",
    x"34B1D5D9",
    x"34B1BFA0",
    x"34B1A969",
    x"34B19335",
    x"34B17D04",
    x"34B166D6",
    x"34B150AB",
    x"34B13A82",
    x"34B1245C",
    x"34B10E39",
    x"34B0F818",
    x"34B0E1FB",
    x"34B0CBE0",
    x"34B0B5C8",
    x"34B09FB2",
    x"34B089A0",
    x"34B07390",
    x"34B05D83",
    x"34B04779",
    x"34B03171",
    x"34B01B6C",
    x"34B0056A",
    x"34AFEF6B",
    x"34AFD96E",
    x"34AFC375",
    x"34AFAD7E",
    x"34AF9789",
    x"34AF8198",
    x"34AF6BA9",
    x"34AF55BD",
    x"34AF3FD3",
    x"34AF29ED",
    x"34AF1409",
    x"34AEFE28",
    x"34AEE849",
    x"34AED26E",
    x"34AEBC95",
    x"34AEA6BF",
    x"34AE90EB",
    x"34AE7B1A",
    x"34AE654C",
    x"34AE4F81",
    x"34AE39B8",
    x"34AE23F3",
    x"34AE0E2F",
    x"34ADF86F",
    x"34ADE2B1",
    x"34ADCCF6",
    x"34ADB73E",
    x"34ADA189",
    x"34AD8BD6",
    x"34AD7626",
    x"34AD6078",
    x"34AD4ACD",
    x"34AD3525",
    x"34AD1F80",
    x"34AD09DE",
    x"34ACF43E",
    x"34ACDEA1",
    x"34ACC906",
    x"34ACB36E",
    x"34AC9DD9",
    x"34AC8847",
    x"34AC72B7",
    x"34AC5D2A",
    x"34AC47A0",
    x"34AC3218",
    x"34AC1C93",
    x"34AC0711",
    x"34ABF192",
    x"34ABDC15",
    x"34ABC69B",
    x"34ABB123",
    x"34AB9BAE",
    x"34AB863C",
    x"34AB70CD",
    x"34AB5B60",
    x"34AB45F6",
    x"34AB308E",
    x"34AB1B2A",
    x"34AB05C8",
    x"34AAF068",
    x"34AADB0C",
    x"34AAC5B1",
    x"34AAB05A",
    x"34AA9B05",
    x"34AA85B3",
    x"34AA7064",
    x"34AA5B17",
    x"34AA45CD",
    x"34AA3086",
    x"34AA1B41",
    x"34AA05FF",
    x"34A9F0C0",
    x"34A9DB83",
    x"34A9C649",
    x"34A9B111",
    x"34A99BDC",
    x"34A986AA",
    x"34A9717B",
    x"34A95C4E",
    x"34A94724",
    x"34A931FC",
    x"34A91CD7",
    x"34A907B5",
    x"34A8F295",
    x"34A8DD78",
    x"34A8C85E",
    x"34A8B346",
    x"34A89E31",
    x"34A8891F",
    x"34A8740F",
    x"34A85F02",
    x"34A849F7",
    x"34A834EF",
    x"34A81FEA",
    x"34A80AE7",
    x"34A7F5E7",
    x"34A7E0EA",
    x"34A7CBEF",
    x"34A7B6F7",
    x"34A7A201",
    x"34A78D0E",
    x"34A7781E",
    x"34A76330",
    x"34A74E45",
    x"34A7395D",
    x"34A72477",
    x"34A70F93",
    x"34A6FAB3",
    x"34A6E5D5",
    x"34A6D0F9",
    x"34A6BC21",
    x"34A6A74A",
    x"34A69277",
    x"34A67DA6",
    x"34A668D7",
    x"34A6540B",
    x"34A63F42",
    x"34A62A7C",
    x"34A615B8",
    x"34A600F6",
    x"34A5EC37",
    x"34A5D77B",
    x"34A5C2C2",
    x"34A5AE0B",
    x"34A59956",
    x"34A584A4",
    x"34A56FF5",
    x"34A55B48",
    x"34A5469E",
    x"34A531F7",
    x"34A51D52",
    x"34A508AF",
    x"34A4F40F",
    x"34A4DF72",
    x"34A4CAD8",
    x"34A4B63F",
    x"34A4A1AA",
    x"34A48D17",
    x"34A47887",
    x"34A463F9",
    x"34A44F6E",
    x"34A43AE5",
    x"34A4265F",
    x"34A411DB",
    x"34A3FD5B",
    x"34A3E8DC",
    x"34A3D460",
    x"34A3BFE7",
    x"34A3AB70",
    x"34A396FC",
    x"34A3828B",
    x"34A36E1C",
    x"34A359AF",
    x"34A34545",
    x"34A330DE",
    x"34A31C79",
    x"34A30817",
    x"34A2F3B7",
    x"34A2DF5A",
    x"34A2CAFF",
    x"34A2B6A7",
    x"34A2A251",
    x"34A28DFE",
    x"34A279AE",
    x"34A26560",
    x"34A25115",
    x"34A23CCC",
    x"34A22885",
    x"34A21442",
    x"34A20000",
    x"34A1EBC2",
    x"34A1D785",
    x"34A1C34C",
    x"34A1AF15",
    x"34A19AE0",
    x"34A186AE",
    x"34A1727E",
    x"34A15E51",
    x"34A14A27",
    x"34A135FF",
    x"34A121D9",
    x"34A10DB6",
    x"34A0F996",
    x"34A0E578",
    x"34A0D15C",
    x"34A0BD43",
    x"34A0A92D",
    x"34A09519",
    x"34A08108",
    x"34A06CF9",
    x"34A058ED",
    x"34A044E3",
    x"34A030DB",
    x"34A01CD6",
    x"34A008D4",
    x"349FF4D4",
    x"349FE0D7",
    x"349FCCDC",
    x"349FB8E4",
    x"349FA4EE",
    x"349F90FA",
    x"349F7D0A",
    x"349F691B",
    x"349F552F",
    x"349F4146",
    x"349F2D5F",
    x"349F197B",
    x"349F0599",
    x"349EF1B9",
    x"349EDDDC",
    x"349ECA02",
    x"349EB62A",
    x"349EA254",
    x"349E8E81",
    x"349E7AB0",
    x"349E66E2",
    x"349E5317",
    x"349E3F4E",
    x"349E2B87",
    x"349E17C3",
    x"349E0401",
    x"349DF042",
    x"349DDC85",
    x"349DC8CB",
    x"349DB513",
    x"349DA15D",
    x"349D8DAA",
    x"349D79FA",
    x"349D664C",
    x"349D52A0",
    x"349D3EF7",
    x"349D2B51",
    x"349D17AC",
    x"349D040B",
    x"349CF06B",
    x"349CDCCF",
    x"349CC934",
    x"349CB59C",
    x"349CA207",
    x"349C8E74",
    x"349C7AE3",
    x"349C6755",
    x"349C53C9",
    x"349C4040",
    x"349C2CB9",
    x"349C1935",
    x"349C05B3",
    x"349BF233",
    x"349BDEB6",
    x"349BCB3C",
    x"349BB7C4",
    x"349BA44E",
    x"349B90DB",
    x"349B7D6A",
    x"349B69FB",
    x"349B568F",
    x"349B4326",
    x"349B2FBE",
    x"349B1C5A",
    x"349B08F7",
    x"349AF597",
    x"349AE23A",
    x"349ACEDF",
    x"349ABB86",
    x"349AA830",
    x"349A94DC",
    x"349A818B",
    x"349A6E3C",
    x"349A5AEF",
    x"349A47A5",
    x"349A345D",
    x"349A2118",
    x"349A0DD5",
    x"3499FA94",
    x"3499E756",
    x"3499D41B",
    x"3499C0E1",
    x"3499ADAA",
    x"34999A76",
    x"34998744",
    x"34997414",
    x"349960E7",
    x"34994DBC",
    x"34993A93",
    x"3499276D",
    x"34991449",
    x"34990128",
    x"3498EE09",
    x"3498DAED",
    x"3498C7D2",
    x"3498B4BB",
    x"3498A1A5",
    x"34988E92",
    x"34987B82",
    x"34986873",
    x"34985568",
    x"3498425E",
    x"34982F57",
    x"34981C52",
    x"34980950",
    x"3497F650",
    x"3497E352",
    x"3497D057",
    x"3497BD5E",
    x"3497AA68",
    x"34979774",
    x"34978482",
    x"34977192",
    x"34975EA5",
    x"34974BBB",
    x"349738D3",
    x"349725ED",
    x"34971309",
    x"34970028",
    x"3496ED49",
    x"3496DA6D",
    x"3496C792",
    x"3496B4BB",
    x"3496A1E5",
    x"34968F12",
    x"34967C41",
    x"34966973",
    x"349656A7",
    x"349643DD",
    x"34963116",
    x"34961E51",
    x"34960B8F",
    x"3495F8CE",
    x"3495E610",
    x"3495D355",
    x"3495C09B",
    x"3495ADE5",
    x"34959B30",
    x"3495887E",
    x"349575CE",
    x"34956320",
    x"34955075",
    x"34953DCC",
    x"34952B26",
    x"34951881",
    x"349505E0",
    x"3494F340",
    x"3494E0A3",
    x"3494CE08",
    x"3494BB6F",
    x"3494A8D9",
    x"34949645",
    x"349483B3",
    x"34947124",
    x"34945E97",
    x"34944C0C",
    x"34943984",
    x"349426FE",
    x"3494147A",
    x"349401F9",
    x"3493EF7A",
    x"3493DCFD",
    x"3493CA83",
    x"3493B80A",
    x"3493A595",
    x"34939321",
    x"349380B0",
    x"34936E41",
    x"34935BD4",
    x"3493496A",
    x"34933702",
    x"3493249C",
    x"34931239",
    x"3492FFD8",
    x"3492ED79",
    x"3492DB1C",
    x"3492C8C2",
    x"3492B66A",
    x"3492A414",
    x"349291C1",
    x"34927F70",
    x"34926D21",
    x"34925AD5",
    x"3492488A",
    x"34923643",
    x"349223FD",
    x"349211BA",
    x"3491FF78",
    x"3491ED3A",
    x"3491DAFD",
    x"3491C8C3",
    x"3491B68B",
    x"3491A455",
    x"34919222",
    x"34917FF1",
    x"34916DC2",
    x"34915B95",
    x"3491496B",
    x"34913743",
    x"3491251D",
    x"349112FA",
    x"349100D8",
    x"3490EEB9",
    x"3490DC9D",
    x"3490CA82",
    x"3490B86A",
    x"3490A654",
    x"34909441",
    x"3490822F",
    x"34907020",
    x"34905E13",
    x"34904C08",
    x"34903A00",
    x"349027FA",
    x"349015F6",
    x"349003F4",
    x"348FF1F5",
    x"348FDFF8",
    x"348FCDFD",
    x"348FBC04",
    x"348FAA0E",
    x"348F981A",
    x"348F8628",
    x"348F7438",
    x"348F624B",
    x"348F5060",
    x"348F3E77",
    x"348F2C90",
    x"348F1AAC",
    x"348F08CA",
    x"348EF6EA",
    x"348EE50C",
    x"348ED330",
    x"348EC157",
    x"348EAF80",
    x"348E9DAB",
    x"348E8BD9",
    x"348E7A08",
    x"348E683A",
    x"348E566E",
    x"348E44A4",
    x"348E32DD",
    x"348E2118",
    x"348E0F55",
    x"348DFD94",
    x"348DEBD5",
    x"348DDA19",
    x"348DC85F",
    x"348DB6A7",
    x"348DA4F1",
    x"348D933E",
    x"348D818C",
    x"348D6FDD",
    x"348D5E30",
    x"348D4C86",
    x"348D3ADD",
    x"348D2937",
    x"348D1793",
    x"348D05F1",
    x"348CF451",
    x"348CE2B4",
    x"348CD119",
    x"348CBF80",
    x"348CADE9",
    x"348C9C54",
    x"348C8AC2",
    x"348C7932",
    x"348C67A4",
    x"348C5618",
    x"348C448E",
    x"348C3307",
    x"348C2181",
    x"348C0FFE",
    x"348BFE7D",
    x"348BECFF",
    x"348BDB82",
    x"348BCA08",
    x"348BB88F",
    x"348BA719",
    x"348B95A6",
    x"348B8434",
    x"348B72C5",
    x"348B6157",
    x"348B4FEC",
    x"348B3E83",
    x"348B2D1D",
    x"348B1BB8",
    x"348B0A56",
    x"348AF8F6",
    x"348AE798",
    x"348AD63C",
    x"348AC4E2",
    x"348AB38A",
    x"348AA235",
    x"348A90E2",
    x"348A7F91",
    x"348A6E42",
    x"348A5CF5",
    x"348A4BAB",
    x"348A3A62",
    x"348A291C",
    x"348A17D8",
    x"348A0696",
    x"3489F556",
    x"3489E419",
    x"3489D2DD",
    x"3489C1A4",
    x"3489B06D",
    x"34899F38",
    x"34898E05",
    x"34897CD5",
    x"34896BA6",
    x"34895A7A",
    x"3489494F",
    x"34893827",
    x"34892701",
    x"348915DE",
    x"348904BC",
    x"3488F39C",
    x"3488E27F",
    x"3488D164",
    x"3488C04B",
    x"3488AF34",
    x"34889E1F",
    x"34888D0C",
    x"34887BFC",
    x"34886AED",
    x"348859E1",
    x"348848D7",
    x"348837CF",
    x"348826C9",
    x"348815C5",
    x"348804C3",
    x"3487F3C4",
    x"3487E2C6",
    x"3487D1CB",
    x"3487C0D2",
    x"3487AFDB",
    x"34879EE6",
    x"34878DF3",
    x"34877D02",
    x"34876C14",
    x"34875B27",
    x"34874A3D",
    x"34873955",
    x"3487286F",
    x"3487178B",
    x"348706A9",
    x"3486F5C9",
    x"3486E4EB",
    x"3486D410",
    x"3486C336",
    x"3486B25F",
    x"3486A18A",
    x"348690B7",
    x"34867FE6",
    x"34866F17",
    x"34865E4A",
    x"34864D7F",
    x"34863CB6",
    x"34862BF0",
    x"34861B2B",
    x"34860A69",
    x"3485F9A9",
    x"3485E8EB",
    x"3485D82F",
    x"3485C775",
    x"3485B6BD",
    x"3485A607",
    x"34859553",
    x"348584A2",
    x"348573F2",
    x"34856345",
    x"34855299",
    x"348541F0",
    x"34853149",
    x"348520A4",
    x"34851001",
    x"3484FF60",
    x"3484EEC1",
    x"3484DE24",
    x"3484CD89",
    x"3484BCF1",
    x"3484AC5A",
    x"34849BC6",
    x"34848B33",
    x"34847AA3",
    x"34846A14",
    x"34845988",
    x"348448FE",
    x"34843876",
    x"348427F0",
    x"3484176C",
    x"348406EA",
    x"3483F66A",
    x"3483E5EC",
    x"3483D571",
    x"3483C4F7",
    x"3483B480",
    x"3483A40A",
    x"34839397",
    x"34838325",
    x"348372B6",
    x"34836248",
    x"348351DD",
    x"34834174",
    x"3483310D",
    x"348320A8",
    x"34831045",
    x"3482FFE4",
    x"3482EF85",
    x"3482DF28",
    x"3482CECD",
    x"3482BE74",
    x"3482AE1D",
    x"34829DC9",
    x"34828D76",
    x"34827D25",
    x"34826CD7",
    x"34825C8A",
    x"34824C3F",
    x"34823BF7",
    x"34822BB0",
    x"34821B6C",
    x"34820B2A",
    x"3481FAE9",
    x"3481EAAB",
    x"3481DA6E",
    x"3481CA34",
    x"3481B9FC",
    x"3481A9C6",
    x"34819991",
    x"3481895F",
    x"3481792F",
    x"34816901",
    x"348158D5",
    x"348148AB",
    x"34813883",
    x"3481285D",
    x"34811839",
    x"34810817",
    x"3480F7F7",
    x"3480E7D9",
    x"3480D7BD",
    x"3480C7A3",
    x"3480B78B",
    x"3480A775",
    x"34809761",
    x"3480874F",
    x"3480773F",
    x"34806731",
    x"34805725",
    x"3480471B",
    x"34803713",
    x"3480270E",
    x"3480170A",
    x"34800708",
    x"347FEE10",
    x"347FCE14",
    x"347FAE1C",
    x"347F8E29",
    x"347F6E39",
    x"347F4E4D",
    x"347F2E65",
    x"347F0E81",
    x"347EEEA2",
    x"347ECEC6",
    x"347EAEEE",
    x"347E8F1A",
    x"347E6F4A",
    x"347E4F7E",
    x"347E2FB6",
    x"347E0FF2",
    x"347DF032",
    x"347DD076",
    x"347DB0BE",
    x"347D910A",
    x"347D715A",
    x"347D51AE",
    x"347D3206",
    x"347D1261",
    x"347CF2C1",
    x"347CD325",
    x"347CB38C",
    x"347C93F8",
    x"347C7467",
    x"347C54DB",
    x"347C3552",
    x"347C15CD",
    x"347BF64C",
    x"347BD6D0",
    x"347BB757",
    x"347B97E2",
    x"347B7871",
    x"347B5904",
    x"347B399B",
    x"347B1A35",
    x"347AFAD4",
    x"347ADB77",
    x"347ABC1D",
    x"347A9CC8",
    x"347A7D76",
    x"347A5E28",
    x"347A3EDE",
    x"347A1F99",
    x"347A0057",
    x"3479E118",
    x"3479C1DE",
    x"3479A2A8",
    x"34798376",
    x"34796447",
    x"3479451D",
    x"347925F6",
    x"347906D3",
    x"3478E7B4",
    x"3478C899",
    x"3478A982",
    x"34788A6F",
    x"34786B5F",
    x"34784C54",
    x"34782D4C",
    x"34780E49",
    x"3477EF49",
    x"3477D04D",
    x"3477B155",
    x"34779260",
    x"34777370",
    x"34775484",
    x"3477359B",
    x"347716B6",
    x"3476F7D5",
    x"3476D8F8",
    x"3476BA1F",
    x"34769B4A",
    x"34767C78",
    x"34765DAB",
    x"34763EE1",
    x"3476201B",
    x"34760159",
    x"3475E29A",
    x"3475C3E0",
    x"3475A529",
    x"34758677",
    x"347567C8",
    x"3475491D",
    x"34752A76",
    x"34750BD2",
    x"3474ED33",
    x"3474CE97",
    x"3474AFFF",
    x"3474916B",
    x"347472DB",
    x"3474544E",
    x"347435C6",
    x"34741741",
    x"3473F8C0",
    x"3473DA43",
    x"3473BBC9",
    x"34739D54",
    x"34737EE2",
    x"34736074",
    x"3473420A",
    x"347323A3",
    x"34730541",
    x"3472E6E2",
    x"3472C887",
    x"3472AA30",
    x"34728BDD",
    x"34726D8D",
    x"34724F41",
    x"347230F9",
    x"347212B5",
    x"3471F474",
    x"3471D638",
    x"3471B7FF",
    x"347199CA",
    x"34717B98",
    x"34715D6B",
    x"34713F41",
    x"3471211B",
    x"347102F9",
    x"3470E4DA",
    x"3470C6C0",
    x"3470A8A9",
    x"34708A95",
    x"34706C86",
    x"34704E7A",
    x"34703072",
    x"3470126E",
    x"346FF46E",
    x"346FD671",
    x"346FB878",
    x"346F9A83",
    x"346F7C92",
    x"346F5EA4",
    x"346F40BA",
    x"346F22D4",
    x"346F04F1",
    x"346EE712",
    x"346EC937",
    x"346EAB60",
    x"346E8D8D",
    x"346E6FBD",
    x"346E51F1",
    x"346E3428",
    x"346E1664",
    x"346DF8A3",
    x"346DDAE5",
    x"346DBD2C",
    x"346D9F76",
    x"346D81C4",
    x"346D6416",
    x"346D466B",
    x"346D28C4",
    x"346D0B21",
    x"346CED81",
    x"346CCFE5",
    x"346CB24D",
    x"346C94B9",
    x"346C7728",
    x"346C599B",
    x"346C3C12",
    x"346C1E8C",
    x"346C010A",
    x"346BE38C",
    x"346BC611",
    x"346BA89A",
    x"346B8B27",
    x"346B6DB8",
    x"346B504C",
    x"346B32E3",
    x"346B157F",
    x"346AF81E",
    x"346ADAC1",
    x"346ABD67",
    x"346AA012",
    x"346A82BF",
    x"346A6571",
    x"346A4826",
    x"346A2ADF",
    x"346A0D9B",
    x"3469F05B",
    x"3469D31F",
    x"3469B5E7",
    x"346998B2",
    x"34697B80",
    x"34695E53",
    x"34694129",
    x"34692403",
    x"346906E0",
    x"3468E9C1",
    x"3468CCA5",
    x"3468AF8E",
    x"3468927A",
    x"34687569",
    x"3468585C",
    x"34683B53",
    x"34681E4D",
    x"3468014B",
    x"3467E44D",
    x"3467C752",
    x"3467AA5B",
    x"34678D68",
    x"34677078",
    x"3467538C",
    x"346736A3",
    x"346719BE",
    x"3466FCDD",
    x"3466DFFF",
    x"3466C325",
    x"3466A64E",
    x"3466897B",
    x"34666CAC",
    x"34664FE0",
    x"34663318",
    x"34661653",
    x"3465F992",
    x"3465DCD5",
    x"3465C01B",
    x"3465A365",
    x"346586B2",
    x"34656A03",
    x"34654D57",
    x"346530B0",
    x"3465140B",
    x"3464F76B",
    x"3464DACD",
    x"3464BE34",
    x"3464A19E",
    x"3464850B",
    x"3464687D",
    x"34644BF1",
    x"34642F6A",
    x"346412E5",
    x"3463F665",
    x"3463D9E8",
    x"3463BD6E",
    x"3463A0F9",
    x"34638486",
    x"34636817",
    x"34634BAC",
    x"34632F44",
    x"346312E0",
    x"3462F680",
    x"3462DA23",
    x"3462BDC9",
    x"3462A173",
    x"34628521",
    x"346268D2",
    x"34624C87",
    x"3462303F",
    x"346213FB",
    x"3461F7BA",
    x"3461DB7D",
    x"3461BF43",
    x"3461A30D",
    x"346186DA",
    x"34616AAB",
    x"34614E80",
    x"34613258",
    x"34611633",
    x"3460FA12",
    x"3460DDF4",
    x"3460C1DA",
    x"3460A5C4",
    x"346089B1",
    x"34606DA2",
    x"34605196",
    x"3460358D",
    x"34601988",
    x"345FFD87",
    x"345FE189",
    x"345FC58E",
    x"345FA997",
    x"345F8DA4",
    x"345F71B4",
    x"345F55C8",
    x"345F39DF",
    x"345F1DF9",
    x"345F0217",
    x"345EE639",
    x"345ECA5E",
    x"345EAE86",
    x"345E92B2",
    x"345E76E1",
    x"345E5B14",
    x"345E3F4B",
    x"345E2384",
    x"345E07C2",
    x"345DEC02",
    x"345DD047",
    x"345DB48E",
    x"345D98DA",
    x"345D7D28",
    x"345D617A",
    x"345D45D0",
    x"345D2A29",
    x"345D0E85",
    x"345CF2E5",
    x"345CD749",
    x"345CBBAF",
    x"345CA01A",
    x"345C8487",
    x"345C68F8",
    x"345C4D6D",
    x"345C31E5",
    x"345C1661",
    x"345BFAE0",
    x"345BDF62",
    x"345BC3E8",
    x"345BA871",
    x"345B8CFE",
    x"345B718E",
    x"345B5621",
    x"345B3AB8",
    x"345B1F52",
    x"345B03F0",
    x"345AE892",
    x"345ACD36",
    x"345AB1DE",
    x"345A968A",
    x"345A7B39",
    x"345A5FEB",
    x"345A44A1",
    x"345A295A",
    x"345A0E16",
    x"3459F2D6",
    x"3459D79A",
    x"3459BC60",
    x"3459A12A",
    x"345985F8",
    x"34596AC9",
    x"34594F9D",
    x"34593475",
    x"34591950",
    x"3458FE2F",
    x"3458E311",
    x"3458C7F6",
    x"3458ACDF",
    x"345891CB",
    x"345876BA",
    x"34585BAD",
    x"345840A3",
    x"3458259D",
    x"34580A9A",
    x"3457EF9A",
    x"3457D49E",
    x"3457B9A5",
    x"34579EB0",
    x"345783BD",
    x"345768CF",
    x"34574DE3",
    x"345732FB",
    x"34571816",
    x"3456FD35",
    x"3456E257",
    x"3456C77D",
    x"3456ACA5",
    x"345691D1",
    x"34567701",
    x"34565C34",
    x"3456416A",
    x"345626A3",
    x"34560BE0",
    x"3455F120",
    x"3455D664",
    x"3455BBAB",
    x"3455A0F5",
    x"34558642",
    x"34556B93",
    x"345550E8",
    x"3455363F",
    x"34551B9A",
    x"345500F8",
    x"3454E65A",
    x"3454CBBF",
    x"3454B127",
    x"34549692",
    x"34547C01",
    x"34546173",
    x"345446E9",
    x"34542C62",
    x"345411DE",
    x"3453F75D",
    x"3453DCE0",
    x"3453C266",
    x"3453A7EF",
    x"34538D7C",
    x"3453730C",
    x"3453589F",
    x"34533E36",
    x"345323D0",
    x"3453096D",
    x"3452EF0D",
    x"3452D4B1",
    x"3452BA58",
    x"3452A002",
    x"345285B0",
    x"34526B61",
    x"34525115",
    x"345236CD",
    x"34521C88",
    x"34520246",
    x"3451E807",
    x"3451CDCC",
    x"3451B394",
    x"3451995F",
    x"34517F2D",
    x"345164FF",
    x"34514AD4",
    x"345130AC",
    x"34511688",
    x"3450FC67",
    x"3450E249",
    x"3450C82E",
    x"3450AE17",
    x"34509403",
    x"345079F2",
    x"34505FE4",
    x"345045DA",
    x"34502BD3",
    x"345011CF",
    x"344FF7CE",
    x"344FDDD1",
    x"344FC3D7",
    x"344FA9E0",
    x"344F8FEC",
    x"344F75FC",
    x"344F5C0F",
    x"344F4225",
    x"344F283E",
    x"344F0E5B",
    x"344EF47B",
    x"344EDA9E",
    x"344EC0C4",
    x"344EA6ED",
    x"344E8D1A",
    x"344E734A",
    x"344E597D",
    x"344E3FB4",
    x"344E25ED",
    x"344E0C2A",
    x"344DF26A",
    x"344DD8AE",
    x"344DBEF4",
    x"344DA53E",
    x"344D8B8B",
    x"344D71DB",
    x"344D582E",
    x"344D3E85",
    x"344D24DF",
    x"344D0B3C",
    x"344CF19C",
    x"344CD7FF",
    x"344CBE66",
    x"344CA4D0",
    x"344C8B3D",
    x"344C71AD",
    x"344C5820",
    x"344C3E97",
    x"344C2511",
    x"344C0B8E",
    x"344BF20E",
    x"344BD891",
    x"344BBF18",
    x"344BA5A1",
    x"344B8C2E",
    x"344B72BE",
    x"344B5952",
    x"344B3FE8",
    x"344B2682",
    x"344B0D1E",
    x"344AF3BE",
    x"344ADA61",
    x"344AC108",
    x"344AA7B1",
    x"344A8E5E",
    x"344A750E",
    x"344A5BC1",
    x"344A4277",
    x"344A2930",
    x"344A0FEC",
    x"3449F6AC",
    x"3449DD6F",
    x"3449C435",
    x"3449AAFE",
    x"344991CA",
    x"34497899",
    x"34495F6C",
    x"34494641",
    x"34492D1A",
    x"344913F6",
    x"3448FAD5",
    x"3448E1B7",
    x"3448C89D",
    x"3448AF85",
    x"34489671",
    x"34487D60",
    x"34486451",
    x"34484B47",
    x"3448323F",
    x"3448193A",
    x"34480038",
    x"3447E73A",
    x"3447CE3F",
    x"3447B546",
    x"34479C51",
    x"3447835F",
    x"34476A70",
    x"34475185",
    x"3447389C",
    x"34471FB6",
    x"344706D4",
    x"3446EDF5",
    x"3446D519",
    x"3446BC40",
    x"3446A36A",
    x"34468A97",
    x"344671C7",
    x"344658FA",
    x"34464031",
    x"3446276A",
    x"34460EA7",
    x"3445F5E7",
    x"3445DD29",
    x"3445C46F",
    x"3445ABB8",
    x"34459304",
    x"34457A53",
    x"344561A6",
    x"344548FB",
    x"34453053",
    x"344517AF",
    x"3444FF0E",
    x"3444E66F",
    x"3444CDD4",
    x"3444B53C",
    x"34449CA7",
    x"34448415",
    x"34446B86",
    x"344452FA",
    x"34443A71",
    x"344421EB",
    x"34440968",
    x"3443F0E9",
    x"3443D86C",
    x"3443BFF3",
    x"3443A77C",
    x"34438F09",
    x"34437698",
    x"34435E2B",
    x"344345C1",
    x"34432D5A",
    x"344314F6",
    x"3442FC94",
    x"3442E436",
    x"3442CBDB",
    x"3442B383",
    x"34429B2E",
    x"344282DD",
    x"34426A8E",
    x"34425242",
    x"344239F9",
    x"344221B3",
    x"34420971",
    x"3441F131",
    x"3441D8F4",
    x"3441C0BB",
    x"3441A884",
    x"34419051",
    x"34417820",
    x"34415FF3",
    x"344147C8",
    x"34412FA1",
    x"3441177C",
    x"3440FF5B",
    x"3440E73C",
    x"3440CF21",
    x"3440B709",
    x"34409EF3",
    x"344086E1",
    x"34406ED2",
    x"344056C5",
    x"34403EBC",
    x"344026B6",
    x"34400EB2",
    x"343FF6B2",
    x"343FDEB5",
    x"343FC6BA",
    x"343FAEC3",
    x"343F96CF",
    x"343F7EDD",
    x"343F66EF",
    x"343F4F03",
    x"343F371B",
    x"343F1F36",
    x"343F0753",
    x"343EEF74",
    x"343ED797",
    x"343EBFBE",
    x"343EA7E7",
    x"343E9014",
    x"343E7843",
    x"343E6076",
    x"343E48AB",
    x"343E30E4",
    x"343E191F",
    x"343E015D",
    x"343DE99F",
    x"343DD1E3",
    x"343DBA2A",
    x"343DA274",
    x"343D8AC2",
    x"343D7312",
    x"343D5B65",
    x"343D43BB",
    x"343D2C14",
    x"343D1470",
    x"343CFCCF",
    x"343CE531",
    x"343CCD96",
    x"343CB5FD",
    x"343C9E68",
    x"343C86D6",
    x"343C6F46",
    x"343C57BA",
    x"343C4030",
    x"343C28AA",
    x"343C1126",
    x"343BF9A6",
    x"343BE228",
    x"343BCAAD",
    x"343BB335",
    x"343B9BC0",
    x"343B844E",
    x"343B6CDF",
    x"343B5573",
    x"343B3E0A",
    x"343B26A4",
    x"343B0F40",
    x"343AF7E0",
    x"343AE082",
    x"343AC928",
    x"343AB1D0",
    x"343A9A7B",
    x"343A8329",
    x"343A6BDA",
    x"343A548E",
    x"343A3D45",
    x"343A25FF",
    x"343A0EBC",
    x"3439F77B",
    x"3439E03E",
    x"3439C903",
    x"3439B1CC",
    x"34399A97",
    x"34398365",
    x"34396C36",
    x"3439550A",
    x"34393DE1",
    x"343926BA",
    x"34390F97",
    x"3438F876",
    x"3438E159",
    x"3438CA3E",
    x"3438B326",
    x"34389C11",
    x"343884FF",
    x"34386DF0",
    x"343856E4",
    x"34383FDA",
    x"343828D4",
    x"343811D0",
    x"3437FACF",
    x"3437E3D1",
    x"3437CCD6",
    x"3437B5DE",
    x"34379EE9",
    x"343787F7",
    x"34377107",
    x"34375A1A",
    x"34374330",
    x"34372C49",
    x"34371565",
    x"3436FE84",
    x"3436E7A6",
    x"3436D0CA",
    x"3436B9F2",
    x"3436A31C",
    x"34368C49",
    x"34367579",
    x"34365EAB",
    x"343647E1",
    x"34363119",
    x"34361A55",
    x"34360393",
    x"3435ECD4",
    x"3435D618",
    x"3435BF5E",
    x"3435A8A8",
    x"343591F4",
    x"34357B43",
    x"34356495",
    x"34354DEA",
    x"34353742",
    x"3435209C",
    x"343509FA",
    x"3434F35A",
    x"3434DCBD",
    x"3434C623",
    x"3434AF8B",
    x"343498F7",
    x"34348265",
    x"34346BD6",
    x"3434554A",
    x"34343EC1",
    x"3434283A",
    x"343411B7",
    x"3433FB36",
    x"3433E4B8",
    x"3433CE3D",
    x"3433B7C4",
    x"3433A14F",
    x"34338ADC",
    x"3433746C",
    x"34335DFF",
    x"34334795",
    x"3433312D",
    x"34331AC8",
    x"34330466",
    x"3432EE07",
    x"3432D7AB",
    x"3432C151",
    x"3432AAFB",
    x"343294A7",
    x"34327E55",
    x"34326807",
    x"343251BB",
    x"34323B73",
    x"3432252D",
    x"34320EE9",
    x"3431F8A9",
    x"3431E26B",
    x"3431CC30",
    x"3431B5F8",
    x"34319FC3",
    x"34318990",
    x"34317360",
    x"34315D33",
    x"34314709",
    x"343130E2",
    x"34311ABD",
    x"3431049B",
    x"3430EE7C",
    x"3430D85F",
    x"3430C246",
    x"3430AC2F",
    x"3430961B",
    x"34308009",
    x"343069FB",
    x"343053EF",
    x"34303DE6",
    x"343027DF",
    x"343011DC",
    x"342FFBDB",
    x"342FE5DD",
    x"342FCFE1",
    x"342FB9E9",
    x"342FA3F3",
    x"342F8E00",
    x"342F780F",
    x"342F6222",
    x"342F4C37",
    x"342F364F",
    x"342F2069",
    x"342F0A86",
    x"342EF4A7",
    x"342EDEC9",
    x"342EC8EF",
    x"342EB317",
    x"342E9D42",
    x"342E8770",
    x"342E71A0",
    x"342E5BD3",
    x"342E4609",
    x"342E3042",
    x"342E1A7D",
    x"342E04BB",
    x"342DEEFC",
    x"342DD93F",
    x"342DC386",
    x"342DADCF",
    x"342D981A",
    x"342D8269",
    x"342D6CBA",
    x"342D570D",
    x"342D4164",
    x"342D2BBD",
    x"342D1619",
    x"342D0078",
    x"342CEAD9",
    x"342CD53D",
    x"342CBFA3",
    x"342CAA0D",
    x"342C9479",
    x"342C7EE8",
    x"342C6959",
    x"342C53CD",
    x"342C3E44",
    x"342C28BE",
    x"342C133A",
    x"342BFDB9",
    x"342BE83B",
    x"342BD2BF",
    x"342BBD46",
    x"342BA7D0",
    x"342B925C",
    x"342B7CEB",
    x"342B677D",
    x"342B5211",
    x"342B3CA8",
    x"342B2742",
    x"342B11DE",
    x"342AFC7E",
    x"342AE71F",
    x"342AD1C4",
    x"342ABC6B",
    x"342AA715",
    x"342A91C1",
    x"342A7C70",
    x"342A6722",
    x"342A51D6",
    x"342A3C8E",
    x"342A2747",
    x"342A1204",
    x"3429FCC3",
    x"3429E785",
    x"3429D249",
    x"3429BD10",
    x"3429A7DA",
    x"342992A6",
    x"34297D75",
    x"34296847",
    x"3429531B",
    x"34293DF2",
    x"342928CB",
    x"342913A8",
    x"3428FE87",
    x"3428E968",
    x"3428D44C",
    x"3428BF33",
    x"3428AA1C",
    x"34289508",
    x"34287FF7",
    x"34286AE8",
    x"342855DC",
    x"342840D3",
    x"34282BCC",
    x"342816C8",
    x"342801C7",
    x"3427ECC8",
    x"3427D7CB",
    x"3427C2D2",
    x"3427ADDB",
    x"342798E6",
    x"342783F4",
    x"34276F05",
    x"34275A19",
    x"3427452F",
    x"34273047",
    x"34271B63",
    x"34270680",
    x"3426F1A1",
    x"3426DCC4",
    x"3426C7EA",
    x"3426B312",
    x"34269E3D",
    x"3426896B",
    x"3426749B",
    x"34265FCD",
    x"34264B03",
    x"3426363B",
    x"34262175",
    x"34260CB2",
    x"3425F7F2",
    x"3425E334",
    x"3425CE79",
    x"3425B9C1",
    x"3425A50B",
    x"34259057",
    x"34257BA7",
    x"342566F8",
    x"3425524D",
    x"34253DA4",
    x"342528FE",
    x"3425145A",
    x"3424FFB8",
    x"3424EB1A",
    x"3424D67E",
    x"3424C1E4",
    x"3424AD4D",
    x"342498B9",
    x"34248427",
    x"34246F98",
    x"34245B0B",
    x"34244681",
    x"342431F9",
    x"34241D75",
    x"342408F2",
    x"3423F472",
    x"3423DFF5",
    x"3423CB7A",
    x"3423B702",
    x"3423A28D",
    x"34238E19",
    x"342379A9",
    x"3423653B",
    x"342350D0",
    x"34233C67",
    x"34232801",
    x"3423139D",
    x"3422FF3C",
    x"3422EADD",
    x"3422D681",
    x"3422C227",
    x"3422ADD0",
    x"3422997C",
    x"3422852A",
    x"342270DB",
    x"34225C8E",
    x"34224844",
    x"342233FC",
    x"34221FB7",
    x"34220B74",
    x"3421F734",
    x"3421E2F6",
    x"3421CEBB",
    x"3421BA82",
    x"3421A64C",
    x"34219219",
    x"34217DE8",
    x"342169B9",
    x"3421558D",
    x"34214164",
    x"34212D3D",
    x"34211919",
    x"342104F7",
    x"3420F0D7",
    x"3420DCBB",
    x"3420C8A0",
    x"3420B488",
    x"3420A073",
    x"34208C60",
    x"34207850",
    x"34206442",
    x"34205037",
    x"34203C2E",
    x"34202828",
    x"34201424",
    x"34200023",
    x"341FEC24",
    x"341FD828",
    x"341FC42E",
    x"341FB037",
    x"341F9C42",
    x"341F8850",
    x"341F7460",
    x"341F6073",
    x"341F4C88",
    x"341F389F",
    x"341F24BA",
    x"341F10D6",
    x"341EFCF5",
    x"341EE917",
    x"341ED53B",
    x"341EC162",
    x"341EAD8B",
    x"341E99B6",
    x"341E85E4",
    x"341E7215",
    x"341E5E48",
    x"341E4A7D",
    x"341E36B5",
    x"341E22F0",
    x"341E0F2C",
    x"341DFB6C",
    x"341DE7AE",
    x"341DD3F2",
    x"341DC039",
    x"341DAC82",
    x"341D98CE",
    x"341D851C",
    x"341D716C",
    x"341D5DBF",
    x"341D4A15",
    x"341D366D",
    x"341D22C7",
    x"341D0F24",
    x"341CFB83",
    x"341CE7E5",
    x"341CD449",
    x"341CC0B0",
    x"341CAD19",
    x"341C9985",
    x"341C85F3",
    x"341C7263",
    x"341C5ED6",
    x"341C4B4C",
    x"341C37C3",
    x"341C243E",
    x"341C10BA",
    x"341BFD3A",
    x"341BE9BB",
    x"341BD63F",
    x"341BC2C6",
    x"341BAF4E",
    x"341B9BDA",
    x"341B8867",
    x"341B74F8",
    x"341B618A",
    x"341B4E1F",
    x"341B3AB7",
    x"341B2751",
    x"341B13ED",
    x"341B008C",
    x"341AED2D",
    x"341AD9D0",
    x"341AC676",
    x"341AB31F",
    x"341A9FC9",
    x"341A8C77",
    x"341A7926",
    x"341A65D8",
    x"341A528D",
    x"341A3F44",
    x"341A2BFD",
    x"341A18B9",
    x"341A0577",
    x"3419F237",
    x"3419DEFA",
    x"3419CBC0",
    x"3419B887",
    x"3419A552",
    x"3419921E",
    x"34197EED",
    x"34196BBE",
    x"34195892",
    x"34194568",
    x"34193241",
    x"34191F1C",
    x"34190BF9",
    x"3418F8D9",
    x"3418E5BB",
    x"3418D29F",
    x"3418BF86",
    x"3418AC6F",
    x"3418995B",
    x"34188649",
    x"34187339",
    x"3418602C",
    x"34184D21",
    x"34183A19",
    x"34182713",
    x"3418140F",
    x"3418010E",
    x"3417EE0F",
    x"3417DB12",
    x"3417C818",
    x"3417B520",
    x"3417A22B",
    x"34178F38",
    x"34177C47",
    x"34176959",
    x"3417566D",
    x"34174383",
    x"3417309C",
    x"34171DB7",
    x"34170AD4",
    x"3416F7F4",
    x"3416E516",
    x"3416D23B",
    x"3416BF62",
    x"3416AC8B",
    x"341699B7",
    x"341686E5",
    x"34167415",
    x"34166148",
    x"34164E7D",
    x"34163BB4",
    x"341628EE",
    x"3416162A",
    x"34160368",
    x"3415F0A9",
    x"3415DDEC",
    x"3415CB31",
    x"3415B879",
    x"3415A5C3",
    x"34159310",
    x"3415805F",
    x"34156DB0",
    x"34155B03",
    x"34154859",
    x"341535B1",
    x"3415230B",
    x"34151068",
    x"3414FDC7",
    x"3414EB29",
    x"3414D88D",
    x"3414C5F3",
    x"3414B35B",
    x"3414A0C6",
    x"34148E33",
    x"34147BA2",
    x"34146914",
    x"34145688",
    x"341443FE",
    x"34143177",
    x"34141EF2",
    x"34140C6F",
    x"3413F9EF",
    x"3413E771",
    x"3413D4F5",
    x"3413C27C",
    x"3413B004",
    x"34139D90",
    x"34138B1D",
    x"341378AD",
    x"3413663F",
    x"341353D3",
    x"3413416A",
    x"34132F03",
    x"34131C9E",
    x"34130A3C",
    x"3412F7DC",
    x"3412E57E",
    x"3412D322",
    x"3412C0C9",
    x"3412AE72",
    x"34129C1D",
    x"341289CB",
    x"3412777B",
    x"3412652D",
    x"341252E2",
    x"34124098",
    x"34122E51",
    x"34121C0D",
    x"341209CA",
    x"3411F78A",
    x"3411E54D",
    x"3411D311",
    x"3411C0D8",
    x"3411AEA1",
    x"34119C6C",
    x"34118A3A",
    x"3411780A",
    x"341165DC",
    x"341153B0",
    x"34114187",
    x"34112F60",
    x"34111D3B",
    x"34110B18",
    x"3410F8F8",
    x"3410E6DA",
    x"3410D4BE",
    x"3410C2A5",
    x"3410B08E",
    x"34109E79",
    x"34108C66",
    x"34107A56",
    x"34106848",
    x"3410563C",
    x"34104432",
    x"3410322B",
    x"34102025",
    x"34100E23",
    x"340FFC22",
    x"340FEA24",
    x"340FD827",
    x"340FC62E",
    x"340FB436",
    x"340FA240",
    x"340F904D",
    x"340F7E5C",
    x"340F6C6E",
    x"340F5A81",
    x"340F4897",
    x"340F36AF",
    x"340F24C9",
    x"340F12E6",
    x"340F0105",
    x"340EEF26",
    x"340EDD49",
    x"340ECB6E",
    x"340EB996",
    x"340EA7C0",
    x"340E95EC",
    x"340E841A",
    x"340E724B",
    x"340E607E",
    x"340E4EB3",
    x"340E3CEA",
    x"340E2B24",
    x"340E195F",
    x"340E079D",
    x"340DF5DE",
    x"340DE420",
    x"340DD265",
    x"340DC0AB",
    x"340DAEF4",
    x"340D9D40",
    x"340D8B8D",
    x"340D79DD",
    x"340D682F",
    x"340D5683",
    x"340D44D9",
    x"340D3331",
    x"340D218C",
    x"340D0FE9",
    x"340CFE48",
    x"340CECA9",
    x"340CDB0D",
    x"340CC973",
    x"340CB7DB",
    x"340CA645",
    x"340C94B1",
    x"340C8320",
    x"340C7190",
    x"340C6003",
    x"340C4E78",
    x"340C3CF0",
    x"340C2B69",
    x"340C19E5",
    x"340C0863",
    x"340BF6E3",
    x"340BE565",
    x"340BD3E9",
    x"340BC270",
    x"340BB0F9",
    x"340B9F84",
    x"340B8E11",
    x"340B7CA0",
    x"340B6B32",
    x"340B59C5",
    x"340B485B",
    x"340B36F3",
    x"340B258D",
    x"340B142A",
    x"340B02C8",
    x"340AF169",
    x"340AE00C",
    x"340ACEB1",
    x"340ABD58",
    x"340AAC02",
    x"340A9AAD",
    x"340A895B",
    x"340A780B",
    x"340A66BD",
    x"340A5571",
    x"340A4428",
    x"340A32E0",
    x"340A219B",
    x"340A1058",
    x"3409FF17",
    x"3409EDD8",
    x"3409DC9B",
    x"3409CB61",
    x"3409BA29",
    x"3409A8F2",
    x"340997BE",
    x"3409868D",
    x"3409755D",
    x"3409642F",
    x"34095304",
    x"340941DA",
    x"340930B3",
    x"34091F8E",
    x"34090E6B",
    x"3408FD4B",
    x"3408EC2C",
    x"3408DB10",
    x"3408C9F5",
    x"3408B8DD",
    x"3408A7C7",
    x"340896B3",
    x"340885A1",
    x"34087492",
    x"34086384",
    x"34085279",
    x"34084170",
    x"34083069",
    x"34081F64",
    x"34080E61",
    x"3407FD60",
    x"3407EC61",
    x"3407DB65",
    x"3407CA6A",
    x"3407B972",
    x"3407A87C",
    x"34079788",
    x"34078696",
    x"340775A6",
    x"340764B9",
    x"340753CD",
    x"340742E4",
    x"340731FD",
    x"34072117",
    x"34071034",
    x"3406FF53",
    x"3406EE74",
    x"3406DD98",
    x"3406CCBD",
    x"3406BBE5",
    x"3406AB0E",
    x"34069A3A",
    x"34068968",
    x"34067897",
    x"340667C9",
    x"340656FD",
    x"34064634",
    x"3406356C",
    x"340624A6",
    x"340613E3",
    x"34060321",
    x"3405F262",
    x"3405E1A5",
    x"3405D0EA",
    x"3405C030",
    x"3405AF7A",
    x"34059EC5",
    x"34058E12",
    x"34057D61",
    x"34056CB2",
    x"34055C06",
    x"34054B5B",
    x"34053AB3",
    x"34052A0D",
    x"34051969",
    x"340508C6",
    x"3404F826",
    x"3404E788",
    x"3404D6EC",
    x"3404C653",
    x"3404B5BB",
    x"3404A525",
    x"34049492",
    x"34048400",
    x"34047371",
    x"340462E3",
    x"34045258",
    x"340441CF",
    x"34043147",
    x"340420C2",
    x"3404103F",
    x"3403FFBE",
    x"3403EF3F",
    x"3403DEC2",
    x"3403CE48",
    x"3403BDCF",
    x"3403AD58",
    x"34039CE4",
    x"34038C71",
    x"34037C00",
    x"34036B92",
    x"34035B26",
    x"34034ABB",
    x"34033A53",
    x"340329ED",
    x"34031988",
    x"34030926",
    x"3402F8C6",
    x"3402E868",
    x"3402D80C",
    x"3402C7B2",
    x"3402B75A",
    x"3402A704",
    x"340296B0",
    x"3402865E",
    x"3402760F",
    x"340265C1",
    x"34025575",
    x"3402452C",
    x"340234E4",
    x"3402249E",
    x"3402145B",
    x"34020419",
    x"3401F3DA",
    x"3401E39C",
    x"3401D361",
    x"3401C327",
    x"3401B2F0",
    x"3401A2BB",
    x"34019287",
    x"34018256",
    x"34017227",
    x"340161FA",
    x"340151CE",
    x"340141A5",
    x"3401317E",
    x"34012159",
    x"34011136",
    x"34010114",
    x"3400F0F5",
    x"3400E0D8",
    x"3400D0BD",
    x"3400C0A4",
    x"3400B08D",
    x"3400A078",
    x"34009065",
    x"34008054",
    x"34007045",
    x"34006038",
    x"3400502D",
    x"34004024",
    x"3400301D",
    x"34002018",
    x"34001015",
    x"34000014",
    x"33FFE029",
    x"33FFC02F",
    x"33FFA039",
    x"33FF8047",
    x"33FF6059",
    x"33FF406F",
    x"33FF2089",
    x"33FF00A7",
    x"33FEE0C9",
    x"33FEC0EF",
    x"33FEA119",
    x"33FE8146",
    x"33FE6178",
    x"33FE41AE",
    x"33FE21E8",
    x"33FE0226",
    x"33FDE267",
    x"33FDC2AD",
    x"33FDA2F7",
    x"33FD8344",
    x"33FD6396",
    x"33FD43EB",
    x"33FD2445",
    x"33FD04A2",
    x"33FCE504",
    x"33FCC569",
    x"33FCA5D2",
    x"33FC8640",
    x"33FC66B1",
    x"33FC4726",
    x"33FC279F",
    x"33FC081C",
    x"33FBE89D",
    x"33FBC922",
    x"33FBA9AB",
    x"33FB8A37",
    x"33FB6AC8",
    x"33FB4B5D",
    x"33FB2BF5",
    x"33FB0C92",
    x"33FAED32",
    x"33FACDD6",
    x"33FAAE7F",
    x"33FA8F2B",
    x"33FA6FDB",
    x"33FA508F",
    x"33FA3147",
    x"33FA1203",
    x"33F9F2C2",
    x"33F9D386",
    x"33F9B44D",
    x"33F99519",
    x"33F975E8",
    x"33F956BB",
    x"33F93792",
    x"33F9186D",
    x"33F8F94C",
    x"33F8DA2F",
    x"33F8BB16",
    x"33F89C00",
    x"33F87CEF",
    x"33F85DE1",
    x"33F83ED7",
    x"33F81FD1",
    x"33F800CF",
    x"33F7E1D1",
    x"33F7C2D7",
    x"33F7A3E0",
    x"33F784EE",
    x"33F765FF",
    x"33F74714",
    x"33F7282D",
    x"33F7094A",
    x"33F6EA6B",
    x"33F6CB90",
    x"33F6ACB8",
    x"33F68DE5",
    x"33F66F15",
    x"33F65049",
    x"33F63181",
    x"33F612BC",
    x"33F5F3FC",
    x"33F5D53F",
    x"33F5B687",
    x"33F597D2",
    x"33F57921",
    x"33F55A74",
    x"33F53BCA",
    x"33F51D25",
    x"33F4FE83",
    x"33F4DFE5",
    x"33F4C14B",
    x"33F4A2B5",
    x"33F48422",
    x"33F46594",
    x"33F44709",
    x"33F42882",
    x"33F409FF",
    x"33F3EB7F",
    x"33F3CD04",
    x"33F3AE8C",
    x"33F39018",
    x"33F371A8",
    x"33F3533C",
    x"33F334D3",
    x"33F3166F",
    x"33F2F80E",
    x"33F2D9B1",
    x"33F2BB57",
    x"33F29D02",
    x"33F27EB0",
    x"33F26062",
    x"33F24218",
    x"33F223D2",
    x"33F2058F",
    x"33F1E750",
    x"33F1C915",
    x"33F1AADE",
    x"33F18CAA",
    x"33F16E7B",
    x"33F1504F",
    x"33F13227",
    x"33F11402",
    x"33F0F5E2",
    x"33F0D7C5",
    x"33F0B9AC",
    x"33F09B96",
    x"33F07D85",
    x"33F05F77",
    x"33F0416D",
    x"33F02367",
    x"33F00564",
    x"33EFE765",
    x"33EFC96A",
    x"33EFAB73",
    x"33EF8D7F",
    x"33EF6F90",
    x"33EF51A3",
    x"33EF33BB",
    x"33EF15D7",
    x"33EEF7F6",
    x"33EEDA19",
    x"33EEBC3F",
    x"33EE9E69",
    x"33EE8098",
    x"33EE62C9",
    x"33EE44FF",
    x"33EE2738",
    x"33EE0975",
    x"33EDEBB6",
    x"33EDCDFA",
    x"33EDB042",
    x"33ED928E",
    x"33ED74DE",
    x"33ED5731",
    x"33ED3988",
    x"33ED1BE2",
    x"33ECFE41",
    x"33ECE0A3",
    x"33ECC309",
    x"33ECA572",
    x"33EC87DF",
    x"33EC6A50",
    x"33EC4CC5",
    x"33EC2F3D",
    x"33EC11B9",
    x"33EBF438",
    x"33EBD6BC",
    x"33EBB943",
    x"33EB9BCD",
    x"33EB7E5C",
    x"33EB60EE",
    x"33EB4384",
    x"33EB261D",
    x"33EB08BA",
    x"33EAEB5B",
    x"33EACDFF",
    x"33EAB0A7",
    x"33EA9353",
    x"33EA7603",
    x"33EA58B6",
    x"33EA3B6C",
    x"33EA1E27",
    x"33EA00E5",
    x"33E9E3A7",
    x"33E9C66C",
    x"33E9A935",
    x"33E98C02",
    x"33E96ED2",
    x"33E951A6",
    x"33E9347D",
    x"33E91759",
    x"33E8FA38",
    x"33E8DD1A",
    x"33E8C000",
    x"33E8A2EA",
    x"33E885D8",
    x"33E868C9",
    x"33E84BBD",
    x"33E82EB6",
    x"33E811B2",
    x"33E7F4B1",
    x"33E7D7B5",
    x"33E7BABB",
    x"33E79DC6",
    x"33E780D4",
    x"33E763E6",
    x"33E746FB",
    x"33E72A14",
    x"33E70D31",
    x"33E6F051",
    x"33E6D374",
    x"33E6B69C",
    x"33E699C7",
    x"33E67CF5",
    x"33E66028",
    x"33E6435D",
    x"33E62697",
    x"33E609D4",
    x"33E5ED14",
    x"33E5D058",
    x"33E5B3A0",
    x"33E596EB",
    x"33E57A3A",
    x"33E55D8D",
    x"33E540E3",
    x"33E5243D",
    x"33E5079A",
    x"33E4EAFB",
    x"33E4CE5F",
    x"33E4B1C7",
    x"33E49533",
    x"33E478A2",
    x"33E45C15",
    x"33E43F8B",
    x"33E42305",
    x"33E40682",
    x"33E3EA03",
    x"33E3CD88",
    x"33E3B110",
    x"33E3949B",
    x"33E3782B",
    x"33E35BBD",
    x"33E33F54",
    x"33E322ED",
    x"33E3068B",
    x"33E2EA2C",
    x"33E2CDD0",
    x"33E2B178",
    x"33E29524",
    x"33E278D3",
    x"33E25C86",
    x"33E2403C",
    x"33E223F6",
    x"33E207B3",
    x"33E1EB74",
    x"33E1CF38",
    x"33E1B300",
    x"33E196CB",
    x"33E17A9A",
    x"33E15E6D",
    x"33E14243",
    x"33E1261C",
    x"33E109F9",
    x"33E0EDDA",
    x"33E0D1BE",
    x"33E0B5A5",
    x"33E09990",
    x"33E07D7F",
    x"33E06171",
    x"33E04566",
    x"33E02960",
    x"33E00D5C",
    x"33DFF15C",
    x"33DFD560",
    x"33DFB967",
    x"33DF9D71",
    x"33DF8180",
    x"33DF6591",
    x"33DF49A6",
    x"33DF2DBF",
    x"33DF11DB",
    x"33DEF5FA",
    x"33DEDA1D",
    x"33DEBE44",
    x"33DEA26E",
    x"33DE869B",
    x"33DE6ACC",
    x"33DE4F00",
    x"33DE3338",
    x"33DE1774",
    x"33DDFBB2",
    x"33DDDFF5",
    x"33DDC43A",
    x"33DDA884",
    x"33DD8CD0",
    x"33DD7120",
    x"33DD5574",
    x"33DD39CB",
    x"33DD1E26",
    x"33DD0283",
    x"33DCE6E5",
    x"33DCCB4A",
    x"33DCAFB2",
    x"33DC941E",
    x"33DC788D",
    x"33DC5D00",
    x"33DC4176",
    x"33DC25EF",
    x"33DC0A6C",
    x"33DBEEED",
    x"33DBD371",
    x"33DBB7F8",
    x"33DB9C83",
    x"33DB8111",
    x"33DB65A2",
    x"33DB4A37",
    x"33DB2ED0",
    x"33DB136C",
    x"33DAF80B",
    x"33DADCAE",
    x"33DAC154",
    x"33DAA5FD",
    x"33DA8AAA",
    x"33DA6F5B",
    x"33DA540E",
    x"33DA38C6",
    x"33DA1D80",
    x"33DA023E",
    x"33D9E700",
    x"33D9CBC4",
    x"33D9B08D",
    x"33D99558",
    x"33D97A27",
    x"33D95EFA",
    x"33D943D0",
    x"33D928A9",
    x"33D90D85",
    x"33D8F265",
    x"33D8D749",
    x"33D8BC30",
    x"33D8A11A",
    x"33D88607",
    x"33D86AF8",
    x"33D84FED",
    x"33D834E4",
    x"33D819DF",
    x"33D7FEDE",
    x"33D7E3E0",
    x"33D7C8E5",
    x"33D7ADED",
    x"33D792F9",
    x"33D77809",
    x"33D75D1B",
    x"33D74231",
    x"33D7274B",
    x"33D70C68",
    x"33D6F188",
    x"33D6D6AB",
    x"33D6BBD2",
    x"33D6A0FC",
    x"33D6862A",
    x"33D66B5B",
    x"33D6508F",
    x"33D635C7",
    x"33D61B02",
    x"33D60040",
    x"33D5E581",
    x"33D5CAC6",
    x"33D5B00F",
    x"33D5955A",
    x"33D57AA9",
    x"33D55FFC",
    x"33D54551",
    x"33D52AAA",
    x"33D51007",
    x"33D4F566",
    x"33D4DAC9",
    x"33D4C030",
    x"33D4A599",
    x"33D48B06",
    x"33D47077",
    x"33D455EA",
    x"33D43B61",
    x"33D420DB",
    x"33D40659",
    x"33D3EBDA",
    x"33D3D15E",
    x"33D3B6E5",
    x"33D39C70",
    x"33D381FE",
    x"33D36790",
    x"33D34D24",
    x"33D332BC",
    x"33D31858",
    x"33D2FDF6",
    x"33D2E398",
    x"33D2C93D",
    x"33D2AEE6",
    x"33D29492",
    x"33D27A41",
    x"33D25FF3",
    x"33D245A9",
    x"33D22B62",
    x"33D2111E",
    x"33D1F6DD",
    x"33D1DCA0",
    x"33D1C266",
    x"33D1A830",
    x"33D18DFC",
    x"33D173CC",
    x"33D1599F",
    x"33D13F76",
    x"33D1254F",
    x"33D10B2C",
    x"33D0F10D",
    x"33D0D6F0",
    x"33D0BCD7",
    x"33D0A2C1",
    x"33D088AE",
    x"33D06E9F",
    x"33D05493",
    x"33D03A8A",
    x"33D02084",
    x"33D00682",
    x"33CFEC82",
    x"33CFD286",
    x"33CFB88E",
    x"33CF9E98",
    x"33CF84A6",
    x"33CF6AB7",
    x"33CF50CB",
    x"33CF36E3",
    x"33CF1CFE",
    x"33CF031C",
    x"33CEE93D",
    x"33CECF61",
    x"33CEB589",
    x"33CE9BB4",
    x"33CE81E2",
    x"33CE6813",
    x"33CE4E48",
    x"33CE3480",
    x"33CE1ABB",
    x"33CE00F9",
    x"33CDE73B",
    x"33CDCD7F",
    x"33CDB3C7",
    x"33CD9A12",
    x"33CD8061",
    x"33CD66B2",
    x"33CD4D07",
    x"33CD335F",
    x"33CD19BA",
    x"33CD0019",
    x"33CCE67A",
    x"33CCCCDF",
    x"33CCB347",
    x"33CC99B2",
    x"33CC8021",
    x"33CC6692",
    x"33CC4D07",
    x"33CC337F",
    x"33CC19FA",
    x"33CC0078",
    x"33CBE6FA",
    x"33CBCD7F",
    x"33CBB407",
    x"33CB9A92",
    x"33CB8120",
    x"33CB67B1",
    x"33CB4E46",
    x"33CB34DE",
    x"33CB1B79",
    x"33CB0217",
    x"33CAE8B8",
    x"33CACF5D",
    x"33CAB604",
    x"33CA9CAF",
    x"33CA835D",
    x"33CA6A0E",
    x"33CA50C3",
    x"33CA377A",
    x"33CA1E35",
    x"33CA04F3",
    x"33C9EBB4",
    x"33C9D278",
    x"33C9B93F",
    x"33C9A009",
    x"33C986D7",
    x"33C96DA8",
    x"33C9547C",
    x"33C93B53",
    x"33C9222D",
    x"33C9090A",
    x"33C8EFEB",
    x"33C8D6CE",
    x"33C8BDB5",
    x"33C8A49F",
    x"33C88B8C",
    x"33C8727C",
    x"33C8596F",
    x"33C84065",
    x"33C8275F",
    x"33C80E5C",
    x"33C7F55B",
    x"33C7DC5E",
    x"33C7C364",
    x"33C7AA6D",
    x"33C7917A",
    x"33C77889",
    x"33C75F9C",
    x"33C746B1",
    x"33C72DCA",
    x"33C714E6",
    x"33C6FC05",
    x"33C6E327",
    x"33C6CA4C",
    x"33C6B174",
    x"33C6989F",
    x"33C67FCE",
    x"33C66700",
    x"33C64E34",
    x"33C6356C",
    x"33C61CA7",
    x"33C603E5",
    x"33C5EB26",
    x"33C5D26A",
    x"33C5B9B1",
    x"33C5A0FC",
    x"33C58849",
    x"33C56F9A",
    x"33C556ED",
    x"33C53E44",
    x"33C5259E",
    x"33C50CFA",
    x"33C4F45A",
    x"33C4DBBD",
    x"33C4C323",
    x"33C4AA8D",
    x"33C491F9",
    x"33C47968",
    x"33C460DA",
    x"33C44850",
    x"33C42FC8",
    x"33C41744",
    x"33C3FEC2",
    x"33C3E644",
    x"33C3CDC9",
    x"33C3B551",
    x"33C39CDC",
    x"33C3846A",
    x"33C36BFA",
    x"33C3538F",
    x"33C33B26",
    x"33C322C0",
    x"33C30A5D",
    x"33C2F1FD",
    x"33C2D9A0",
    x"33C2C147",
    x"33C2A8F0",
    x"33C2909D",
    x"33C2784C",
    x"33C25FFE",
    x"33C247B4",
    x"33C22F6D",
    x"33C21728",
    x"33C1FEE7",
    x"33C1E6A8",
    x"33C1CE6D",
    x"33C1B635",
    x"33C19DFF",
    x"33C185CD",
    x"33C16D9E",
    x"33C15572",
    x"33C13D49",
    x"33C12523",
    x"33C10CFF",
    x"33C0F4DF",
    x"33C0DCC2",
    x"33C0C4A8",
    x"33C0AC91",
    x"33C0947D",
    x"33C07C6C",
    x"33C0645E",
    x"33C04C53",
    x"33C0344B",
    x"33C01C46",
    x"33C00444",
    x"33BFEC45",
    x"33BFD449",
    x"33BFBC50",
    x"33BFA45A",
    x"33BF8C67",
    x"33BF7476",
    x"33BF5C89",
    x"33BF449F",
    x"33BF2CB8",
    x"33BF14D4",
    x"33BEFCF3",
    x"33BEE515",
    x"33BECD3A",
    x"33BEB562",
    x"33BE9D8C",
    x"33BE85BA",
    x"33BE6DEB",
    x"33BE561F",
    x"33BE3E55",
    x"33BE268F",
    x"33BE0ECC",
    x"33BDF70B",
    x"33BDDF4E",
    x"33BDC794",
    x"33BDAFDC",
    x"33BD9828",
    x"33BD8076",
    x"33BD68C8",
    x"33BD511C",
    x"33BD3973",
    x"33BD21CE",
    x"33BD0A2B",
    x"33BCF28B",
    x"33BCDAEE",
    x"33BCC354",
    x"33BCABBD",
    x"33BC9429",
    x"33BC7C98",
    x"33BC650A",
    x"33BC4D7F",
    x"33BC35F7",
    x"33BC1E72",
    x"33BC06EF",
    x"33BBEF70",
    x"33BBD7F3",
    x"33BBC07A",
    x"33BBA903",
    x"33BB9190",
    x"33BB7A1F",
    x"33BB62B1",
    x"33BB4B46",
    x"33BB33DE",
    x"33BB1C79",
    x"33BB0517",
    x"33BAEDB8",
    x"33BAD65C",
    x"33BABF02",
    x"33BAA7AC",
    x"33BA9058",
    x"33BA7908",
    x"33BA61BA",
    x"33BA4A6F",
    x"33BA3328",
    x"33BA1BE3",
    x"33BA04A1",
    x"33B9ED61",
    x"33B9D625",
    x"33B9BEEC",
    x"33B9A7B5",
    x"33B99082",
    x"33B97951",
    x"33B96224",
    x"33B94AF9",
    x"33B933D1",
    x"33B91CAC",
    x"33B9058A",
    x"33B8EE6A",
    x"33B8D74E",
    x"33B8C035",
    x"33B8A91E",
    x"33B8920A",
    x"33B87AFA",
    x"33B863EC",
    x"33B84CE1",
    x"33B835D8",
    x"33B81ED3",
    x"33B807D1",
    x"33B7F0D1",
    x"33B7D9D5",
    x"33B7C2DB",
    x"33B7ABE4",
    x"33B794F0",
    x"33B77DFF",
    x"33B76710",
    x"33B75025",
    x"33B7393C",
    x"33B72256",
    x"33B70B74",
    x"33B6F494",
    x"33B6DDB6",
    x"33B6C6DC",
    x"33B6B005",
    x"33B69930",
    x"33B6825E",
    x"33B66B90",
    x"33B654C4",
    x"33B63DFA",
    x"33B62734",
    x"33B61071",
    x"33B5F9B0",
    x"33B5E2F2",
    x"33B5CC37",
    x"33B5B57F",
    x"33B59ECA",
    x"33B58817",
    x"33B57168",
    x"33B55ABB",
    x"33B54411",
    x"33B52D6A",
    x"33B516C6",
    x"33B50024",
    x"33B4E986",
    x"33B4D2EA",
    x"33B4BC51",
    x"33B4A5BB",
    x"33B48F28",
    x"33B47897",
    x"33B46209",
    x"33B44B7F",
    x"33B434F7",
    x"33B41E71",
    x"33B407EF",
    x"33B3F16F",
    x"33B3DAF3",
    x"33B3C479",
    x"33B3AE01",
    x"33B3978D",
    x"33B3811C",
    x"33B36AAD",
    x"33B35441",
    x"33B33DD8",
    x"33B32771",
    x"33B3110E",
    x"33B2FAAD",
    x"33B2E44F",
    x"33B2CDF4",
    x"33B2B79C",
    x"33B2A146",
    x"33B28AF3",
    x"33B274A3",
    x"33B25E56",
    x"33B2480C",
    x"33B231C4",
    x"33B21B7F",
    x"33B2053D",
    x"33B1EEFE",
    x"33B1D8C2",
    x"33B1C288",
    x"33B1AC51",
    x"33B1961D",
    x"33B17FEC",
    x"33B169BD",
    x"33B15391",
    x"33B13D68",
    x"33B12742",
    x"33B1111E",
    x"33B0FAFD",
    x"33B0E4DF",
    x"33B0CEC4",
    x"33B0B8AC",
    x"33B0A296",
    x"33B08C83",
    x"33B07673",
    x"33B06065",
    x"33B04A5B",
    x"33B03453",
    x"33B01E4E",
    x"33B0084B",
    x"33AFF24C",
    x"33AFDC4F",
    x"33AFC655",
    x"33AFB05D",
    x"33AF9A69",
    x"33AF8477",
    x"33AF6E87",
    x"33AF589B",
    x"33AF42B1",
    x"33AF2CCA",
    x"33AF16E6",
    x"33AF0105",
    x"33AEEB26",
    x"33AED54A",
    x"33AEBF70",
    x"33AEA99A",
    x"33AE93C6",
    x"33AE7DF5",
    x"33AE6827",
    x"33AE525B",
    x"33AE3C92",
    x"33AE26CC",
    x"33AE1108",
    x"33ADFB48",
    x"33ADE589",
    x"33ADCFCE",
    x"33ADBA16",
    x"33ADA460",
    x"33AD8EAC",
    x"33AD78FC",
    x"33AD634E",
    x"33AD4DA3",
    x"33AD37FB",
    x"33AD2255",
    x"33AD0CB2",
    x"33ACF712",
    x"33ACE174",
    x"33ACCBDA",
    x"33ACB641",
    x"33ACA0AC",
    x"33AC8B19",
    x"33AC7589",
    x"33AC5FFC",
    x"33AC4A71",
    x"33AC34E9",
    x"33AC1F64",
    x"33AC09E1",
    x"33ABF462",
    x"33ABDEE4",
    x"33ABC96A",
    x"33ABB3F2",
    x"33AB9E7D",
    x"33AB890A",
    x"33AB739B",
    x"33AB5E2D",
    x"33AB48C3",
    x"33AB335B",
    x"33AB1DF6",
    x"33AB0894",
    x"33AAF334",
    x"33AADDD7",
    x"33AAC87D",
    x"33AAB325",
    x"33AA9DD0",
    x"33AA887D",
    x"33AA732E",
    x"33AA5DE1",
    x"33AA4896",
    x"33AA334E",
    x"33AA1E09",
    x"33AA08C7",
    x"33A9F387",
    x"33A9DE4A",
    x"33A9C910",
    x"33A9B3D8",
    x"33A99EA3",
    x"33A98970",
    x"33A97440",
    x"33A95F13",
    x"33A949E9",
    x"33A934C1",
    x"33A91F9B",
    x"33A90A79",
    x"33A8F559",
    x"33A8E03B",
    x"33A8CB21",
    x"33A8B609",
    x"33A8A0F3",
    x"33A88BE0",
    x"33A876D0",
    x"33A861C3",
    x"33A84CB8",
    x"33A837AF",
    x"33A822AA",
    x"33A80DA7",
    x"33A7F8A6",
    x"33A7E3A9",
    x"33A7CEAD",
    x"33A7B9B5",
    x"33A7A4BF",
    x"33A78FCC",
    x"33A77ADB",
    x"33A765ED",
    x"33A75102",
    x"33A73C19",
    x"33A72733",
    x"33A7124F",
    x"33A6FD6E",
    x"33A6E890",
    x"33A6D3B4",
    x"33A6BEDB",
    x"33A6AA04",
    x"33A69530",
    x"33A6805F",
    x"33A66B90",
    x"33A656C4",
    x"33A641FA",
    x"33A62D33",
    x"33A6186F",
    x"33A603AD",
    x"33A5EEEE",
    x"33A5DA32",
    x"33A5C578",
    x"33A5B0C0",
    x"33A59C0B",
    x"33A58759",
    x"33A572AA",
    x"33A55DFD",
    x"33A54952",
    x"33A534AA",
    x"33A52005",
    x"33A50B62",
    x"33A4F6C2",
    x"33A4E225",
    x"33A4CD8A",
    x"33A4B8F1",
    x"33A4A45B",
    x"33A48FC8",
    x"33A47B37",
    x"33A466A9",
    x"33A4521E",
    x"33A43D95",
    x"33A4290E",
    x"33A4148A",
    x"33A40009",
    x"33A3EB8A",
    x"33A3D70E",
    x"33A3C295",
    x"33A3AE1E",
    x"33A399A9",
    x"33A38537",
    x"33A370C8",
    x"33A35C5B",
    x"33A347F1",
    x"33A33389",
    x"33A31F24",
    x"33A30AC1",
    x"33A2F661",
    x"33A2E204",
    x"33A2CDA9",
    x"33A2B950",
    x"33A2A4FA",
    x"33A290A7",
    x"33A27C56",
    x"33A26808",
    x"33A253BC",
    x"33A23F73",
    x"33A22B2C",
    x"33A216E8",
    x"33A202A7",
    x"33A1EE68",
    x"33A1DA2B",
    x"33A1C5F1",
    x"33A1B1BA",
    x"33A19D85",
    x"33A18952",
    x"33A17522",
    x"33A160F5",
    x"33A14CCA",
    x"33A138A2",
    x"33A1247C",
    x"33A11059",
    x"33A0FC38",
    x"33A0E81A",
    x"33A0D3FE",
    x"33A0BFE5",
    x"33A0ABCE",
    x"33A097BA",
    x"33A083A8",
    x"33A06F99",
    x"33A05B8C",
    x"33A04782",
    x"33A0337A",
    x"33A01F75",
    x"33A00B72",
    x"339FF772",
    x"339FE374",
    x"339FCF79",
    x"339FBB80",
    x"339FA78A",
    x"339F9397",
    x"339F7FA5",
    x"339F6BB7",
    x"339F57CA",
    x"339F43E1",
    x"339F2FF9",
    x"339F1C15",
    x"339F0832",
    x"339EF453",
    x"339EE075",
    x"339ECC9B",
    x"339EB8C2",
    x"339EA4EC",
    x"339E9119",
    x"339E7D48",
    x"339E697A",
    x"339E55AE",
    x"339E41E4",
    x"339E2E1D",
    x"339E1A59",
    x"339E0697",
    x"339DF2D7",
    x"339DDF1A",
    x"339DCB5F",
    x"339DB7A7",
    x"339DA3F1",
    x"339D903E",
    x"339D7C8D",
    x"339D68DF",
    x"339D5533",
    x"339D418A",
    x"339D2DE3",
    x"339D1A3E",
    x"339D069C",
    x"339CF2FD",
    x"339CDF5F",
    x"339CCBC5",
    x"339CB82C",
    x"339CA497",
    x"339C9103",
    x"339C7D72",
    x"339C69E4",
    x"339C5658",
    x"339C42CE",
    x"339C2F47",
    x"339C1BC3",
    x"339C0840",
    x"339BF4C1",
    x"339BE143",
    x"339BCDC8",
    x"339BBA50",
    x"339BA6DA",
    x"339B9366",
    x"339B7FF5",
    x"339B6C86",
    x"339B591A",
    x"339B45B0",
    x"339B3248",
    x"339B1EE3",
    x"339B0B80",
    x"339AF820",
    x"339AE4C2",
    x"339AD167",
    x"339ABE0E",
    x"339AAAB8",
    x"339A9763",
    x"339A8412",
    x"339A70C2",
    x"339A5D76",
    x"339A4A2B",
    x"339A36E3",
    x"339A239D",
    x"339A105A",
    x"3399FD19",
    x"3399E9DB",
    x"3399D69F",
    x"3399C365",
    x"3399B02E",
    x"33999CF9",
    x"339989C7",
    x"33997697",
    x"33996369",
    x"3399503E",
    x"33993D15",
    x"339929EF",
    x"339916CA",
    x"339903A9",
    x"3398F08A",
    x"3398DD6D",
    x"3398CA52",
    x"3398B73A",
    x"3398A424",
    x"33989111",
    x"33987E00",
    x"33986AF2",
    x"339857E5",
    x"339844DC",
    x"339831D4",
    x"33981ECF",
    x"33980BCC",
    x"3397F8CC",
    x"3397E5CE",
    x"3397D2D3",
    x"3397BFDA",
    x"3397ACE3",
    x"339799EE",
    x"339786FC",
    x"3397740D",
    x"3397611F",
    x"33974E34",
    x"33973B4C",
    x"33972866",
    x"33971582",
    x"339702A0",
    x"3396EFC1",
    x"3396DCE4",
    x"3396CA0A",
    x"3396B732",
    x"3396A45C",
    x"33969189",
    x"33967EB8",
    x"33966BE9",
    x"3396591D",
    x"33964653",
    x"3396338B",
    x"339620C6",
    x"33960E03",
    x"3395FB42",
    x"3395E884",
    x"3395D5C8",
    x"3395C30F",
    x"3395B057",
    x"33959DA2",
    x"33958AF0",
    x"33957840",
    x"33956592",
    x"339552E6",
    x"3395403D",
    x"33952D96",
    x"33951AF2",
    x"33950850",
    x"3394F5B0",
    x"3394E312",
    x"3394D077",
    x"3394BDDE",
    x"3394AB47",
    x"339498B3",
    x"33948621",
    x"33947392",
    x"33946104",
    x"33944E79",
    x"33943BF1",
    x"3394296A",
    x"339416E6",
    x"33940465",
    x"3393F1E5",
    x"3393DF68",
    x"3393CCED",
    x"3393BA75",
    x"3393A7FF",
    x"3393958B",
    x"33938319",
    x"339370AA",
    x"33935E3D",
    x"33934BD3",
    x"3393396A",
    x"33932704",
    x"339314A1",
    x"3393023F",
    x"3392EFE0",
    x"3392DD83",
    x"3392CB29",
    x"3392B8D0",
    x"3392A67A",
    x"33929427",
    x"339281D5",
    x"33926F86",
    x"33925D3A",
    x"33924AEF",
    x"339238A7",
    x"33922661",
    x"3392141D",
    x"339201DC",
    x"3391EF9D",
    x"3391DD60",
    x"3391CB25",
    x"3391B8ED",
    x"3391A6B7",
    x"33919483",
    x"33918252",
    x"33917023",
    x"33915DF6",
    x"33914BCB",
    x"339139A3",
    x"3391277D",
    x"33911559",
    x"33910338",
    x"3390F118",
    x"3390DEFB",
    x"3390CCE1",
    x"3390BAC8",
    x"3390A8B2",
    x"3390969E",
    x"3390848C",
    x"3390727D",
    x"33906070",
    x"33904E65",
    x"33903C5C",
    x"33902A56",
    x"33901851",
    x"33900650",
    x"338FF450",
    x"338FE252",
    x"338FD057",
    x"338FBE5E",
    x"338FAC68",
    x"338F9A73",
    x"338F8881",
    x"338F7691",
    x"338F64A3",
    x"338F52B8",
    x"338F40CF",
    x"338F2EE8",
    x"338F1D03",
    x"338F0B21",
    x"338EF940",
    x"338EE762",
    x"338ED586",
    x"338EC3AD",
    x"338EB1D5",
    x"338EA000",
    x"338E8E2D",
    x"338E7C5D",
    x"338E6A8E",
    x"338E58C2",
    x"338E46F8",
    x"338E3530",
    x"338E236B",
    x"338E11A8",
    x"338DFFE6",
    x"338DEE28",
    x"338DDC6B",
    x"338DCAB1",
    x"338DB8F8",
    x"338DA742",
    x"338D958E",
    x"338D83DD",
    x"338D722D",
    x"338D6080",
    x"338D4ED5",
    x"338D3D2D",
    x"338D2B86",
    x"338D19E2",
    x"338D0840",
    x"338CF6A0",
    x"338CE502",
    x"338CD366",
    x"338CC1CD",
    x"338CB036",
    x"338C9EA1",
    x"338C8D0E",
    x"338C7B7E",
    x"338C69EF",
    x"338C5863",
    x"338C46D9",
    x"338C3552",
    x"338C23CC",
    x"338C1249",
    x"338C00C7",
    x"338BEF48",
    x"338BDDCC",
    x"338BCC51",
    x"338BBAD9",
    x"338BA962",
    x"338B97EE",
    x"338B867C",
    x"338B750D",
    x"338B639F",
    x"338B5234",
    x"338B40CA",
    x"338B2F63",
    x"338B1DFF",
    x"338B0C9C",
    x"338AFB3B",
    x"338AE9DD",
    x"338AD881",
    x"338AC727",
    x"338AB5CF",
    x"338AA47A",
    x"338A9326",
    x"338A81D5",
    x"338A7086",
    x"338A5F39",
    x"338A4DEE",
    x"338A3CA5",
    x"338A2B5F",
    x"338A1A1A",
    x"338A08D8",
    x"3389F798",
    x"3389E65A",
    x"3389D51F",
    x"3389C3E5",
    x"3389B2AE",
    x"3389A178",
    x"33899045",
    x"33897F14",
    x"33896DE5",
    x"33895CB9",
    x"33894B8E",
    x"33893A66",
    x"33892940",
    x"3389181C",
    x"338906FA",
    x"3388F5DA",
    x"3388E4BC",
    x"3388D3A1",
    x"3388C287",
    x"3388B170",
    x"3388A05B",
    x"33888F48",
    x"33887E37",
    x"33886D28",
    x"33885C1C",
    x"33884B11",
    x"33883A09",
    x"33882903",
    x"338817FF",
    x"338806FD",
    x"3387F5FD",
    x"3387E4FF",
    x"3387D404",
    x"3387C30A",
    x"3387B213",
    x"3387A11E",
    x"3387902B",
    x"33877F3A",
    x"33876E4B",
    x"33875D5E",
    x"33874C74",
    x"33873B8B",
    x"33872AA5",
    x"338719C0",
    x"338708DE",
    x"3386F7FE",
    x"3386E720",
    x"3386D644",
    x"3386C56B",
    x"3386B493",
    x"3386A3BE",
    x"338692EA",
    x"33868219",
    x"3386714A",
    x"3386607C",
    x"33864FB1",
    x"33863EE9",
    x"33862E22",
    x"33861D5D",
    x"33860C9A",
    x"3385FBDA",
    x"3385EB1B",
    x"3385DA5F",
    x"3385C9A5",
    x"3385B8ED",
    x"3385A837",
    x"33859783",
    x"338586D1",
    x"33857621",
    x"33856573",
    x"338554C8",
    x"3385441E",
    x"33853377",
    x"338522D1",
    x"3385122E",
    x"3385018D",
    x"3384F0ED",
    x"3384E050",
    x"3384CFB5",
    x"3384BF1C",
    x"3384AE86",
    x"33849DF1",
    x"33848D5E",
    x"33847CCD",
    x"33846C3F",
    x"33845BB2",
    x"33844B28",
    x"33843AA0",
    x"33842A19",
    x"33841995",
    x"33840913",
    x"3383F893",
    x"3383E815",
    x"3383D799",
    x"3383C71F",
    x"3383B6A7",
    x"3383A631",
    x"338395BD",
    x"3383854C",
    x"338374DC",
    x"3383646F",
    x"33835403",
    x"3383439A",
    x"33833332",
    x"338322CD",
    x"33831269",
    x"33830208",
    x"3382F1A9",
    x"3382E14C",
    x"3382D0F1",
    x"3382C098",
    x"3382B040",
    x"33829FEB",
    x"33828F98",
    x"33827F48",
    x"33826EF9",
    x"33825EAC",
    x"33824E61",
    x"33823E18",
    x"33822DD1",
    x"33821D8D",
    x"33820D4A",
    x"3381FD09",
    x"3381ECCB",
    x"3381DC8E",
    x"3381CC54",
    x"3381BC1B",
    x"3381ABE5",
    x"33819BB0",
    x"33818B7E",
    x"33817B4D",
    x"33816B1F",
    x"33815AF3",
    x"33814AC8",
    x"33813AA0",
    x"33812A7A",
    x"33811A55",
    x"33810A33",
    x"3380FA13",
    x"3380E9F4",
    x"3380D9D8",
    x"3380C9BE",
    x"3380B9A6",
    x"3380A990",
    x"3380997B",
    x"33808969",
    x"33807959",
    x"3380694B",
    x"3380593F",
    x"33804935",
    x"3380392C",
    x"33802926",
    x"33801922",
    x"33800920",
    x"337FF240",
    x"337FD243",
    x"337FB24B",
    x"337F9257",
    x"337F7266",
    x"337F527A",
    x"337F3292",
    x"337F12AE",
    x"337EF2CD",
    x"337ED2F1",
    x"337EB318",
    x"337E9344",
    x"337E7374",
    x"337E53A7",
    x"337E33DF",
    x"337E141A",
    x"337DF45A",
    x"337DD49D",
    x"337DB4E5",
    x"337D9530",
    x"337D757F",
    x"337D55D3",
    x"337D362A",
    x"337D1685",
    x"337CF6E4",
    x"337CD747",
    x"337CB7AE",
    x"337C9819",
    x"337C7888",
    x"337C58FB",
    x"337C3972",
    x"337C19ED",
    x"337BFA6C",
    x"337BDAEE",
    x"337BBB75",
    x"337B9BFF",
    x"337B7C8E",
    x"337B5D20",
    x"337B3DB7",
    x"337B1E51",
    x"337AFEEF",
    x"337ADF91",
    x"337AC037",
    x"337AA0E1",
    x"337A818F",
    x"337A6241",
    x"337A42F6",
    x"337A23B0",
    x"337A046D",
    x"3379E52F",
    x"3379C5F4",
    x"3379A6BD",
    x"3379878A",
    x"3379685B",
    x"33794930",
    x"33792A09",
    x"33790AE6",
    x"3378EBC6",
    x"3378CCAB",
    x"3378AD93",
    x"33788E7F",
    x"33786F70",
    x"33785064",
    x"3378315B",
    x"33781257",
    x"3377F357",
    x"3377D45A",
    x"3377B562",
    x"3377966D",
    x"3377777C",
    x"3377588F",
    x"337739A6",
    x"33771AC1",
    x"3376FBDF",
    x"3376DD02",
    x"3376BE28",
    x"33769F52",
    x"33768080",
    x"337661B2",
    x"337642E8",
    x"33762421",
    x"3376055F",
    x"3375E6A0",
    x"3375C7E5",
    x"3375A92E",
    x"33758A7B",
    x"33756BCB",
    x"33754D20",
    x"33752E78",
    x"33750FD4",
    x"3374F134",
    x"3374D298",
    x"3374B400",
    x"3374956B",
    x"337476DA",
    x"3374584D",
    x"337439C4",
    x"33741B3F",
    x"3373FCBD",
    x"3373DE40",
    x"3373BFC6",
    x"3373A150",
    x"337382DD",
    x"3373646F",
    x"33734604",
    x"3373279D",
    x"3373093A",
    x"3372EADB",
    x"3372CC80",
    x"3372AE28",
    x"33728FD4",
    x"33727184",
    x"33725338",
    x"337234EF",
    x"337216AB",
    x"3371F86A",
    x"3371DA2C",
    x"3371BBF3",
    x"33719DBD",
    x"33717F8C",
    x"3371615E",
    x"33714333",
    x"3371250D",
    x"337106EA",
    x"3370E8CB",
    x"3370CAB0",
    x"3370AC98",
    x"33708E85",
    x"33707075",
    x"33705269",
    x"33703460",
    x"3370165B",
    x"336FF85B",
    x"336FDA5D",
    x"336FBC64",
    x"336F9E6E",
    x"336F807C",
    x"336F628E",
    x"336F44A4",
    x"336F26BD",
    x"336F08DA",
    x"336EEAFB",
    x"336ECD1F",
    x"336EAF48",
    x"336E9173",
    x"336E73A3",
    x"336E55D7",
    x"336E380E",
    x"336E1A49",
    x"336DFC87",
    x"336DDEC9",
    x"336DC10F",
    x"336DA359",
    x"336D85A7",
    x"336D67F8",
    x"336D4A4D",
    x"336D2CA5",
    x"336D0F01",
    x"336CF161",
    x"336CD3C5",
    x"336CB62C",
    x"336C9898",
    x"336C7B06",
    x"336C5D79",
    x"336C3FEF",
    x"336C2269",
    x"336C04E6",
    x"336BE768",
    x"336BC9EC",
    x"336BAC75",
    x"336B8F01",
    x"336B7191",
    x"336B5425",
    x"336B36BC",
    x"336B1957",
    x"336AFBF6",
    x"336ADE98",
    x"336AC13E",
    x"336AA3E8",
    x"336A8695",
    x"336A6946",
    x"336A4BFB",
    x"336A2EB3",
    x"336A116F",
    x"3369F42F",
    x"3369D6F2",
    x"3369B9B9",
    x"33699C84",
    x"33697F52",
    x"33696224",
    x"336944FA",
    x"336927D3",
    x"33690AB0",
    x"3368ED90",
    x"3368D074",
    x"3368B35C",
    x"33689647",
    x"33687936",
    x"33685C29",
    x"33683F1F",
    x"33682219",
    x"33680517",
    x"3367E818",
    x"3367CB1D",
    x"3367AE25",
    x"33679131",
    x"33677441",
    x"33675754",
    x"33673A6B",
    x"33671D86",
    x"336700A4",
    x"3366E3C5",
    x"3366C6EB",
    x"3366AA14",
    x"33668D40",
    x"33667070",
    x"336653A4",
    x"336636DC",
    x"33661A16",
    x"3365FD55",
    x"3365E097",
    x"3365C3DD",
    x"3365A726",
    x"33658A73",
    x"33656DC4",
    x"33655118",
    x"3365346F",
    x"336517CB",
    x"3364FB29",
    x"3364DE8C",
    x"3364C1F2",
    x"3364A55B",
    x"336488C8",
    x"33646C39",
    x"33644FAD",
    x"33643325",
    x"336416A1",
    x"3363FA1F",
    x"3363DDA2",
    x"3363C128",
    x"3363A4B2",
    x"3363883F",
    x"33636BD0",
    x"33634F64",
    x"336332FC",
    x"33631697",
    x"3362FA36",
    x"3362DDD9",
    x"3362C17F",
    x"3362A528",
    x"336288D5",
    x"33626C86",
    x"3362503A",
    x"336233F2",
    x"336217AD",
    x"3361FB6C",
    x"3361DF2E",
    x"3361C2F4",
    x"3361A6BE",
    x"33618A8B",
    x"33616E5B",
    x"3361522F",
    x"33613606",
    x"336119E1",
    x"3360FDC0",
    x"3360E1A2",
    x"3360C588",
    x"3360A971",
    x"33608D5D",
    x"3360714D",
    x"33605541",
    x"33603938",
    x"33601D33",
    x"33600131",
    x"335FE532",
    x"335FC937",
    x"335FAD40",
    x"335F914C",
    x"335F755C",
    x"335F596F",
    x"335F3D85",
    x"335F219F",
    x"335F05BD",
    x"335EE9DE",
    x"335ECE02",
    x"335EB22A",
    x"335E9656",
    x"335E7A85",
    x"335E5EB7",
    x"335E42ED",
    x"335E2727",
    x"335E0B63",
    x"335DEFA4",
    x"335DD3E7",
    x"335DB82F",
    x"335D9C79",
    x"335D80C8",
    x"335D6519",
    x"335D496E",
    x"335D2DC7",
    x"335D1223",
    x"335CF682",
    x"335CDAE5",
    x"335CBF4C",
    x"335CA3B5",
    x"335C8823",
    x"335C6C93",
    x"335C5108",
    x"335C357F",
    x"335C19FA",
    x"335BFE79",
    x"335BE2FB",
    x"335BC780",
    x"335BAC09",
    x"335B9095",
    x"335B7525",
    x"335B59B8",
    x"335B3E4E",
    x"335B22E8",
    x"335B0785",
    x"335AEC26",
    x"335AD0CA",
    x"335AB572",
    x"335A9A1D",
    x"335A7ECB",
    x"335A637D",
    x"335A4833",
    x"335A2CEB",
    x"335A11A7",
    x"3359F667",
    x"3359DB2A",
    x"3359BFF0",
    x"3359A4BA",
    x"33598987",
    x"33596E57",
    x"3359532B",
    x"33593803",
    x"33591CDD",
    x"335901BB",
    x"3358E69D",
    x"3358CB82",
    x"3358B06A",
    x"33589556",
    x"33587A45",
    x"33585F37",
    x"3358442D",
    x"33582926",
    x"33580E23",
    x"3357F322",
    x"3357D826",
    x"3357BD2C",
    x"3357A236",
    x"33578744",
    x"33576C55",
    x"33575169",
    x"33573680",
    x"33571B9B",
    x"335700B9",
    x"3356E5DB",
    x"3356CB00",
    x"3356B028",
    x"33569554",
    x"33567A83",
    x"33565FB5",
    x"335644EB",
    x"33562A24",
    x"33560F60",
    x"3355F4A0",
    x"3355D9E3",
    x"3355BF2A",
    x"3355A473",
    x"335589C1",
    x"33556F11",
    x"33555465",
    x"335539BC",
    x"33551F16",
    x"33550474",
    x"3354E9D5",
    x"3354CF3A",
    x"3354B4A1",
    x"33549A0D",
    x"33547F7B",
    x"335464ED",
    x"33544A62",
    x"33542FDA",
    x"33541556",
    x"3353FAD5",
    x"3353E057",
    x"3353C5DD",
    x"3353AB66",
    x"335390F2",
    x"33537681",
    x"33535C14",
    x"335341AA",
    x"33532744",
    x"33530CE1",
    x"3352F281",
    x"3352D824",
    x"3352BDCB",
    x"3352A374",
    x"33528922",
    x"33526ED2",
    x"33525486",
    x"33523A3D",
    x"33521FF7",
    x"335205B5",
    x"3351EB76",
    x"3351D13A",
    x"3351B702",
    x"33519CCC",
    x"3351829A",
    x"3351686C",
    x"33514E40",
    x"33513418",
    x"335119F3",
    x"3350FFD2",
    x"3350E5B3",
    x"3350CB98",
    x"3350B180",
    x"3350976C",
    x"33507D5B",
    x"3350634D",
    x"33504942",
    x"33502F3A",
    x"33501536",
    x"334FFB35",
    x"334FE137",
    x"334FC73D",
    x"334FAD45",
    x"334F9351",
    x"334F7961",
    x"334F5F73",
    x"334F4589",
    x"334F2BA2",
    x"334F11BE",
    x"334EF7DD",
    x"334EDE00",
    x"334EC426",
    x"334EAA4F",
    x"334E907B",
    x"334E76AB",
    x"334E5CDD",
    x"334E4313",
    x"334E294D",
    x"334E0F89",
    x"334DF5C9",
    x"334DDC0C",
    x"334DC252",
    x"334DA89B",
    x"334D8EE8",
    x"334D7537",
    x"334D5B8A",
    x"334D41E0",
    x"334D283A",
    x"334D0E96",
    x"334CF4F6",
    x"334CDB59",
    x"334CC1BF",
    x"334CA829",
    x"334C8E95",
    x"334C7505",
    x"334C5B78",
    x"334C41EE",
    x"334C2868",
    x"334C0EE4",
    x"334BF564",
    x"334BDBE7",
    x"334BC26D",
    x"334BA8F6",
    x"334B8F83",
    x"334B7612",
    x"334B5CA5",
    x"334B433B",
    x"334B29D4",
    x"334B1071",
    x"334AF710",
    x"334ADDB3",
    x"334AC459",
    x"334AAB02",
    x"334A91AE",
    x"334A785D",
    x"334A5F10",
    x"334A45C6",
    x"334A2C7E",
    x"334A133A",
    x"3349F9FA",
    x"3349E0BC",
    x"3349C781",
    x"3349AE4A",
    x"33499516",
    x"33497BE5",
    x"334962B7",
    x"3349498C",
    x"33493065",
    x"33491740",
    x"3348FE1F",
    x"3348E501",
    x"3348CBE5",
    x"3348B2CE",
    x"334899B9",
    x"334880A7",
    x"33486799",
    x"33484E8D",
    x"33483585",
    x"33481C80",
    x"3348037E",
    x"3347EA7F",
    x"3347D183",
    x"3347B88B",
    x"33479F95",
    x"334786A3",
    x"33476DB3",
    x"334754C7",
    x"33473BDE",
    x"334722F8",
    x"33470A15",
    x"3346F136",
    x"3346D859",
    x"3346BF80",
    x"3346A6A9",
    x"33468DD6",
    x"33467506",
    x"33465C39",
    x"3346436F",
    x"33462AA8",
    x"334611E4",
    x"3345F923",
    x"3345E066",
    x"3345C7AB",
    x"3345AEF4",
    x"33459640",
    x"33457D8E",
    x"334564E0",
    x"33454C35",
    x"3345338D",
    x"33451AE8",
    x"33450246",
    x"3344E9A8",
    x"3344D10C",
    x"3344B873",
    x"33449FDE",
    x"3344874B",
    x"33446EBC",
    x"33445630",
    x"33443DA7",
    x"33442520",
    x"33440C9D",
    x"3343F41D",
    x"3343DBA0",
    x"3343C326",
    x"3343AAAF",
    x"3343923C",
    x"334379CB",
    x"3343615D",
    x"334348F3",
    x"3343308B",
    x"33431826",
    x"3342FFC5",
    x"3342E766",
    x"3342CF0B",
    x"3342B6B3",
    x"33429E5D",
    x"3342860B",
    x"33426DBC",
    x"33425570",
    x"33423D27",
    x"334224E0",
    x"33420C9D",
    x"3341F45D",
    x"3341DC20",
    x"3341C3E6",
    x"3341ABAF",
    x"3341937B",
    x"33417B4A",
    x"3341631C",
    x"33414AF2",
    x"334132CA",
    x"33411AA5",
    x"33410283",
    x"3340EA64",
    x"3340D248",
    x"3340BA30",
    x"3340A21A",
    x"33408A07",
    x"334071F7",
    x"334059EB",
    x"334041E1",
    x"334029DA",
    x"334011D6",
    x"333FF9D6",
    x"333FE1D8",
    x"333FC9DD",
    x"333FB1E6",
    x"333F99F1",
    x"333F81FF",
    x"333F6A10",
    x"333F5225",
    x"333F3A3C",
    x"333F2256",
    x"333F0A73",
    x"333EF293",
    x"333EDAB7",
    x"333EC2DD",
    x"333EAB06",
    x"333E9332",
    x"333E7B61",
    x"333E6393",
    x"333E4BC8",
    x"333E3400",
    x"333E1C3B",
    x"333E0479",
    x"333DECBA",
    x"333DD4FE",
    x"333DBD45",
    x"333DA58F",
    x"333D8DDB",
    x"333D762B",
    x"333D5E7E",
    x"333D46D3",
    x"333D2F2C",
    x"333D1788",
    x"333CFFE6",
    x"333CE848",
    x"333CD0AC",
    x"333CB914",
    x"333CA17E",
    x"333C89EB",
    x"333C725B",
    x"333C5ACF",
    x"333C4345",
    x"333C2BBE",
    x"333C143A",
    x"333BFCB9",
    x"333BE53B",
    x"333BCDBF",
    x"333BB647",
    x"333B9ED2",
    x"333B875F",
    x"333B6FF0",
    x"333B5883",
    x"333B411A",
    x"333B29B3",
    x"333B124F",
    x"333AFAEF",
    x"333AE391",
    x"333ACC36",
    x"333AB4DE",
    x"333A9D88",
    x"333A8636",
    x"333A6EE7",
    x"333A579B",
    x"333A4051",
    x"333A290A",
    x"333A11C7",
    x"3339FA86",
    x"3339E348",
    x"3339CC0D",
    x"3339B4D5",
    x"33399DA0",
    x"3339866E",
    x"33396F3E",
    x"33395812",
    x"333940E8",
    x"333929C2",
    x"3339129E",
    x"3338FB7D",
    x"3338E45F",
    x"3338CD44",
    x"3338B62C",
    x"33389F16",
    x"33388804",
    x"333870F4",
    x"333859E8",
    x"333842DE",
    x"33382BD7",
    x"333814D3",
    x"3337FDD2",
    x"3337E6D4",
    x"3337CFD8",
    x"3337B8E0",
    x"3337A1EA",
    x"33378AF7",
    x"33377407",
    x"33375D1A",
    x"33374630",
    x"33372F49",
    x"33371864",
    x"33370182",
    x"3336EAA4",
    x"3336D3C8",
    x"3336BCEF",
    x"3336A619",
    x"33368F45",
    x"33367875",
    x"333661A7",
    x"33364ADC",
    x"33363414",
    x"33361D4F",
    x"3336068D",
    x"3335EFCE",
    x"3335D911",
    x"3335C257",
    x"3335ABA0",
    x"333594EC",
    x"33357E3B",
    x"3335678D",
    x"333550E1",
    x"33353A39",
    x"33352393",
    x"33350CF0",
    x"3334F650",
    x"3334DFB2",
    x"3334C918",
    x"3334B280",
    x"33349BEB",
    x"33348559",
    x"33346ECA",
    x"3334583D",
    x"333441B4",
    x"33342B2D",
    x"333414A9",
    x"3333FE28",
    x"3333E7A9",
    x"3333D12E",
    x"3333BAB5",
    x"3333A43F",
    x"33338DCC",
    x"3333775C",
    x"333360EE",
    x"33334A83",
    x"3333341B",
    x"33331DB6",
    x"33330754",
    x"3332F0F5",
    x"3332DA98",
    x"3332C43E",
    x"3332ADE7",
    x"33329792",
    x"33328141",
    x"33326AF2",
    x"333254A6",
    x"33323E5D",
    x"33322817",
    x"333211D3",
    x"3331FB92",
    x"3331E554",
    x"3331CF19",
    x"3331B8E0",
    x"3331A2AB",
    x"33318C78",
    x"33317647",
    x"3331601A",
    x"333149EF",
    x"333133C8",
    x"33311DA2",
    x"33310780",
    x"3330F161",
    x"3330DB44",
    x"3330C52A",
    x"3330AF12",
    x"333098FE",
    x"333082EC",
    x"33306CDD",
    x"333056D1",
    x"333040C8",
    x"33302AC1",
    x"333014BD",
    x"332FFEBC",
    x"332FE8BD",
    x"332FD2C1",
    x"332FBCC8",
    x"332FA6D2",
    x"332F90DF",
    x"332F7AEE",
    x"332F6500",
    x"332F4F15",
    x"332F392C",
    x"332F2346",
    x"332F0D63",
    x"332EF783",
    x"332EE1A6",
    x"332ECBCB",
    x"332EB5F3",
    x"332EA01D",
    x"332E8A4B",
    x"332E747B",
    x"332E5EAD",
    x"332E48E3",
    x"332E331B",
    x"332E1D56",
    x"332E0794",
    x"332DF1D4",
    x"332DDC17",
    x"332DC65D",
    x"332DB0A6",
    x"332D9AF1",
    x"332D853F",
    x"332D6F90",
    x"332D59E3",
    x"332D4439",
    x"332D2E92",
    x"332D18EE",
    x"332D034C",
    x"332CEDAD",
    x"332CD811",
    x"332CC277",
    x"332CACE0",
    x"332C974C",
    x"332C81BA",
    x"332C6C2B",
    x"332C569F",
    x"332C4116",
    x"332C2B8F",
    x"332C160B",
    x"332C0089",
    x"332BEB0B",
    x"332BD58E",
    x"332BC015",
    x"332BAA9E",
    x"332B952A",
    x"332B7FB9",
    x"332B6A4B",
    x"332B54DF",
    x"332B3F75",
    x"332B2A0F",
    x"332B14AB",
    x"332AFF4A",
    x"332AE9EB",
    x"332AD48F",
    x"332ABF36",
    x"332AA9DF",
    x"332A948B",
    x"332A7F3A",
    x"332A69EC",
    x"332A54A0",
    x"332A3F56",
    x"332A2A10",
    x"332A14CC",
    x"3329FF8B",
    x"3329EA4C",
    x"3329D510",
    x"3329BFD7",
    x"3329AAA0",
    x"3329956C",
    x"3329803B",
    x"33296B0C",
    x"332955E0",
    x"332940B7",
    x"33292B90",
    x"3329166C",
    x"3329014A",
    x"3328EC2B",
    x"3328D70F",
    x"3328C1F6",
    x"3328ACDF",
    x"332897CA",
    x"332882B9",
    x"33286DAA",
    x"3328589D",
    x"33284394",
    x"33282E8C",
    x"33281988",
    x"33280486",
    x"3327EF87",
    x"3327DA8A",
    x"3327C590",
    x"3327B099",
    x"33279BA4",
    x"332786B2",
    x"332771C2",
    x"33275CD5",
    x"332747EB",
    x"33273303",
    x"33271E1E",
    x"3327093C",
    x"3326F45C",
    x"3326DF7F",
    x"3326CAA4",
    x"3326B5CC",
    x"3326A0F7",
    x"33268C24",
    x"33267754",
    x"33266286",
    x"33264DBB",
    x"332638F3",
    x"3326242D",
    x"33260F6A",
    x"3325FAA9",
    x"3325E5EB",
    x"3325D12F",
    x"3325BC77",
    x"3325A7C0",
    x"3325930D",
    x"33257E5C",
    x"332569AD",
    x"33255501",
    x"33254058",
    x"33252BB1",
    x"3325170D",
    x"3325026B",
    x"3324EDCC",
    x"3324D930",
    x"3324C496",
    x"3324AFFF",
    x"33249B6A",
    x"332486D8",
    x"33247248",
    x"33245DBB",
    x"33244931",
    x"332434A9",
    x"33242024",
    x"33240BA1",
    x"3323F721",
    x"3323E2A3",
    x"3323CE28",
    x"3323B9B0",
    x"3323A53A",
    x"332390C6",
    x"33237C56",
    x"332367E7",
    x"3323537C",
    x"33233F12",
    x"33232AAC",
    x"33231648",
    x"332301E6",
    x"3322ED87",
    x"3322D92B",
    x"3322C4D1",
    x"3322B07A",
    x"33229C25",
    x"332287D3",
    x"33227383",
    x"33225F36",
    x"33224AEB",
    x"332236A3",
    x"3322225D",
    x"33220E1A",
    x"3321F9DA",
    x"3321E59C",
    x"3321D160",
    x"3321BD28",
    x"3321A8F1",
    x"332194BD",
    x"3321808C",
    x"33216C5D",
    x"33215831",
    x"33214407",
    x"33212FE0",
    x"33211BBB",
    x"33210799",
    x"3320F379",
    x"3320DF5C",
    x"3320CB41",
    x"3320B729",
    x"3320A314",
    x"33208F01",
    x"33207AF0",
    x"332066E2",
    x"332052D6",
    x"33203ECD",
    x"33202AC6",
    x"332016C2",
    x"332002C1",
    x"331FEEC2",
    x"331FDAC5",
    x"331FC6CB",
    x"331FB2D3",
    x"331F9EDE",
    x"331F8AEC",
    x"331F76FC",
    x"331F630E",
    x"331F4F23",
    x"331F3B3A",
    x"331F2754",
    x"331F1370",
    x"331EFF8F",
    x"331EEBB0",
    x"331ED7D4",
    x"331EC3FA",
    x"331EB023",
    x"331E9C4E",
    x"331E887C",
    x"331E74AC",
    x"331E60DF",
    x"331E4D14",
    x"331E394C",
    x"331E2586",
    x"331E11C2",
    x"331DFE01",
    x"331DEA43",
    x"331DD687",
    x"331DC2CD",
    x"331DAF16",
    x"331D9B61",
    x"331D87AF",
    x"331D7400",
    x"331D6052",
    x"331D4CA7",
    x"331D38FF",
    x"331D2559",
    x"331D11B6",
    x"331CFE15",
    x"331CEA76",
    x"331CD6DA",
    x"331CC340",
    x"331CAFA9",
    x"331C9C15",
    x"331C8882",
    x"331C74F2",
    x"331C6165",
    x"331C4DDA",
    x"331C3A52",
    x"331C26CC",
    x"331C1348",
    x"331BFFC7",
    x"331BEC48",
    x"331BD8CC",
    x"331BC552",
    x"331BB1DA",
    x"331B9E65",
    x"331B8AF3",
    x"331B7783",
    x"331B6415",
    x"331B50AA",
    x"331B3D41",
    x"331B29DA",
    x"331B1676",
    x"331B0315",
    x"331AEFB5",
    x"331ADC59",
    x"331AC8FE",
    x"331AB5A6",
    x"331AA251",
    x"331A8EFE",
    x"331A7BAD",
    x"331A685F",
    x"331A5513",
    x"331A41CA",
    x"331A2E83",
    x"331A1B3E",
    x"331A07FC",
    x"3319F4BC",
    x"3319E17F",
    x"3319CE44",
    x"3319BB0B",
    x"3319A7D5",
    x"331994A1",
    x"33198170",
    x"33196E41",
    x"33195B14",
    x"331947EA",
    x"331934C2",
    x"3319219D",
    x"33190E7A",
    x"3318FB59",
    x"3318E83B",
    x"3318D51F",
    x"3318C206",
    x"3318AEEF",
    x"33189BDA",
    x"331888C8",
    x"331875B8",
    x"331862AA",
    x"33184F9F",
    x"33183C96",
    x"33182990",
    x"3318168C",
    x"3318038A",
    x"3317F08B",
    x"3317DD8E",
    x"3317CA94",
    x"3317B79C",
    x"3317A4A6",
    x"331791B2",
    x"33177EC1",
    x"33176BD3",
    x"331758E6",
    x"331745FC",
    x"33173315",
    x"33172030",
    x"33170D4D",
    x"3316FA6C",
    x"3316E78E",
    x"3316D4B2",
    x"3316C1D9",
    x"3316AF02",
    x"33169C2D",
    x"3316895B",
    x"3316768B",
    x"331663BD",
    x"331650F2",
    x"33163E29",
    x"33162B62",
    x"3316189E",
    x"331605DC",
    x"3315F31D",
    x"3315E060",
    x"3315CDA5",
    x"3315BAEC",
    x"3315A836",
    x"33159582",
    x"331582D1",
    x"33157021",
    x"33155D75",
    x"33154ACA",
    x"33153822",
    x"3315257C",
    x"331512D8",
    x"33150037",
    x"3314ED98",
    x"3314DAFC",
    x"3314C862",
    x"3314B5CA",
    x"3314A334",
    x"331490A1",
    x"33147E10",
    x"33146B81",
    x"331458F5",
    x"3314466B",
    x"331433E4",
    x"3314215E",
    x"33140EDB",
    x"3313FC5B",
    x"3313E9DC",
    x"3313D760",
    x"3313C4E6",
    x"3313B26F",
    x"33139FFA",
    x"33138D87",
    x"33137B16",
    x"331368A8",
    x"3313563C",
    x"331343D3",
    x"3313316B",
    x"33131F06",
    x"33130CA3",
    x"3312FA43",
    x"3312E7E5",
    x"3312D589",
    x"3312C32F",
    x"3312B0D8",
    x"33129E83",
    x"33128C31",
    x"331279E0",
    x"33126792",
    x"33125546",
    x"331242FD",
    x"331230B6",
    x"33121E71",
    x"33120C2E",
    x"3311F9EE",
    x"3311E7AF",
    x"3311D574",
    x"3311C33A",
    x"3311B103",
    x"33119ECE",
    x"33118C9B",
    x"33117A6B",
    x"3311683D",
    x"33115611",
    x"331143E7",
    x"331131C0",
    x"33111F9B",
    x"33110D78",
    x"3310FB57",
    x"3310E939",
    x"3310D71D",
    x"3310C503",
    x"3310B2EC",
    x"3310A0D6",
    x"33108EC3",
    x"33107CB3",
    x"33106AA4",
    x"33105898",
    x"3310468E",
    x"33103486",
    x"33102281",
    x"3310107E",
    x"330FFE7D",
    x"330FEC7E",
    x"330FDA82",
    x"330FC888",
    x"330FB690",
    x"330FA49A",
    x"330F92A6",
    x"330F80B5",
    x"330F6EC6",
    x"330F5CDA",
    x"330F4AEF",
    x"330F3907",
    x"330F2721",
    x"330F153D",
    x"330F035C",
    x"330EF17C",
    x"330EDF9F",
    x"330ECDC4",
    x"330EBBEC",
    x"330EAA15",
    x"330E9841",
    x"330E866F",
    x"330E74A0",
    x"330E62D2",
    x"330E5107",
    x"330E3F3E",
    x"330E2D77",
    x"330E1BB2",
    x"330E09F0",
    x"330DF830",
    x"330DE672",
    x"330DD4B6",
    x"330DC2FD",
    x"330DB146",
    x"330D9F91",
    x"330D8DDE",
    x"330D7C2D",
    x"330D6A7F",
    x"330D58D2",
    x"330D4728",
    x"330D3581",
    x"330D23DB",
    x"330D1238",
    x"330D0097",
    x"330CEEF8",
    x"330CDD5B",
    x"330CCBC0",
    x"330CBA28",
    x"330CA892",
    x"330C96FE",
    x"330C856C",
    x"330C73DC",
    x"330C624F",
    x"330C50C4",
    x"330C3F3B",
    x"330C2DB4",
    x"330C1C2F",
    x"330C0AAD",
    x"330BF92D",
    x"330BE7AF",
    x"330BD633",
    x"330BC4B9",
    x"330BB342",
    x"330BA1CC",
    x"330B9059",
    x"330B7EE8",
    x"330B6D79",
    x"330B5C0D",
    x"330B4AA2",
    x"330B393A",
    x"330B27D4",
    x"330B1670",
    x"330B050F",
    x"330AF3AF",
    x"330AE252",
    x"330AD0F6",
    x"330ABF9D",
    x"330AAE46",
    x"330A9CF2",
    x"330A8B9F",
    x"330A7A4F",
    x"330A6901",
    x"330A57B5",
    x"330A466B",
    x"330A3523",
    x"330A23DD",
    x"330A129A",
    x"330A0159",
    x"3309F01A",
    x"3309DEDD",
    x"3309CDA2",
    x"3309BC69",
    x"3309AB33",
    x"330999FF",
    x"330988CC",
    x"3309779C",
    x"3309666E",
    x"33095543",
    x"33094419",
    x"330932F2",
    x"330921CC",
    x"330910A9",
    x"3308FF88",
    x"3308EE69",
    x"3308DD4D",
    x"3308CC32",
    x"3308BB1A",
    x"3308AA03",
    x"330898EF",
    x"330887DD",
    x"330876CD",
    x"330865BF",
    x"330854B4",
    x"330843AA",
    x"330832A3",
    x"3308219E",
    x"3308109A",
    x"3307FF99",
    x"3307EE9A",
    x"3307DD9E",
    x"3307CCA3",
    x"3307BBAB",
    x"3307AAB4",
    x"330799C0",
    x"330788CE",
    x"330777DE",
    x"330766F0",
    x"33075604",
    x"3307451A",
    x"33073433",
    x"3307234D",
    x"3307126A",
    x"33070189",
    x"3306F0A9",
    x"3306DFCC",
    x"3306CEF2",
    x"3306BE19",
    x"3306AD42",
    x"33069C6D",
    x"33068B9B",
    x"33067ACA",
    x"330669FC",
    x"33065930",
    x"33064866",
    x"3306379E",
    x"330626D8",
    x"33061614",
    x"33060552",
    x"3305F493",
    x"3305E3D5",
    x"3305D31A",
    x"3305C261",
    x"3305B1A9",
    x"3305A0F4",
    x"33059041",
    x"33057F90",
    x"33056EE1",
    x"33055E34",
    x"33054D8A",
    x"33053CE1",
    x"33052C3A",
    x"33051B96",
    x"33050AF3",
    x"3304FA53",
    x"3304E9B5",
    x"3304D919",
    x"3304C87F",
    x"3304B7E7",
    x"3304A751",
    x"330496BD",
    x"3304862B",
    x"3304759B",
    x"3304650E",
    x"33045482",
    x"330443F8",
    x"33043371",
    x"330422EC",
    x"33041268",
    x"330401E7",
    x"3303F168",
    x"3303E0EB",
    x"3303D070",
    x"3303BFF7",
    x"3303AF80",
    x"33039F0B",
    x"33038E98",
    x"33037E27",
    x"33036DB8",
    x"33035D4C",
    x"33034CE1",
    x"33033C78",
    x"33032C12",
    x"33031BAD",
    x"33030B4B",
    x"3302FAEB",
    x"3302EA8C",
    x"3302DA30",
    x"3302C9D6",
    x"3302B97D",
    x"3302A927",
    x"330298D3",
    x"33028881",
    x"33027831",
    x"330267E3",
    x"33025797",
    x"3302474D",
    x"33023705",
    x"330226BF",
    x"3302167C",
    x"3302063A",
    x"3301F5FA",
    x"3301E5BC",
    x"3301D581",
    x"3301C547",
    x"3301B50F",
    x"3301A4DA",
    x"330194A6",
    x"33018474",
    x"33017445",
    x"33016417",
    x"330153EC",
    x"330143C2",
    x"3301339B",
    x"33012375",
    x"33011352",
    x"33010331",
    x"3300F311",
    x"3300E2F4",
    x"3300D2D9",
    x"3300C2BF",
    x"3300B2A8",
    x"3300A293",
    x"3300927F",
    x"3300826E",
    x"3300725F",
    x"33006251",
    x"33005246",
    x"3300423D",
    x"33003235",
    x"33002230",
    x"3300122D",
    x"3300022C",
    x"32FFE459",
    x"32FFC45E",
    x"32FFA468",
    x"32FF8475",
    x"32FF6486",
    x"32FF449C",
    x"32FF24B5",
    x"32FF04D3",
    x"32FEE4F4",
    x"32FEC51A",
    x"32FEA543",
    x"32FE8570",
    x"32FE65A1",
    x"32FE45D7",
    x"32FE2610",
    x"32FE064D",
    x"32FDE68E",
    x"32FDC6D4",
    x"32FDA71D",
    x"32FD876A",
    x"32FD67BB",
    x"32FD4810",
    x"32FD2869",
    x"32FD08C6",
    x"32FCE927",
    x"32FCC98C",
    x"32FCA9F4",
    x"32FC8A61",
    x"32FC6AD2",
    x"32FC4B46",
    x"32FC2BBF",
    x"32FC0C3B",
    x"32FBECBC",
    x"32FBCD40",
    x"32FBADC9",
    x"32FB8E55",
    x"32FB6EE5",
    x"32FB4F79",
    x"32FB3011",
    x"32FB10AD",
    x"32FAF14D",
    x"32FAD1F1",
    x"32FAB298",
    x"32FA9344",
    x"32FA73F4",
    x"32FA54A7",
    x"32FA355E",
    x"32FA161A",
    x"32F9F6D9",
    x"32F9D79C",
    x"32F9B863",
    x"32F9992E",
    x"32F979FD",
    x"32F95ACF",
    x"32F93BA6",
    x"32F91C80",
    x"32F8FD5F",
    x"32F8DE41",
    x"32F8BF27",
    x"32F8A011",
    x"32F880FF",
    x"32F861F1",
    x"32F842E7",
    x"32F823E0",
    x"32F804DE",
    x"32F7E5DF",
    x"32F7C6E4",
    x"32F7A7ED",
    x"32F788FA",
    x"32F76A0B",
    x"32F74B20",
    x"32F72C38",
    x"32F70D55",
    x"32F6EE75",
    x"32F6CF99",
    x"32F6B0C1",
    x"32F691ED",
    x"32F6731D",
    x"32F65450",
    x"32F63588",
    x"32F616C3",
    x"32F5F802",
    x"32F5D945",
    x"32F5BA8C",
    x"32F59BD6",
    x"32F57D25",
    x"32F55E77",
    x"32F53FCD",
    x"32F52127",
    x"32F50285",
    x"32F4E3E6",
    x"32F4C54C",
    x"32F4A6B5",
    x"32F48822",
    x"32F46993",
    x"32F44B08",
    x"32F42C80",
    x"32F40DFD",
    x"32F3EF7D",
    x"32F3D101",
    x"32F3B288",
    x"32F39414",
    x"32F375A3",
    x"32F35737",
    x"32F338CE",
    x"32F31A68",
    x"32F2FC07",
    x"32F2DDA9",
    x"32F2BF50",
    x"32F2A0FA",
    x"32F282A7",
    x"32F26459",
    x"32F2460E",
    x"32F227C7",
    x"32F20984",
    x"32F1EB45",
    x"32F1CD0A",
    x"32F1AED2",
    x"32F1909E",
    x"32F1726E",
    x"32F15441",
    x"32F13619",
    x"32F117F4",
    x"32F0F9D3",
    x"32F0DBB5",
    x"32F0BD9C",
    x"32F09F86",
    x"32F08174",
    x"32F06365",
    x"32F0455B",
    x"32F02754",
    x"32F00951",
    x"32EFEB52",
    x"32EFCD56",
    x"32EFAF5E",
    x"32EF916A",
    x"32EF737A",
    x"32EF558E",
    x"32EF37A5",
    x"32EF19C0",
    x"32EEFBDE",
    x"32EEDE01",
    x"32EEC027",
    x"32EEA251",
    x"32EE847E",
    x"32EE66B0",
    x"32EE48E5",
    x"32EE2B1D",
    x"32EE0D5A",
    x"32EDEF9A",
    x"32EDD1DE",
    x"32EDB425",
    x"32ED9671",
    x"32ED78C0",
    x"32ED5B13",
    x"32ED3D69",
    x"32ED1FC3",
    x"32ED0221",
    x"32ECE483",
    x"32ECC6E8",
    x"32ECA951",
    x"32EC8BBE",
    x"32EC6E2E",
    x"32EC50A2",
    x"32EC331A",
    x"32EC1595",
    x"32EBF815",
    x"32EBDA97",
    x"32EBBD1E",
    x"32EB9FA8",
    x"32EB8236",
    x"32EB64C8",
    x"32EB475D",
    x"32EB29F6",
    x"32EB0C92",
    x"32EAEF33",
    x"32EAD1D6",
    x"32EAB47E",
    x"32EA9729",
    x"32EA79D8",
    x"32EA5C8B",
    x"32EA3F41",
    x"32EA21FB",
    x"32EA04B9",
    x"32E9E77A",
    x"32E9CA3F",
    x"32E9AD07",
    x"32E98FD4",
    x"32E972A3",
    x"32E95577",
    x"32E9384E",
    x"32E91B29",
    x"32E8FE07",
    x"32E8E0E9",
    x"32E8C3CF",
    x"32E8A6B8",
    x"32E889A5",
    x"32E86C96",
    x"32E84F8A",
    x"32E83282",
    x"32E8157E",
    x"32E7F87D",
    x"32E7DB7F",
    x"32E7BE86",
    x"32E7A190",
    x"32E7849D",
    x"32E767AF",
    x"32E74AC3",
    x"32E72DDC",
    x"32E710F8",
    x"32E6F418",
    x"32E6D73B",
    x"32E6BA62",
    x"32E69D8C",
    x"32E680BB",
    x"32E663EC",
    x"32E64722",
    x"32E62A5A",
    x"32E60D97",
    x"32E5F0D7",
    x"32E5D41B",
    x"32E5B762",
    x"32E59AAD",
    x"32E57DFB",
    x"32E5614D",
    x"32E544A3",
    x"32E527FC",
    x"32E50B59",
    x"32E4EEB9",
    x"32E4D21D",
    x"32E4B585",
    x"32E498F0",
    x"32E47C5F",
    x"32E45FD1",
    x"32E44347",
    x"32E426C0",
    x"32E40A3D",
    x"32E3EDBD",
    x"32E3D142",
    x"32E3B4C9",
    x"32E39854",
    x"32E37BE3",
    x"32E35F75",
    x"32E3430B",
    x"32E326A5",
    x"32E30A42",
    x"32E2EDE2",
    x"32E2D186",
    x"32E2B52E",
    x"32E298D9",
    x"32E27C87",
    x"32E2603A",
    x"32E243EF",
    x"32E227A9",
    x"32E20B65",
    x"32E1EF26",
    x"32E1D2EA",
    x"32E1B6B1",
    x"32E19A7C",
    x"32E17E4A",
    x"32E1621C",
    x"32E145F2",
    x"32E129CB",
    x"32E10DA7",
    x"32E0F188",
    x"32E0D56B",
    x"32E0B952",
    x"32E09D3D",
    x"32E0812B",
    x"32E0651C",
    x"32E04912",
    x"32E02D0A",
    x"32E01106",
    x"32DFF506",
    x"32DFD909",
    x"32DFBD10",
    x"32DFA11A",
    x"32DF8527",
    x"32DF6939",
    x"32DF4D4D",
    x"32DF3165",
    x"32DF1581",
    x"32DEF9A0",
    x"32DEDDC2",
    x"32DEC1E8",
    x"32DEA612",
    x"32DE8A3F",
    x"32DE6E6F",
    x"32DE52A3",
    x"32DE36DB",
    x"32DE1B16",
    x"32DDFF54",
    x"32DDE396",
    x"32DDC7DB",
    x"32DDAC24",
    x"32DD9070",
    x"32DD74C0",
    x"32DD5913",
    x"32DD3D69",
    x"32DD21C3",
    x"32DD0621",
    x"32DCEA82",
    x"32DCCEE6",
    x"32DCB34E",
    x"32DC97B9",
    x"32DC7C28",
    x"32DC609A",
    x"32DC4510",
    x"32DC2989",
    x"32DC0E06",
    x"32DBF286",
    x"32DBD709",
    x"32DBBB90",
    x"32DBA01A",
    x"32DB84A8",
    x"32DB6939",
    x"32DB4DCE",
    x"32DB3266",
    x"32DB1701",
    x"32DAFBA0",
    x"32DAE042",
    x"32DAC4E8",
    x"32DAA991",
    x"32DA8E3D",
    x"32DA72ED",
    x"32DA57A1",
    x"32DA3C57",
    x"32DA2112",
    x"32DA05CF",
    x"32D9EA90",
    x"32D9CF54",
    x"32D9B41C",
    x"32D998E7",
    x"32D97DB6",
    x"32D96288",
    x"32D9475D",
    x"32D92C36",
    x"32D91112",
    x"32D8F5F2",
    x"32D8DAD5",
    x"32D8BFBB",
    x"32D8A4A5",
    x"32D88992",
    x"32D86E83",
    x"32D85376",
    x"32D8386E",
    x"32D81D68",
    x"32D80266",
    x"32D7E768",
    x"32D7CC6C",
    x"32D7B175",
    x"32D79680",
    x"32D77B8F",
    x"32D760A1",
    x"32D745B7",
    x"32D72AD0",
    x"32D70FEC",
    x"32D6F50C",
    x"32D6DA2F",
    x"32D6BF55",
    x"32D6A47F",
    x"32D689AC",
    x"32D66EDD",
    x"32D65410",
    x"32D63948",
    x"32D61E82",
    x"32D603C0",
    x"32D5E901",
    x"32D5CE46",
    x"32D5B38E",
    x"32D598D9",
    x"32D57E27",
    x"32D56379",
    x"32D548CE",
    x"32D52E27",
    x"32D51383",
    x"32D4F8E2",
    x"32D4DE45",
    x"32D4C3AB",
    x"32D4A914",
    x"32D48E80",
    x"32D473F0",
    x"32D45963",
    x"32D43EDA",
    x"32D42454",
    x"32D409D1",
    x"32D3EF51",
    x"32D3D4D5",
    x"32D3BA5C",
    x"32D39FE6",
    x"32D38574",
    x"32D36B05",
    x"32D35099",
    x"32D33631",
    x"32D31BCC",
    x"32D3016A",
    x"32D2E70B",
    x"32D2CCB0",
    x"32D2B258",
    x"32D29804",
    x"32D27DB2",
    x"32D26364",
    x"32D24919",
    x"32D22ED2",
    x"32D2148E",
    x"32D1FA4D",
    x"32D1E00F",
    x"32D1C5D5",
    x"32D1AB9E",
    x"32D1916A",
    x"32D17739",
    x"32D15D0C",
    x"32D142E2",
    x"32D128BB",
    x"32D10E98",
    x"32D0F478",
    x"32D0DA5B",
    x"32D0C041",
    x"32D0A62B",
    x"32D08C17",
    x"32D07208",
    x"32D057FB",
    x"32D03DF2",
    x"32D023EB",
    x"32D009E9",
    x"32CFEFE9",
    x"32CFD5ED",
    x"32CFBBF4",
    x"32CFA1FE",
    x"32CF880B",
    x"32CF6E1C",
    x"32CF542F",
    x"32CF3A47",
    x"32CF2061",
    x"32CF067E",
    x"32CEEC9F",
    x"32CED2C3",
    x"32CEB8EB",
    x"32CE9F15",
    x"32CE8543",
    x"32CE6B74",
    x"32CE51A8",
    x"32CE37DF",
    x"32CE1E1A",
    x"32CE0458",
    x"32CDEA99",
    x"32CDD0DD",
    x"32CDB725",
    x"32CD9D6F",
    x"32CD83BD",
    x"32CD6A0E",
    x"32CD5063",
    x"32CD36BA",
    x"32CD1D15",
    x"32CD0373",
    x"32CCE9D4",
    x"32CCD039",
    x"32CCB6A0",
    x"32CC9D0B",
    x"32CC8379",
    x"32CC69EA",
    x"32CC505E",
    x"32CC36D6",
    x"32CC1D51",
    x"32CC03CF",
    x"32CBEA50",
    x"32CBD0D4",
    x"32CBB75C",
    x"32CB9DE6",
    x"32CB8474",
    x"32CB6B05",
    x"32CB5199",
    x"32CB3831",
    x"32CB1ECB",
    x"32CB0569",
    x"32CAEC0A",
    x"32CAD2AE",
    x"32CAB955",
    x"32CAA000",
    x"32CA86AD",
    x"32CA6D5E",
    x"32CA5412",
    x"32CA3AC9",
    x"32CA2183",
    x"32CA0841",
    x"32C9EF01",
    x"32C9D5C5",
    x"32C9BC8C",
    x"32C9A356",
    x"32C98A23",
    x"32C970F3",
    x"32C957C7",
    x"32C93E9D",
    x"32C92577",
    x"32C90C54",
    x"32C8F334",
    x"32C8DA17",
    x"32C8C0FD",
    x"32C8A7E7",
    x"32C88ED3",
    x"32C875C3",
    x"32C85CB6",
    x"32C843AC",
    x"32C82AA5",
    x"32C811A1",
    x"32C7F8A1",
    x"32C7DFA3",
    x"32C7C6A9",
    x"32C7ADB1",
    x"32C794BD",
    x"32C77BCC",
    x"32C762DE",
    x"32C749F4",
    x"32C7310C",
    x"32C71827",
    x"32C6FF46",
    x"32C6E668",
    x"32C6CD8C",
    x"32C6B4B4",
    x"32C69BDF",
    x"32C6830D",
    x"32C66A3E",
    x"32C65173",
    x"32C638AA",
    x"32C61FE4",
    x"32C60722",
    x"32C5EE63",
    x"32C5D5A6",
    x"32C5BCED",
    x"32C5A437",
    x"32C58B84",
    x"32C572D4",
    x"32C55A27",
    x"32C5417E",
    x"32C528D7",
    x"32C51034",
    x"32C4F793",
    x"32C4DEF6",
    x"32C4C65B",
    x"32C4ADC4",
    x"32C49530",
    x"32C47C9F",
    x"32C46411",
    x"32C44B86",
    x"32C432FE",
    x"32C41A79",
    x"32C401F7",
    x"32C3E978",
    x"32C3D0FD",
    x"32C3B884",
    x"32C3A00F",
    x"32C3879C",
    x"32C36F2D",
    x"32C356C0",
    x"32C33E57",
    x"32C325F1",
    x"32C30D8E",
    x"32C2F52D",
    x"32C2DCD0",
    x"32C2C476",
    x"32C2AC1F",
    x"32C293CB",
    x"32C27B7A",
    x"32C2632C",
    x"32C24AE1",
    x"32C2329A",
    x"32C21A55",
    x"32C20213",
    x"32C1E9D4",
    x"32C1D199",
    x"32C1B960",
    x"32C1A12A",
    x"32C188F8",
    x"32C170C8",
    x"32C1589B",
    x"32C14072",
    x"32C1284B",
    x"32C11028",
    x"32C0F807",
    x"32C0DFEA",
    x"32C0C7CF",
    x"32C0AFB8",
    x"32C097A3",
    x"32C07F92",
    x"32C06783",
    x"32C04F78",
    x"32C03770",
    x"32C01F6A",
    x"32C00768",
    x"32BFEF68",
    x"32BFD76C",
    x"32BFBF72",
    x"32BFA77C",
    x"32BF8F89",
    x"32BF7798",
    x"32BF5FAB",
    x"32BF47C0",
    x"32BF2FD9",
    x"32BF17F4",
    x"32BF0013",
    x"32BEE834",
    x"32BED059",
    x"32BEB880",
    x"32BEA0AB",
    x"32BE88D8",
    x"32BE7108",
    x"32BE593C",
    x"32BE4172",
    x"32BE29AB",
    x"32BE11E8",
    x"32BDFA27",
    x"32BDE269",
    x"32BDCAAE",
    x"32BDB2F6",
    x"32BD9B42",
    x"32BD8390",
    x"32BD6BE1",
    x"32BD5435",
    x"32BD3C8C",
    x"32BD24E6",
    x"32BD0D42",
    x"32BCF5A2",
    x"32BCDE05",
    x"32BCC66B",
    x"32BCAED3",
    x"32BC973F",
    x"32BC7FAE",
    x"32BC681F",
    x"32BC5094",
    x"32BC390B",
    x"32BC2185",
    x"32BC0A03",
    x"32BBF283",
    x"32BBDB06",
    x"32BBC38C",
    x"32BBAC15",
    x"32BB94A1",
    x"32BB7D30",
    x"32BB65C2",
    x"32BB4E56",
    x"32BB36EE",
    x"32BB1F89",
    x"32BB0826",
    x"32BAF0C7",
    x"32BAD96A",
    x"32BAC210",
    x"32BAAABA",
    x"32BA9366",
    x"32BA7C15",
    x"32BA64C7",
    x"32BA4D7B",
    x"32BA3633",
    x"32BA1EEE",
    x"32BA07AC",
    x"32B9F06C",
    x"32B9D92F",
    x"32B9C1F6",
    x"32B9AABF",
    x"32B9938B",
    x"32B97C5A",
    x"32B9652C",
    x"32B94E01",
    x"32B936D8",
    x"32B91FB3",
    x"32B90890",
    x"32B8F171",
    x"32B8DA54",
    x"32B8C33A",
    x"32B8AC23",
    x"32B8950F",
    x"32B87DFE",
    x"32B866F0",
    x"32B84FE4",
    x"32B838DC",
    x"32B821D6",
    x"32B80AD3",
    x"32B7F3D3",
    x"32B7DCD6",
    x"32B7C5DC",
    x"32B7AEE5",
    x"32B797F0",
    x"32B780FF",
    x"32B76A10",
    x"32B75324",
    x"32B73C3B",
    x"32B72555",
    x"32B70E72",
    x"32B6F792",
    x"32B6E0B4",
    x"32B6C9DA",
    x"32B6B302",
    x"32B69C2D",
    x"32B6855B",
    x"32B66E8B",
    x"32B657BF",
    x"32B640F6",
    x"32B62A2F",
    x"32B6136B",
    x"32B5FCAA",
    x"32B5E5EC",
    x"32B5CF30",
    x"32B5B878",
    x"32B5A1C2",
    x"32B58B10",
    x"32B57460",
    x"32B55DB2",
    x"32B54708",
    x"32B53061",
    x"32B519BC",
    x"32B5031A",
    x"32B4EC7B",
    x"32B4D5DF",
    x"32B4BF46",
    x"32B4A8AF",
    x"32B4921C",
    x"32B47B8B",
    x"32B464FD",
    x"32B44E72",
    x"32B437E9",
    x"32B42164",
    x"32B40AE1",
    x"32B3F461",
    x"32B3DDE4",
    x"32B3C769",
    x"32B3B0F2",
    x"32B39A7D",
    x"32B3840B",
    x"32B36D9C",
    x"32B35730",
    x"32B340C6",
    x"32B32A60",
    x"32B313FC",
    x"32B2FD9B",
    x"32B2E73C",
    x"32B2D0E1",
    x"32B2BA88",
    x"32B2A432",
    x"32B28DDF",
    x"32B2778F",
    x"32B26141",
    x"32B24AF6",
    x"32B234AE",
    x"32B21E69",
    x"32B20827",
    x"32B1F1E7",
    x"32B1DBAA",
    x"32B1C570",
    x"32B1AF39",
    x"32B19905",
    x"32B182D3",
    x"32B16CA4",
    x"32B15678",
    x"32B1404E",
    x"32B12A28",
    x"32B11404",
    x"32B0FDE3",
    x"32B0E7C4",
    x"32B0D1A9",
    x"32B0BB90",
    x"32B0A57A",
    x"32B08F66",
    x"32B07956",
    x"32B06348",
    x"32B04D3D",
    x"32B03735",
    x"32B0212F",
    x"32B00B2C",
    x"32AFF52C",
    x"32AFDF2F",
    x"32AFC935",
    x"32AFB33D",
    x"32AF9D48",
    x"32AF8756",
    x"32AF7166",
    x"32AF5B79",
    x"32AF458F",
    x"32AF2FA8",
    x"32AF19C3",
    x"32AF03E1",
    x"32AEEE02",
    x"32AED826",
    x"32AEC24C",
    x"32AEAC75",
    x"32AE96A1",
    x"32AE80D0",
    x"32AE6B01",
    x"32AE5535",
    x"32AE3F6C",
    x"32AE29A5",
    x"32AE13E1",
    x"32ADFE20",
    x"32ADE862",
    x"32ADD2A6",
    x"32ADBCED",
    x"32ADA737",
    x"32AD9183",
    x"32AD7BD2",
    x"32AD6624",
    x"32AD5079",
    x"32AD3AD0",
    x"32AD252A",
    x"32AD0F87",
    x"32ACF9E6",
    x"32ACE448",
    x"32ACCEAD",
    x"32ACB915",
    x"32ACA37F",
    x"32AC8DEC",
    x"32AC785B",
    x"32AC62CE",
    x"32AC4D43",
    x"32AC37BA",
    x"32AC2235",
    x"32AC0CB2",
    x"32ABF732",
    x"32ABE1B4",
    x"32ABCC39",
    x"32ABB6C1",
    x"32ABA14B",
    x"32AB8BD9",
    x"32AB7669",
    x"32AB60FB",
    x"32AB4B90",
    x"32AB3628",
    x"32AB20C3",
    x"32AB0B60",
    x"32AAF600",
    x"32AAE0A2",
    x"32AACB48",
    x"32AAB5F0",
    x"32AAA09A",
    x"32AA8B47",
    x"32AA75F7",
    x"32AA60AA",
    x"32AA4B5F",
    x"32AA3617",
    x"32AA20D2",
    x"32AA0B8F",
    x"32A9F64F",
    x"32A9E111",
    x"32A9CBD7",
    x"32A9B69E",
    x"32A9A169",
    x"32A98C36",
    x"32A97706",
    x"32A961D8",
    x"32A94CAD",
    x"32A93785",
    x"32A92260",
    x"32A90D3D",
    x"32A8F81C",
    x"32A8E2FF",
    x"32A8CDE3",
    x"32A8B8CB",
    x"32A8A3B5",
    x"32A88EA2",
    x"32A87992",
    x"32A86484",
    x"32A84F78",
    x"32A83A70",
    x"32A8256A",
    x"32A81066",
    x"32A7FB66",
    x"32A7E668",
    x"32A7D16C",
    x"32A7BC73",
    x"32A7A77D",
    x"32A79289",
    x"32A77D98",
    x"32A768AA",
    x"32A753BE",
    x"32A73ED5",
    x"32A729EF",
    x"32A7150B",
    x"32A70029",
    x"32A6EB4B",
    x"32A6D66E",
    x"32A6C195",
    x"32A6ACBE",
    x"32A697EA",
    x"32A68318",
    x"32A66E49",
    x"32A6597D",
    x"32A644B3",
    x"32A62FEB",
    x"32A61B27",
    x"32A60665",
    x"32A5F1A5",
    x"32A5DCE8",
    x"32A5C82E",
    x"32A5B376",
    x"32A59EC1",
    x"32A58A0E",
    x"32A5755E",
    x"32A560B1",
    x"32A54C06",
    x"32A5375E",
    x"32A522B8",
    x"32A50E15",
    x"32A4F975",
    x"32A4E4D7",
    x"32A4D03C",
    x"32A4BBA3",
    x"32A4A70D",
    x"32A49279",
    x"32A47DE8",
    x"32A4695A",
    x"32A454CE",
    x"32A44044",
    x"32A42BBE",
    x"32A4173A",
    x"32A402B8",
    x"32A3EE39",
    x"32A3D9BC",
    x"32A3C542",
    x"32A3B0CB",
    x"32A39C56",
    x"32A387E4",
    x"32A37374",
    x"32A35F07",
    x"32A34A9D",
    x"32A33634",
    x"32A321CF",
    x"32A30D6C",
    x"32A2F90C",
    x"32A2E4AE",
    x"32A2D052",
    x"32A2BBFA",
    x"32A2A7A3",
    x"32A29350",
    x"32A27EFF",
    x"32A26AB0",
    x"32A25664",
    x"32A2421A",
    x"32A22DD3",
    x"32A2198F",
    x"32A2054D",
    x"32A1F10E",
    x"32A1DCD1",
    x"32A1C896",
    x"32A1B45F",
    x"32A1A029",
    x"32A18BF7",
    x"32A177C6",
    x"32A16399",
    x"32A14F6D",
    x"32A13B45",
    x"32A1271F",
    x"32A112FB",
    x"32A0FEDA",
    x"32A0EABB",
    x"32A0D69F",
    x"32A0C286",
    x"32A0AE6F",
    x"32A09A5A",
    x"32A08648",
    x"32A07238",
    x"32A05E2B",
    x"32A04A21",
    x"32A03619",
    x"32A02213",
    x"32A00E10",
    x"329FFA10",
    x"329FE612",
    x"329FD216",
    x"329FBE1D",
    x"329FAA27",
    x"329F9633",
    x"329F8241",
    x"329F6E52",
    x"329F5A66",
    x"329F467C",
    x"329F3294",
    x"329F1EAF",
    x"329F0ACC",
    x"329EF6EC",
    x"329EE30F",
    x"329ECF34",
    x"329EBB5B",
    x"329EA785",
    x"329E93B1",
    x"329E7FE0",
    x"329E6C11",
    x"329E5845",
    x"329E447B",
    x"329E30B4",
    x"329E1CEF",
    x"329E092C",
    x"329DF56C",
    x"329DE1AF",
    x"329DCDF4",
    x"329DBA3C",
    x"329DA685",
    x"329D92D2",
    x"329D7F21",
    x"329D6B72",
    x"329D57C6",
    x"329D441C",
    x"329D3075",
    x"329D1CD0",
    x"329D092E",
    x"329CF58E",
    x"329CE1F0",
    x"329CCE55",
    x"329CBABD",
    x"329CA727",
    x"329C9393",
    x"329C8002",
    x"329C6C73",
    x"329C58E7",
    x"329C455D",
    x"329C31D5",
    x"329C1E50",
    x"329C0ACE",
    x"329BF74E",
    x"329BE3D0",
    x"329BD055",
    x"329BBCDC",
    x"329BA965",
    x"329B95F1",
    x"329B8280",
    x"329B6F11",
    x"329B5BA4",
    x"329B483A",
    x"329B34D2",
    x"329B216D",
    x"329B0E0A",
    x"329AFAA9",
    x"329AE74B",
    x"329AD3EF",
    x"329AC096",
    x"329AAD3F",
    x"329A99EB",
    x"329A8699",
    x"329A7349",
    x"329A5FFC",
    x"329A4CB1",
    x"329A3969",
    x"329A2623",
    x"329A12DF",
    x"3299FF9E",
    x"3299EC5F",
    x"3299D923",
    x"3299C5E9",
    x"3299B2B1",
    x"32999F7C",
    x"32998C4A",
    x"32997919",
    x"329965EB",
    x"329952C0",
    x"32993F97",
    x"32992C70",
    x"3299194C",
    x"3299062A",
    x"3298F30A",
    x"3298DFED",
    x"3298CCD2",
    x"3298B9BA",
    x"3298A6A4",
    x"32989390",
    x"3298807F",
    x"32986D70",
    x"32985A63",
    x"32984759",
    x"32983451",
    x"3298214C",
    x"32980E49",
    x"3297FB49",
    x"3297E84A",
    x"3297D54E",
    x"3297C255",
    x"3297AF5E",
    x"32979C69",
    x"32978977",
    x"32977687",
    x"32976399",
    x"329750AE",
    x"32973DC5",
    x"32972ADE",
    x"329717FA",
    x"32970518",
    x"3296F239",
    x"3296DF5C",
    x"3296CC81",
    x"3296B9A9",
    x"3296A6D3",
    x"329693FF",
    x"3296812E",
    x"32966E5F",
    x"32965B92",
    x"329648C8",
    x"32963600",
    x"3296233A",
    x"32961077",
    x"3295FDB6",
    x"3295EAF8",
    x"3295D83C",
    x"3295C582",
    x"3295B2CA",
    x"3295A015",
    x"32958D62",
    x"32957AB2",
    x"32956803",
    x"32955558",
    x"329542AE",
    x"32953007",
    x"32951D62",
    x"32950AC0",
    x"3294F81F",
    x"3294E582",
    x"3294D2E6",
    x"3294C04D",
    x"3294ADB6",
    x"32949B21",
    x"3294888F",
    x"329475FF",
    x"32946372",
    x"329450E6",
    x"32943E5D",
    x"32942BD7",
    x"32941953",
    x"329406D0",
    x"3293F451",
    x"3293E1D3",
    x"3293CF58",
    x"3293BCE0",
    x"3293AA69",
    x"329397F5",
    x"32938583",
    x"32937314",
    x"329360A6",
    x"32934E3B",
    x"32933BD3",
    x"3293296C",
    x"32931708",
    x"329304A7",
    x"3292F247",
    x"3292DFEA",
    x"3292CD8F",
    x"3292BB37",
    x"3292A8E1",
    x"3292968D",
    x"3292843B",
    x"329271EB",
    x"32925F9E",
    x"32924D54",
    x"32923B0B",
    x"329228C5",
    x"32921681",
    x"3292043F",
    x"3291F200",
    x"3291DFC3",
    x"3291CD88",
    x"3291BB4F",
    x"3291A919",
    x"329196E5",
    x"329184B3",
    x"32917284",
    x"32916057",
    x"32914E2C",
    x"32913C03",
    x"329129DD",
    x"329117B9",
    x"32910597",
    x"3290F377",
    x"3290E15A",
    x"3290CF3F",
    x"3290BD26",
    x"3290AB10",
    x"329098FB",
    x"329086E9",
    x"329074DA",
    x"329062CC",
    x"329050C1",
    x"32903EB8",
    x"32902CB1",
    x"32901AAD",
    x"329008AB",
    x"328FF6AB",
    x"328FE4AD",
    x"328FD2B1",
    x"328FC0B8",
    x"328FAEC1",
    x"328F9CCD",
    x"328F8ADA",
    x"328F78EA",
    x"328F66FC",
    x"328F5510",
    x"328F4327",
    x"328F313F",
    x"328F1F5A",
    x"328F0D77",
    x"328EFB97",
    x"328EE9B9",
    x"328ED7DD",
    x"328EC603",
    x"328EB42B",
    x"328EA256",
    x"328E9082",
    x"328E7EB1",
    x"328E6CE3",
    x"328E5B16",
    x"328E494C",
    x"328E3784",
    x"328E25BE",
    x"328E13FA",
    x"328E0239",
    x"328DF07A",
    x"328DDEBD",
    x"328DCD02",
    x"328DBB4A",
    x"328DA993",
    x"328D97DF",
    x"328D862D",
    x"328D747E",
    x"328D62D0",
    x"328D5125",
    x"328D3F7C",
    x"328D2DD5",
    x"328D1C31",
    x"328D0A8E",
    x"328CF8EE",
    x"328CE750",
    x"328CD5B4",
    x"328CC41B",
    x"328CB283",
    x"328CA0EE",
    x"328C8F5B",
    x"328C7DCA",
    x"328C6C3B",
    x"328C5AAF",
    x"328C4925",
    x"328C379D",
    x"328C2617",
    x"328C1493",
    x"328C0312",
    x"328BF192",
    x"328BE015",
    x"328BCE9A",
    x"328BBD22",
    x"328BABAB",
    x"328B9A37",
    x"328B88C5",
    x"328B7755",
    x"328B65E7",
    x"328B547B",
    x"328B4312",
    x"328B31AA",
    x"328B2045",
    x"328B0EE2",
    x"328AFD81",
    x"328AEC23",
    x"328ADAC6",
    x"328AC96C",
    x"328AB814",
    x"328AA6BE",
    x"328A956A",
    x"328A8419",
    x"328A72C9",
    x"328A617C",
    x"328A5031",
    x"328A3EE8",
    x"328A2DA1",
    x"328A1C5D",
    x"328A0B1A",
    x"3289F9DA",
    x"3289E89C",
    x"3289D760",
    x"3289C626",
    x"3289B4EE",
    x"3289A3B9",
    x"32899285",
    x"32898154",
    x"32897025",
    x"32895EF8",
    x"32894DCD",
    x"32893CA5",
    x"32892B7E",
    x"32891A5A",
    x"32890937",
    x"3288F817",
    x"3288E6F9",
    x"3288D5DE",
    x"3288C4C4",
    x"3288B3AC",
    x"3288A297",
    x"32889184",
    x"32888073",
    x"32886F64",
    x"32885E57",
    x"32884D4C",
    x"32883C43",
    x"32882B3D",
    x"32881A39",
    x"32880936",
    x"3287F836",
    x"3287E738",
    x"3287D63D",
    x"3287C543",
    x"3287B44B",
    x"3287A356",
    x"32879262",
    x"32878171",
    x"32877082",
    x"32875F95",
    x"32874EAA",
    x"32873DC1",
    x"32872CDB",
    x"32871BF6",
    x"32870B14",
    x"3286FA33",
    x"3286E955",
    x"3286D879",
    x"3286C79F",
    x"3286B6C7",
    x"3286A5F1",
    x"3286951E",
    x"3286844C",
    x"3286737D",
    x"328662AF",
    x"328651E4",
    x"3286411B",
    x"32863054",
    x"32861F8F",
    x"32860ECC",
    x"3285FE0B",
    x"3285ED4C",
    x"3285DC90",
    x"3285CBD5",
    x"3285BB1D",
    x"3285AA66",
    x"328599B2",
    x"32858900",
    x"32857850",
    x"328567A2",
    x"328556F6",
    x"3285464C",
    x"328535A4",
    x"328524FF",
    x"3285145B",
    x"328503BA",
    x"3284F31A",
    x"3284E27D",
    x"3284D1E2",
    x"3284C148",
    x"3284B0B1",
    x"3284A01C",
    x"32848F89",
    x"32847EF8",
    x"32846E69",
    x"32845DDD",
    x"32844D52",
    x"32843CC9",
    x"32842C43",
    x"32841BBE",
    x"32840B3C",
    x"3283FABB",
    x"3283EA3D",
    x"3283D9C1",
    x"3283C947",
    x"3283B8CF",
    x"3283A858",
    x"328397E4",
    x"32838773",
    x"32837703",
    x"32836695",
    x"32835629",
    x"328345BF",
    x"32833558",
    x"328324F2",
    x"3283148E",
    x"3283042D",
    x"3282F3CD",
    x"3282E370",
    x"3282D314",
    x"3282C2BB",
    x"3282B264",
    x"3282A20E",
    x"328291BB",
    x"3282816A",
    x"3282711B",
    x"328260CE",
    x"32825083",
    x"3282403A",
    x"32822FF3",
    x"32821FAE",
    x"32820F6B",
    x"3281FF2A",
    x"3281EEEB",
    x"3281DEAE",
    x"3281CE73",
    x"3281BE3A",
    x"3281AE04",
    x"32819DCF",
    x"32818D9C",
    x"32817D6B",
    x"32816D3D",
    x"32815D10",
    x"32814CE6",
    x"32813CBD",
    x"32812C96",
    x"32811C72",
    x"32810C4F",
    x"3280FC2F",
    x"3280EC10",
    x"3280DBF4",
    x"3280CBD9",
    x"3280BBC1",
    x"3280ABAA",
    x"32809B96",
    x"32808B83",
    x"32807B73",
    x"32806B65",
    x"32805B58",
    x"32804B4E",
    x"32803B45",
    x"32802B3F",
    x"32801B3A",
    x"32800B38",
    x"327FF66F",
    x"327FD673",
    x"327FB67A",
    x"327F9685",
    x"327F7694",
    x"327F56A7",
    x"327F36BE",
    x"327F16DA",
    x"327EF6F9",
    x"327ED71C",
    x"327EB743",
    x"327E976E",
    x"327E779D",
    x"327E57D0",
    x"327E3807",
    x"327E1842",
    x"327DF881",
    x"327DD8C4",
    x"327DB90B",
    x"327D9956",
    x"327D79A5",
    x"327D59F7",
    x"327D3A4E",
    x"327D1AA9",
    x"327CFB07",
    x"327CDB6A",
    x"327CBBD1",
    x"327C9C3B",
    x"327C7CA9",
    x"327C5D1C",
    x"327C3D92",
    x"327C1E0C",
    x"327BFE8B",
    x"327BDF0D",
    x"327BBF93",
    x"327BA01D",
    x"327B80AB",
    x"327B613D",
    x"327B41D3",
    x"327B226C",
    x"327B030A",
    x"327AE3AC",
    x"327AC451",
    x"327AA4FA",
    x"327A85A8",
    x"327A6659",
    x"327A470E",
    x"327A27C7",
    x"327A0884",
    x"3279E945",
    x"3279CA0A",
    x"3279AAD3",
    x"32798B9F",
    x"32796C70",
    x"32794D44",
    x"32792E1C",
    x"32790EF9",
    x"3278EFD9",
    x"3278D0BD",
    x"3278B1A5",
    x"32789290",
    x"32787380",
    x"32785473",
    x"3278356B",
    x"32781666",
    x"3277F765",
    x"3277D868",
    x"3277B96F",
    x"32779A7A",
    x"32777B88",
    x"32775C9B",
    x"32773DB1",
    x"32771ECB",
    x"3276FFEA",
    x"3276E10C",
    x"3276C231",
    x"3276A35B",
    x"32768488",
    x"327665BA",
    x"327646EF",
    x"32762828",
    x"32760965",
    x"3275EAA6",
    x"3275CBEA",
    x"3275AD33",
    x"32758E7F",
    x"32756FCF",
    x"32755123",
    x"3275327B",
    x"327513D6",
    x"3274F536",
    x"3274D699",
    x"3274B800",
    x"3274996B",
    x"32747ADA",
    x"32745C4C",
    x"32743DC3",
    x"32741F3D",
    x"327400BB",
    x"3273E23D",
    x"3273C3C2",
    x"3273A54C",
    x"327386D9",
    x"3273686A",
    x"327349FF",
    x"32732B98",
    x"32730D34",
    x"3272EED4",
    x"3272D078",
    x"3272B220",
    x"327293CC",
    x"3272757B",
    x"3272572F",
    x"327238E6",
    x"32721AA0",
    x"3271FC5F",
    x"3271DE21",
    x"3271BFE7",
    x"3271A1B1",
    x"3271837F",
    x"32716550",
    x"32714726",
    x"327128FF",
    x"32710ADB",
    x"3270ECBC",
    x"3270CEA0",
    x"3270B088",
    x"32709274",
    x"32707464",
    x"32705657",
    x"3270384E",
    x"32701A49",
    x"326FFC47",
    x"326FDE4A",
    x"326FC050",
    x"326FA25A",
    x"326F8467",
    x"326F6679",
    x"326F488E",
    x"326F2AA6",
    x"326F0CC3",
    x"326EEEE3",
    x"326ED107",
    x"326EB32F",
    x"326E955A",
    x"326E778A",
    x"326E59BD",
    x"326E3BF3",
    x"326E1E2E",
    x"326E006C",
    x"326DE2AD",
    x"326DC4F3",
    x"326DA73C",
    x"326D8989",
    x"326D6BDA",
    x"326D4E2E",
    x"326D3086",
    x"326D12E2",
    x"326CF542",
    x"326CD7A5",
    x"326CBA0C",
    x"326C9C76",
    x"326C7EE5",
    x"326C6157",
    x"326C43CC",
    x"326C2646",
    x"326C08C3",
    x"326BEB43",
    x"326BCDC8",
    x"326BB050",
    x"326B92DC",
    x"326B756B",
    x"326B57FE",
    x"326B3A95",
    x"326B1D30",
    x"326AFFCE",
    x"326AE270",
    x"326AC515",
    x"326AA7BF",
    x"326A8A6B",
    x"326A6D1C",
    x"326A4FD0",
    x"326A3288",
    x"326A1543",
    x"3269F803",
    x"3269DAC5",
    x"3269BD8C",
    x"3269A056",
    x"32698324",
    x"326965F5",
    x"326948CA",
    x"32692BA3",
    x"32690E7F",
    x"3268F15F",
    x"3268D443",
    x"3268B72A",
    x"32689A15",
    x"32687D04",
    x"32685FF6",
    x"326842EC",
    x"326825E5",
    x"326808E2",
    x"3267EBE3",
    x"3267CEE7",
    x"3267B1EF",
    x"326794FB",
    x"3267780A",
    x"32675B1D",
    x"32673E33",
    x"3267214D",
    x"3267046B",
    x"3266E78C",
    x"3266CAB1",
    x"3266ADDA",
    x"32669106",
    x"32667435",
    x"32665769",
    x"32663AA0",
    x"32661DDA",
    x"32660118",
    x"3265E45A",
    x"3265C79F",
    x"3265AAE8",
    x"32658E34",
    x"32657184",
    x"326554D8",
    x"3265382F",
    x"32651B8A",
    x"3264FEE8",
    x"3264E24A",
    x"3264C5B0",
    x"3264A919",
    x"32648C85",
    x"32646FF6",
    x"32645369",
    x"326436E1",
    x"32641A5C",
    x"3263FDDA",
    x"3263E15C",
    x"3263C4E2",
    x"3263A86B",
    x"32638BF8",
    x"32636F88",
    x"3263531C",
    x"326336B3",
    x"32631A4E",
    x"3262FDED",
    x"3262E18F",
    x"3262C534",
    x"3262A8DD",
    x"32628C8A",
    x"3262703A",
    x"326253EE",
    x"326237A5",
    x"32621B60",
    x"3261FF1E",
    x"3261E2E0",
    x"3261C6A6",
    x"3261AA6F",
    x"32618E3B",
    x"3261720B",
    x"326155DF",
    x"326139B6",
    x"32611D90",
    x"3261016E",
    x"3260E550",
    x"3260C935",
    x"3260AD1D",
    x"3260910A",
    x"326074F9",
    x"326058EC",
    x"32603CE3",
    x"326020DD",
    x"326004DB",
    x"325FE8DC",
    x"325FCCE1",
    x"325FB0E9",
    x"325F94F4",
    x"325F7903",
    x"325F5D16",
    x"325F412C",
    x"325F2546",
    x"325F0963",
    x"325EED83",
    x"325ED1A7",
    x"325EB5CF",
    x"325E99FA",
    x"325E7E28",
    x"325E625A",
    x"325E4690",
    x"325E2AC9",
    x"325E0F05",
    x"325DF345",
    x"325DD788",
    x"325DBBCF",
    x"325DA019",
    x"325D8467",
    x"325D68B8",
    x"325D4D0D",
    x"325D3165",
    x"325D15C1",
    x"325CFA20",
    x"325CDE82",
    x"325CC2E8",
    x"325CA751",
    x"325C8BBE",
    x"325C702E",
    x"325C54A2",
    x"325C3919",
    x"325C1D94",
    x"325C0212",
    x"325BE693",
    x"325BCB18",
    x"325BAFA1",
    x"325B942C",
    x"325B78BB",
    x"325B5D4E",
    x"325B41E4",
    x"325B267E",
    x"325B0B1B",
    x"325AEFBB",
    x"325AD45F",
    x"325AB906",
    x"325A9DB0",
    x"325A825E",
    x"325A6710",
    x"325A4BC5",
    x"325A307D",
    x"325A1538",
    x"3259F9F8",
    x"3259DEBA",
    x"3259C380",
    x"3259A849",
    x"32598D16",
    x"325971E6",
    x"325956B9",
    x"32593B90",
    x"3259206A",
    x"32590548",
    x"3258EA29",
    x"3258CF0D",
    x"3258B3F5",
    x"325898E1",
    x"32587DCF",
    x"325862C1",
    x"325847B6",
    x"32582CAF",
    x"325811AB",
    x"3257F6AB",
    x"3257DBAE",
    x"3257C0B4",
    x"3257A5BD",
    x"32578ACA",
    x"32576FDB",
    x"325754EE",
    x"32573A05",
    x"32571F20",
    x"3257043E",
    x"3256E95F",
    x"3256CE83",
    x"3256B3AB",
    x"325698D6",
    x"32567E05",
    x"32566337",
    x"3256486C",
    x"32562DA5",
    x"325612E1",
    x"3255F820",
    x"3255DD63",
    x"3255C2A9",
    x"3255A7F2",
    x"32558D3F",
    x"3255728F",
    x"325557E2",
    x"32553D39",
    x"32552293",
    x"325507F0",
    x"3254ED51",
    x"3254D2B5",
    x"3254B81C",
    x"32549D87",
    x"325482F5",
    x"32546866",
    x"32544DDB",
    x"32543353",
    x"325418CE",
    x"3253FE4C",
    x"3253E3CE",
    x"3253C953",
    x"3253AEDC",
    x"32539468",
    x"325379F7",
    x"32535F89",
    x"3253451F",
    x"32532AB8",
    x"32531054",
    x"3252F5F4",
    x"3252DB97",
    x"3252C13D",
    x"3252A6E6",
    x"32528C93",
    x"32527243",
    x"325257F7",
    x"32523DAD",
    x"32522367",
    x"32520924",
    x"3251EEE5",
    x"3251D4A9",
    x"3251BA70",
    x"3251A03A",
    x"32518608",
    x"32516BD9",
    x"325151AD",
    x"32513784",
    x"32511D5F",
    x"3251033D",
    x"3250E91E",
    x"3250CF03",
    x"3250B4EA",
    x"32509AD5",
    x"325080C4",
    x"325066B5",
    x"32504CAA",
    x"325032A2",
    x"3250189D",
    x"324FFE9C",
    x"324FE49E",
    x"324FCAA3",
    x"324FB0AB",
    x"324F96B7",
    x"324F7CC5",
    x"324F62D7",
    x"324F48ED",
    x"324F2F05",
    x"324F1521",
    x"324EFB40",
    x"324EE162",
    x"324EC787",
    x"324EADB0",
    x"324E93DC",
    x"324E7A0B",
    x"324E603E",
    x"324E4673",
    x"324E2CAC",
    x"324E12E8",
    x"324DF927",
    x"324DDF6A",
    x"324DC5AF",
    x"324DABF8",
    x"324D9244",
    x"324D7894",
    x"324D5EE6",
    x"324D453C",
    x"324D2B95",
    x"324D11F1",
    x"324CF850",
    x"324CDEB3",
    x"324CC519",
    x"324CAB82",
    x"324C91EE",
    x"324C785D",
    x"324C5ED0",
    x"324C4546",
    x"324C2BBE",
    x"324C123B",
    x"324BF8BA",
    x"324BDF3C",
    x"324BC5C2",
    x"324BAC4B",
    x"324B92D7",
    x"324B7966",
    x"324B5FF9",
    x"324B468E",
    x"324B2D27",
    x"324B13C3",
    x"324AFA62",
    x"324AE104",
    x"324AC7AA",
    x"324AAE52",
    x"324A94FE",
    x"324A7BAD",
    x"324A625F",
    x"324A4915",
    x"324A2FCD",
    x"324A1689",
    x"3249FD47",
    x"3249E409",
    x"3249CACE",
    x"3249B197",
    x"32499862",
    x"32497F31",
    x"32496602",
    x"32494CD7",
    x"324933AF",
    x"32491A8A",
    x"32490168",
    x"3248E84A",
    x"3248CF2E",
    x"3248B616",
    x"32489D01",
    x"324883EF",
    x"32486AE0",
    x"324851D4",
    x"324838CB",
    x"32481FC6",
    x"324806C3",
    x"3247EDC4",
    x"3247D4C8",
    x"3247BBCF",
    x"3247A2D9",
    x"324789E6",
    x"324770F7",
    x"3247580A",
    x"32473F20",
    x"3247263A",
    x"32470D57",
    x"3246F477",
    x"3246DB9A",
    x"3246C2C0",
    x"3246A9E9",
    x"32469115",
    x"32467845",
    x"32465F77",
    x"324646AD",
    x"32462DE6",
    x"32461522",
    x"3245FC60",
    x"3245E3A2",
    x"3245CAE8",
    x"3245B230",
    x"3245997B",
    x"324580C9",
    x"3245681B",
    x"32454F6F",
    x"324536C7",
    x"32451E22",
    x"3245057F",
    x"3244ECE0",
    x"3244D444",
    x"3244BBAB",
    x"3244A315",
    x"32448A82",
    x"324471F3",
    x"32445966",
    x"324440DC",
    x"32442856",
    x"32440FD2",
    x"3243F752",
    x"3243DED4",
    x"3243C65A",
    x"3243ADE3",
    x"3243956F",
    x"32437CFD",
    x"3243648F",
    x"32434C24",
    x"324333BC",
    x"32431B57",
    x"324302F5",
    x"3242EA97",
    x"3242D23B",
    x"3242B9E2",
    x"3242A18C",
    x"3242893A",
    x"324270EA",
    x"3242589D",
    x"32424054",
    x"3242280D",
    x"32420FCA",
    x"3241F789",
    x"3241DF4C",
    x"3241C712",
    x"3241AEDA",
    x"324196A6",
    x"32417E75",
    x"32416646",
    x"32414E1B",
    x"324135F3",
    x"32411DCD",
    x"324105AB",
    x"3240ED8C",
    x"3240D570",
    x"3240BD57",
    x"3240A541",
    x"32408D2D",
    x"3240751D",
    x"32405D10",
    x"32404506",
    x"32402CFF",
    x"324014FB",
    x"323FFCFA",
    x"323FE4FB",
    x"323FCD00",
    x"323FB508",
    x"323F9D13",
    x"323F8521",
    x"323F6D32",
    x"323F5546",
    x"323F3D5C",
    x"323F2576",
    x"323F0D93",
    x"323EF5B3",
    x"323EDDD6",
    x"323EC5FB",
    x"323EAE24",
    x"323E9650",
    x"323E7E7F",
    x"323E66B0",
    x"323E4EE5",
    x"323E371D",
    x"323E1F57",
    x"323E0795",
    x"323DEFD5",
    x"323DD819",
    x"323DC05F",
    x"323DA8A9",
    x"323D90F5",
    x"323D7944",
    x"323D6197",
    x"323D49EC",
    x"323D3244",
    x"323D1A9F",
    x"323D02FE",
    x"323CEB5F",
    x"323CD3C3",
    x"323CBC2A",
    x"323CA494",
    x"323C8D01",
    x"323C7571",
    x"323C5DE3",
    x"323C4659",
    x"323C2ED2",
    x"323C174D",
    x"323BFFCC",
    x"323BE84D",
    x"323BD0D2",
    x"323BB959",
    x"323BA1E3",
    x"323B8A71",
    x"323B7301",
    x"323B5B94",
    x"323B442A",
    x"323B2CC3",
    x"323B155F",
    x"323AFDFE",
    x"323AE69F",
    x"323ACF44",
    x"323AB7EB",
    x"323AA096",
    x"323A8943",
    x"323A71F4",
    x"323A5AA7",
    x"323A435D",
    x"323A2C16",
    x"323A14D2",
    x"3239FD91",
    x"3239E653",
    x"3239CF17",
    x"3239B7DF",
    x"3239A0A9",
    x"32398977",
    x"32397247",
    x"32395B1A",
    x"323943F0",
    x"32392CC9",
    x"323915A5",
    x"3238FE84",
    x"3238E765",
    x"3238D04A",
    x"3238B931",
    x"3238A21B",
    x"32388B09",
    x"323873F9",
    x"32385CEC",
    x"323845E1",
    x"32382EDA",
    x"323817D6",
    x"323800D4",
    x"3237E9D6",
    x"3237D2DA",
    x"3237BBE1",
    x"3237A4EB",
    x"32378DF8",
    x"32377707",
    x"3237601A",
    x"3237492F",
    x"32373248",
    x"32371B63",
    x"32370481",
    x"3236EDA2",
    x"3236D6C5",
    x"3236BFEC",
    x"3236A915",
    x"32369242",
    x"32367B71",
    x"323664A3",
    x"32364DD8",
    x"3236370F",
    x"3236204A",
    x"32360987",
    x"3235F2C7",
    x"3235DC0B",
    x"3235C550",
    x"3235AE99",
    x"323597E5",
    x"32358133",
    x"32356A85",
    x"323553D9",
    x"32353D30",
    x"32352689",
    x"32350FE6",
    x"3234F945",
    x"3234E2A8",
    x"3234CC0D",
    x"3234B575",
    x"32349EDF",
    x"3234884D",
    x"323471BD",
    x"32345B30",
    x"323444A6",
    x"32342E1F",
    x"3234179B",
    x"32340119",
    x"3233EA9B",
    x"3233D41F",
    x"3233BDA6",
    x"3233A72F",
    x"323390BC",
    x"32337A4B",
    x"323363DD",
    x"32334D72",
    x"3233370A",
    x"323320A4",
    x"32330A42",
    x"3232F3E2",
    x"3232DD85",
    x"3232C72A",
    x"3232B0D3",
    x"32329A7E",
    x"3232842C",
    x"32326DDD",
    x"32325791",
    x"32324147",
    x"32322B01",
    x"323214BD",
    x"3231FE7B",
    x"3231E83D",
    x"3231D201",
    x"3231BBC8",
    x"3231A592",
    x"32318F5F",
    x"3231792E",
    x"32316301",
    x"32314CD6",
    x"323136AE",
    x"32312088",
    x"32310A65",
    x"3230F445",
    x"3230DE28",
    x"3230C80E",
    x"3230B1F6",
    x"32309BE1",
    x"323085CF",
    x"32306FC0",
    x"323059B3",
    x"323043AA",
    x"32302DA2",
    x"3230179E",
    x"3230019D",
    x"322FEB9E",
    x"322FD5A2",
    x"322FBFA8",
    x"322FA9B2",
    x"322F93BE",
    x"322F7DCD",
    x"322F67DE",
    x"322F51F3",
    x"322F3C0A",
    x"322F2624",
    x"322F1040",
    x"322EFA60",
    x"322EE482",
    x"322ECEA7",
    x"322EB8CE",
    x"322EA2F8",
    x"322E8D25",
    x"322E7755",
    x"322E6188",
    x"322E4BBD",
    x"322E35F5",
    x"322E202F",
    x"322E0A6D",
    x"322DF4AD",
    x"322DDEEF",
    x"322DC935",
    x"322DB37D",
    x"322D9DC8",
    x"322D8816",
    x"322D7266",
    x"322D5CB9",
    x"322D470F",
    x"322D3167",
    x"322D1BC3",
    x"322D0620",
    x"322CF081",
    x"322CDAE4",
    x"322CC54A",
    x"322CAFB3",
    x"322C9A1E",
    x"322C848C",
    x"322C6EFD",
    x"322C5971",
    x"322C43E7",
    x"322C2E60",
    x"322C18DB",
    x"322C0359",
    x"322BEDDA",
    x"322BD85E",
    x"322BC2E4",
    x"322BAD6D",
    x"322B97F9",
    x"322B8287",
    x"322B6D18",
    x"322B57AC",
    x"322B4242",
    x"322B2CDB",
    x"322B1777",
    x"322B0216",
    x"322AECB7",
    x"322AD75A",
    x"322AC201",
    x"322AACAA",
    x"322A9756",
    x"322A8204",
    x"322A6CB5",
    x"322A5769",
    x"322A421F",
    x"322A2CD8",
    x"322A1794",
    x"322A0252",
    x"3229ED14",
    x"3229D7D7",
    x"3229C29E",
    x"3229AD67",
    x"32299832",
    x"32298301",
    x"32296DD1",
    x"322958A5",
    x"3229437B",
    x"32292E54",
    x"32291930",
    x"3229040E",
    x"3228EEEF",
    x"3228D9D2",
    x"3228C4B8",
    x"3228AFA1",
    x"32289A8C",
    x"3228857A",
    x"3228706B",
    x"32285B5E",
    x"32284654",
    x"3228314D",
    x"32281C48",
    x"32280746",
    x"3227F246",
    x"3227DD49",
    x"3227C84F",
    x"3227B357",
    x"32279E62",
    x"3227896F",
    x"3227747F",
    x"32275F92",
    x"32274AA8",
    x"322735C0",
    x"322720DA",
    x"32270BF7",
    x"3226F717",
    x"3226E23A",
    x"3226CD5F",
    x"3226B886",
    x"3226A3B0",
    x"32268EDD",
    x"32267A0D",
    x"3226653F",
    x"32265073",
    x"32263BAB",
    x"322626E5",
    x"32261221",
    x"3225FD60",
    x"3225E8A2",
    x"3225D3E6",
    x"3225BF2D",
    x"3225AA76",
    x"322595C2",
    x"32258111",
    x"32256C62",
    x"322557B5",
    x"3225430C",
    x"32252E65",
    x"322519C0",
    x"3225051E",
    x"3224F07F",
    x"3224DBE2",
    x"3224C748",
    x"3224B2B0",
    x"32249E1B",
    x"32248989",
    x"322474F9",
    x"3224606C",
    x"32244BE1",
    x"32243759",
    x"322422D3",
    x"32240E50",
    x"3223F9CF",
    x"3223E551",
    x"3223D0D6",
    x"3223BC5D",
    x"3223A7E7",
    x"32239373",
    x"32237F02",
    x"32236A94",
    x"32235627",
    x"322341BE",
    x"32232D57",
    x"322318F3",
    x"32230491",
    x"3222F031",
    x"3222DBD5",
    x"3222C77B",
    x"3222B323",
    x"32229ECE",
    x"32228A7B",
    x"3222762B",
    x"322261DE",
    x"32224D93",
    x"3222394A",
    x"32222504",
    x"322210C1",
    x"3221FC80",
    x"3221E842",
    x"3221D406",
    x"3221BFCD",
    x"3221AB96",
    x"32219762",
    x"32218330",
    x"32216F01",
    x"32215AD5",
    x"322146AA",
    x"32213283",
    x"32211E5E",
    x"32210A3B",
    x"3220F61B",
    x"3220E1FE",
    x"3220CDE3",
    x"3220B9CA",
    x"3220A5B4",
    x"322091A1",
    x"32207D90",
    x"32206981",
    x"32205576",
    x"3220416C",
    x"32202D65",
    x"32201961",
    x"3220055F",
    x"321FF15F",
    x"321FDD62",
    x"321FC968",
    x"321FB570",
    x"321FA17B",
    x"321F8D88",
    x"321F7997",
    x"321F65A9",
    x"321F51BE",
    x"321F3DD5",
    x"321F29EE",
    x"321F160A",
    x"321F0229",
    x"321EEE4A",
    x"321EDA6D",
    x"321EC693",
    x"321EB2BC",
    x"321E9EE7",
    x"321E8B14",
    x"321E7744",
    x"321E6376",
    x"321E4FAB",
    x"321E3BE2",
    x"321E281C",
    x"321E1458",
    x"321E0097",
    x"321DECD8",
    x"321DD91C",
    x"321DC562",
    x"321DB1AA",
    x"321D9DF5",
    x"321D8A43",
    x"321D7693",
    x"321D62E5",
    x"321D4F3A",
    x"321D3B91",
    x"321D27EB",
    x"321D1447",
    x"321D00A6",
    x"321CED07",
    x"321CD96B",
    x"321CC5D1",
    x"321CB239",
    x"321C9EA4",
    x"321C8B12",
    x"321C7782",
    x"321C63F4",
    x"321C5069",
    x"321C3CE0",
    x"321C2959",
    x"321C15D5",
    x"321C0254",
    x"321BEED5",
    x"321BDB58",
    x"321BC7DE",
    x"321BB466",
    x"321BA0F1",
    x"321B8D7E",
    x"321B7A0E",
    x"321B66A0",
    x"321B5334",
    x"321B3FCB",
    x"321B2C64",
    x"321B1900",
    x"321B059E",
    x"321AF23E",
    x"321ADEE1",
    x"321ACB86",
    x"321AB82E",
    x"321AA4D8",
    x"321A9185",
    x"321A7E34",
    x"321A6AE5",
    x"321A5799",
    x"321A4450",
    x"321A3108",
    x"321A1DC3",
    x"321A0A81",
    x"3219F741",
    x"3219E403",
    x"3219D0C8",
    x"3219BD8F",
    x"3219AA58",
    x"32199724",
    x"321983F3",
    x"321970C3",
    x"32195D96",
    x"32194A6C",
    x"32193744",
    x"3219241E",
    x"321910FB",
    x"3218FDDA",
    x"3218EABB",
    x"3218D79F",
    x"3218C485",
    x"3218B16E",
    x"32189E59",
    x"32188B46",
    x"32187836",
    x"32186528",
    x"3218521D",
    x"32183F14",
    x"32182C0D",
    x"32181909",
    x"32180607",
    x"3217F307",
    x"3217E00A",
    x"3217CD0F",
    x"3217BA17",
    x"3217A721",
    x"3217942D",
    x"3217813C",
    x"32176E4D",
    x"32175B60",
    x"32174876",
    x"3217358E",
    x"321722A8",
    x"32170FC5",
    x"3216FCE5",
    x"3216EA06",
    x"3216D72A",
    x"3216C450",
    x"3216B179",
    x"32169EA4",
    x"32168BD1",
    x"32167901",
    x"32166633",
    x"32165367",
    x"3216409E",
    x"32162DD7",
    x"32161B13",
    x"32160851",
    x"3215F591",
    x"3215E2D3",
    x"3215D018",
    x"3215BD5F",
    x"3215AAA9",
    x"321597F4",
    x"32158543",
    x"32157293",
    x"32155FE6",
    x"32154D3B",
    x"32153A93",
    x"321527ED",
    x"32151549",
    x"321502A7",
    x"3214F008",
    x"3214DD6B",
    x"3214CAD1",
    x"3214B838",
    x"3214A5A3",
    x"3214930F",
    x"3214807E",
    x"32146DEF",
    x"32145B62",
    x"321448D8",
    x"32143650",
    x"321423CB",
    x"32141147",
    x"3213FEC6",
    x"3213EC48",
    x"3213D9CB",
    x"3213C751",
    x"3213B4D9",
    x"3213A264",
    x"32138FF1",
    x"32137D80",
    x"32136B11",
    x"321358A5",
    x"3213463B",
    x"321333D4",
    x"3213216E",
    x"32130F0B",
    x"3212FCAA",
    x"3212EA4C",
    x"3212D7F0",
    x"3212C596",
    x"3212B33E",
    x"3212A0E9",
    x"32128E96",
    x"32127C46",
    x"321269F7",
    x"321257AB",
    x"32124561",
    x"3212331A",
    x"321220D4",
    x"32120E92",
    x"3211FC51",
    x"3211EA12",
    x"3211D7D6",
    x"3211C59C",
    x"3211B365",
    x"3211A130",
    x"32118EFD",
    x"32117CCC",
    x"32116A9D",
    x"32115871",
    x"32114647",
    x"32113420",
    x"321121FA",
    x"32110FD7",
    x"3210FDB6",
    x"3210EB98",
    x"3210D97B",
    x"3210C761",
    x"3210B54A",
    x"3210A334",
    x"32109121",
    x"32107F10",
    x"32106D01",
    x"32105AF5",
    x"321048EA",
    x"321036E2",
    x"321024DD",
    x"321012D9",
    x"321000D8",
    x"320FEED9",
    x"320FDCDC",
    x"320FCAE2",
    x"320FB8E9",
    x"320FA6F3",
    x"320F9500",
    x"320F830E",
    x"320F711F",
    x"320F5F32",
    x"320F4D47",
    x"320F3B5F",
    x"320F2978",
    x"320F1794",
    x"320F05B2",
    x"320EF3D3",
    x"320EE1F5",
    x"320ED01A",
    x"320EBE41",
    x"320EAC6B",
    x"320E9A96",
    x"320E88C4",
    x"320E76F4",
    x"320E6526",
    x"320E535B",
    x"320E4191",
    x"320E2FCA",
    x"320E1E06",
    x"320E0C43",
    x"320DFA82",
    x"320DE8C4",
    x"320DD708",
    x"320DC54F",
    x"320DB397",
    x"320DA1E2",
    x"320D902E",
    x"320D7E7E",
    x"320D6CCF",
    x"320D5B22",
    x"320D4978",
    x"320D37D0",
    x"320D262A",
    x"320D1486",
    x"320D02E5",
    x"320CF146",
    x"320CDFA9",
    x"320CCE0E",
    x"320CBC75",
    x"320CAADF",
    x"320C994A",
    x"320C87B8",
    x"320C7629",
    x"320C649B",
    x"320C530F",
    x"320C4186",
    x"320C2FFF",
    x"320C1E7A",
    x"320C0CF7",
    x"320BFB77",
    x"320BE9F8",
    x"320BD87C",
    x"320BC702",
    x"320BB58B",
    x"320BA415",
    x"320B92A2",
    x"320B8130",
    x"320B6FC1",
    x"320B5E54",
    x"320B4CEA",
    x"320B3B81",
    x"320B2A1B",
    x"320B18B7",
    x"320B0755",
    x"320AF5F5",
    x"320AE497",
    x"320AD33C",
    x"320AC1E2",
    x"320AB08B",
    x"320A9F36",
    x"320A8DE3",
    x"320A7C93",
    x"320A6B44",
    x"320A59F8",
    x"320A48AE",
    x"320A3766",
    x"320A2620",
    x"320A14DC",
    x"320A039B",
    x"3209F25B",
    x"3209E11E",
    x"3209CFE3",
    x"3209BEAA",
    x"3209AD73",
    x"32099C3F",
    x"32098B0C",
    x"320979DC",
    x"320968AE",
    x"32095782",
    x"32094658",
    x"32093530",
    x"3209240B",
    x"320912E7",
    x"320901C6",
    x"3208F0A7",
    x"3208DF8A",
    x"3208CE6F",
    x"3208BD56",
    x"3208AC40",
    x"32089B2B",
    x"32088A19",
    x"32087909",
    x"320867FB",
    x"320856EF",
    x"320845E5",
    x"320834DD",
    x"320823D8",
    x"320812D4",
    x"320801D3",
    x"3207F0D4",
    x"3207DFD7",
    x"3207CEDC",
    x"3207BDE3",
    x"3207ACEC",
    x"32079BF8",
    x"32078B05",
    x"32077A15",
    x"32076927",
    x"3207583B",
    x"32074751",
    x"32073669",
    x"32072583",
    x"3207149F",
    x"320703BE",
    x"3206F2DF",
    x"3206E201",
    x"3206D126",
    x"3206C04D",
    x"3206AF76",
    x"32069EA1",
    x"32068DCE",
    x"32067CFE",
    x"32066C2F",
    x"32065B63",
    x"32064A98",
    x"320639D0",
    x"3206290A",
    x"32061846",
    x"32060784",
    x"3205F6C4",
    x"3205E606",
    x"3205D54A",
    x"3205C491",
    x"3205B3D9",
    x"3205A324",
    x"32059270",
    x"320581BF",
    x"32057110",
    x"32056063",
    x"32054FB8",
    x"32053F0F",
    x"32052E68",
    x"32051DC3",
    x"32050D21",
    x"3204FC80",
    x"3204EBE1",
    x"3204DB45",
    x"3204CAAB",
    x"3204BA12",
    x"3204A97C",
    x"320498E8",
    x"32048856",
    x"320477C6",
    x"32046738",
    x"320456AC",
    x"32044622",
    x"3204359B",
    x"32042515",
    x"32041491",
    x"32040410",
    x"3203F390",
    x"3203E313",
    x"3203D298",
    x"3203C21E",
    x"3203B1A7",
    x"3203A132",
    x"320390BF",
    x"3203804E",
    x"32036FDF",
    x"32035F72",
    x"32034F07",
    x"32033E9E",
    x"32032E37",
    x"32031DD2",
    x"32030D70",
    x"3202FD0F",
    x"3202ECB0",
    x"3202DC54",
    x"3202CBF9",
    x"3202BBA1",
    x"3202AB4A",
    x"32029AF6",
    x"32028AA4",
    x"32027A53",
    x"32026A05",
    x"320259B9",
    x"3202496F",
    x"32023926",
    x"320228E0",
    x"3202189C",
    x"3202085A",
    x"3201F81A",
    x"3201E7DC",
    x"3201D7A0",
    x"3201C766",
    x"3201B72E",
    x"3201A6F8",
    x"320196C5",
    x"32018693",
    x"32017663",
    x"32016635",
    x"32015609",
    x"320145E0",
    x"320135B8",
    x"32012592",
    x"3201156F",
    x"3201054D",
    x"3200F52D",
    x"3200E510",
    x"3200D4F4",
    x"3200C4DA",
    x"3200B4C3",
    x"3200A4AD",
    x"3200949A",
    x"32008488",
    x"32007478",
    x"3200646B",
    x"3200545F",
    x"32004456",
    x"3200344E",
    x"32002449",
    x"32001445",
    x"32000444",
    x"31FFE888",
    x"31FFC88D",
    x"31FFA896",
    x"31FF88A3",
    x"31FF68B4",
    x"31FF48C9",
    x"31FF28E2",
    x"31FF08FF",
    x"31FEE91F",
    x"31FEC944",
    x"31FEA96D",
    x"31FE899A",
    x"31FE69CB",
    x"31FE4A00",
    x"31FE2A38",
    x"31FE0A75",
    x"31FDEAB6",
    x"31FDCAFA",
    x"31FDAB43",
    x"31FD8B8F",
    x"31FD6BE0",
    x"31FD4C34",
    x"31FD2C8D",
    x"31FD0CE9",
    x"31FCED4A",
    x"31FCCDAE",
    x"31FCAE16",
    x"31FC8E83",
    x"31FC6EF3",
    x"31FC4F67",
    x"31FC2FDF",
    x"31FC105B",
    x"31FBF0DB",
    x"31FBD15F",
    x"31FBB1E6",
    x"31FB9272",
    x"31FB7302",
    x"31FB5395",
    x"31FB342D",
    x"31FB14C8",
    x"31FAF568",
    x"31FAD60B",
    x"31FAB6B2",
    x"31FA975D",
    x"31FA780C",
    x"31FA58BF",
    x"31FA3976",
    x"31FA1A31",
    x"31F9FAF0",
    x"31F9DBB2",
    x"31F9BC79",
    x"31F99D43",
    x"31F97E11",
    x"31F95EE4",
    x"31F93FBA",
    x"31F92094",
    x"31F90171",
    x"31F8E253",
    x"31F8C339",
    x"31F8A422",
    x"31F88510",
    x"31F86601",
    x"31F846F6",
    x"31F827EF",
    x"31F808EC",
    x"31F7E9ED",
    x"31F7CAF2",
    x"31F7ABFA",
    x"31F78D07",
    x"31F76E17",
    x"31F74F2B",
    x"31F73043",
    x"31F7115F",
    x"31F6F27F",
    x"31F6D3A3",
    x"31F6B4CA",
    x"31F695F5",
    x"31F67725",
    x"31F65858",
    x"31F6398F",
    x"31F61AC9",
    x"31F5FC08",
    x"31F5DD4A",
    x"31F5BE91",
    x"31F59FDB",
    x"31F58129",
    x"31F5627A",
    x"31F543D0",
    x"31F52529",
    x"31F50687",
    x"31F4E7E8",
    x"31F4C94D",
    x"31F4AAB5",
    x"31F48C22",
    x"31F46D92",
    x"31F44F07",
    x"31F4307F",
    x"31F411FB",
    x"31F3F37A",
    x"31F3D4FE",
    x"31F3B685",
    x"31F39810",
    x"31F3799F",
    x"31F35B32",
    x"31F33CC8",
    x"31F31E62",
    x"31F30001",
    x"31F2E1A2",
    x"31F2C348",
    x"31F2A4F2",
    x"31F2869F",
    x"31F26850",
    x"31F24A05",
    x"31F22BBD",
    x"31F20D7A",
    x"31F1EF3A",
    x"31F1D0FE",
    x"31F1B2C6",
    x"31F19491",
    x"31F17661",
    x"31F15834",
    x"31F13A0B",
    x"31F11BE5",
    x"31F0FDC4",
    x"31F0DFA6",
    x"31F0C18C",
    x"31F0A375",
    x"31F08563",
    x"31F06754",
    x"31F04949",
    x"31F02B42",
    x"31F00D3E",
    x"31EFEF3E",
    x"31EFD142",
    x"31EFB34A",
    x"31EF9556",
    x"31EF7765",
    x"31EF5978",
    x"31EF3B8E",
    x"31EF1DA9",
    x"31EEFFC7",
    x"31EEE1E9",
    x"31EEC40F",
    x"31EEA638",
    x"31EE8865",
    x"31EE6A96",
    x"31EE4CCA",
    x"31EE2F03",
    x"31EE113F",
    x"31EDF37E",
    x"31EDD5C2",
    x"31EDB809",
    x"31ED9A54",
    x"31ED7CA2",
    x"31ED5EF5",
    x"31ED414B",
    x"31ED23A4",
    x"31ED0602",
    x"31ECE863",
    x"31ECCAC8",
    x"31ECAD30",
    x"31EC8F9C",
    x"31EC720C",
    x"31EC5480",
    x"31EC36F7",
    x"31EC1972",
    x"31EBFBF1",
    x"31EBDE73",
    x"31EBC0F9",
    x"31EBA383",
    x"31EB8610",
    x"31EB68A1",
    x"31EB4B36",
    x"31EB2DCE",
    x"31EB106B",
    x"31EAF30A",
    x"31EAD5AE",
    x"31EAB855",
    x"31EA9B00",
    x"31EA7DAE",
    x"31EA6060",
    x"31EA4316",
    x"31EA25CF",
    x"31EA088D",
    x"31E9EB4D",
    x"31E9CE12",
    x"31E9B0DA",
    x"31E993A6",
    x"31E97675",
    x"31E95948",
    x"31E93C1F",
    x"31E91EF9",
    x"31E901D7",
    x"31E8E4B8",
    x"31E8C79E",
    x"31E8AA87",
    x"31E88D73",
    x"31E87063",
    x"31E85357",
    x"31E8364E",
    x"31E81949",
    x"31E7FC48",
    x"31E7DF4A",
    x"31E7C250",
    x"31E7A55A",
    x"31E78867",
    x"31E76B78",
    x"31E74E8C",
    x"31E731A4",
    x"31E714C0",
    x"31E6F7DF",
    x"31E6DB02",
    x"31E6BE28",
    x"31E6A152",
    x"31E68480",
    x"31E667B1",
    x"31E64AE6",
    x"31E62E1E",
    x"31E6115A",
    x"31E5F49A",
    x"31E5D7DD",
    x"31E5BB24",
    x"31E59E6E",
    x"31E581BC",
    x"31E5650E",
    x"31E54863",
    x"31E52BBC",
    x"31E50F18",
    x"31E4F278",
    x"31E4D5DB",
    x"31E4B943",
    x"31E49CAD",
    x"31E4801B",
    x"31E4638D",
    x"31E44702",
    x"31E42A7B",
    x"31E40DF8",
    x"31E3F178",
    x"31E3D4FB",
    x"31E3B883",
    x"31E39C0D",
    x"31E37F9C",
    x"31E3632D",
    x"31E346C3",
    x"31E32A5C",
    x"31E30DF8",
    x"31E2F198",
    x"31E2D53C",
    x"31E2B8E3",
    x"31E29C8E",
    x"31E2803C",
    x"31E263EE",
    x"31E247A3",
    x"31E22B5C",
    x"31E20F18",
    x"31E1F2D8",
    x"31E1D69B",
    x"31E1BA62",
    x"31E19E2D",
    x"31E181FB",
    x"31E165CC",
    x"31E149A1",
    x"31E12D7A",
    x"31E11156",
    x"31E0F535",
    x"31E0D919",
    x"31E0BCFF",
    x"31E0A0E9",
    x"31E084D7",
    x"31E068C8",
    x"31E04CBD",
    x"31E030B5",
    x"31E014B1",
    x"31DFF8B0",
    x"31DFDCB2",
    x"31DFC0B9",
    x"31DFA4C2",
    x"31DF88CF",
    x"31DF6CE0",
    x"31DF50F4",
    x"31DF350C",
    x"31DF1927",
    x"31DEFD46",
    x"31DEE168",
    x"31DEC58D",
    x"31DEA9B6",
    x"31DE8DE3",
    x"31DE7213",
    x"31DE5646",
    x"31DE3A7D",
    x"31DE1EB8",
    x"31DE02F5",
    x"31DDE737",
    x"31DDCB7C",
    x"31DDAFC4",
    x"31DD9410",
    x"31DD785F",
    x"31DD5CB2",
    x"31DD4108",
    x"31DD2561",
    x"31DD09BE",
    x"31DCEE1F",
    x"31DCD283",
    x"31DCB6EA",
    x"31DC9B55",
    x"31DC7FC3",
    x"31DC6435",
    x"31DC48AA",
    x"31DC2D23",
    x"31DC119F",
    x"31DBF61F",
    x"31DBDAA2",
    x"31DBBF28",
    x"31DBA3B2",
    x"31DB883F",
    x"31DB6CD0",
    x"31DB5164",
    x"31DB35FB",
    x"31DB1A96",
    x"31DAFF35",
    x"31DAE3D7",
    x"31DAC87C",
    x"31DAAD24",
    x"31DA91D1",
    x"31DA7680",
    x"31DA5B33",
    x"31DA3FE9",
    x"31DA24A3",
    x"31DA0960",
    x"31D9EE21",
    x"31D9D2E5",
    x"31D9B7AC",
    x"31D99C77",
    x"31D98145",
    x"31D96616",
    x"31D94AEB",
    x"31D92FC4",
    x"31D9149F",
    x"31D8F97E",
    x"31D8DE61",
    x"31D8C347",
    x"31D8A830",
    x"31D88D1D",
    x"31D8720D",
    x"31D85700",
    x"31D83BF7",
    x"31D820F1",
    x"31D805EF",
    x"31D7EAF0",
    x"31D7CFF4",
    x"31D7B4FC",
    x"31D79A07",
    x"31D77F15",
    x"31D76427",
    x"31D7493C",
    x"31D72E55",
    x"31D71371",
    x"31D6F890",
    x"31D6DDB2",
    x"31D6C2D8",
    x"31D6A802",
    x"31D68D2E",
    x"31D6725E",
    x"31D65792",
    x"31D63CC9",
    x"31D62203",
    x"31D60740",
    x"31D5EC81",
    x"31D5D1C5",
    x"31D5B70C",
    x"31D59C57",
    x"31D581A5",
    x"31D566F7",
    x"31D54C4C",
    x"31D531A4",
    x"31D516FF",
    x"31D4FC5E",
    x"31D4E1C0",
    x"31D4C726",
    x"31D4AC8E",
    x"31D491FA",
    x"31D4776A",
    x"31D45CDD",
    x"31D44253",
    x"31D427CC",
    x"31D40D49",
    x"31D3F2C9",
    x"31D3D84C",
    x"31D3BDD3",
    x"31D3A35C",
    x"31D388EA",
    x"31D36E7A",
    x"31D3540E",
    x"31D339A5",
    x"31D31F40",
    x"31D304DD",
    x"31D2EA7E",
    x"31D2D023",
    x"31D2B5CA",
    x"31D29B75",
    x"31D28124",
    x"31D266D5",
    x"31D24C8A",
    x"31D23242",
    x"31D217FD",
    x"31D1FDBC",
    x"31D1E37E",
    x"31D1C943",
    x"31D1AF0C",
    x"31D194D7",
    x"31D17AA6",
    x"31D16079",
    x"31D1464E",
    x"31D12C27",
    x"31D11203",
    x"31D0F7E3",
    x"31D0DDC5",
    x"31D0C3AB",
    x"31D0A994",
    x"31D08F81",
    x"31D07570",
    x"31D05B63",
    x"31D0415A",
    x"31D02753",
    x"31D00D50",
    x"31CFF350",
    x"31CFD953",
    x"31CFBF59",
    x"31CFA563",
    x"31CF8B70",
    x"31CF7180",
    x"31CF5794",
    x"31CF3DAA",
    x"31CF23C4",
    x"31CF09E1",
    x"31CEF002",
    x"31CED625",
    x"31CEBC4C",
    x"31CEA276",
    x"31CE88A4",
    x"31CE6ED4",
    x"31CE5508",
    x"31CE3B3F",
    x"31CE2179",
    x"31CE07B7",
    x"31CDEDF7",
    x"31CDD43B",
    x"31CDBA82",
    x"31CDA0CC",
    x"31CD871A",
    x"31CD6D6B",
    x"31CD53BF",
    x"31CD3A16",
    x"31CD2070",
    x"31CD06CE",
    x"31CCED2E",
    x"31CCD392",
    x"31CCB9F9",
    x"31CCA064",
    x"31CC86D1",
    x"31CC6D42",
    x"31CC53B6",
    x"31CC3A2D",
    x"31CC20A7",
    x"31CC0725",
    x"31CBEDA6",
    x"31CBD42A",
    x"31CBBAB1",
    x"31CBA13B",
    x"31CB87C8",
    x"31CB6E59",
    x"31CB54ED",
    x"31CB3B84",
    x"31CB221E",
    x"31CB08BB",
    x"31CAEF5C",
    x"31CAD5FF",
    x"31CABCA6",
    x"31CAA350",
    x"31CA89FD",
    x"31CA70AE",
    x"31CA5761",
    x"31CA3E18",
    x"31CA24D2",
    x"31CA0B8F",
    x"31C9F24F",
    x"31C9D912",
    x"31C9BFD8",
    x"31C9A6A2",
    x"31C98D6F",
    x"31C9743F",
    x"31C95B12",
    x"31C941E8",
    x"31C928C1",
    x"31C90F9E",
    x"31C8F67D",
    x"31C8DD60",
    x"31C8C446",
    x"31C8AB2F",
    x"31C8921B",
    x"31C8790B",
    x"31C85FFD",
    x"31C846F3",
    x"31C82DEB",
    x"31C814E7",
    x"31C7FBE6",
    x"31C7E2E8",
    x"31C7C9ED",
    x"31C7B0F6",
    x"31C79801",
    x"31C77F10",
    x"31C76621",
    x"31C74D36",
    x"31C7344E",
    x"31C71B69",
    x"31C70287",
    x"31C6E9A8",
    x"31C6D0CD",
    x"31C6B7F4",
    x"31C69F1F",
    x"31C6864C",
    x"31C66D7D",
    x"31C654B1",
    x"31C63BE8",
    x"31C62322",
    x"31C60A5F",
    x"31C5F19F",
    x"31C5D8E3",
    x"31C5C029",
    x"31C5A773",
    x"31C58EBF",
    x"31C5760F",
    x"31C55D62",
    x"31C544B8",
    x"31C52C11",
    x"31C5136D",
    x"31C4FACC",
    x"31C4E22E",
    x"31C4C993",
    x"31C4B0FC",
    x"31C49867",
    x"31C47FD6",
    x"31C46747",
    x"31C44EBC",
    x"31C43633",
    x"31C41DAE",
    x"31C4052C",
    x"31C3ECAD",
    x"31C3D431",
    x"31C3BBB8",
    x"31C3A342",
    x"31C38ACF",
    x"31C3725F",
    x"31C359F2",
    x"31C34189",
    x"31C32922",
    x"31C310BE",
    x"31C2F85E",
    x"31C2E000",
    x"31C2C7A6",
    x"31C2AF4E",
    x"31C296FA",
    x"31C27EA9",
    x"31C2665A",
    x"31C24E0F",
    x"31C235C7",
    x"31C21D82",
    x"31C2053F",
    x"31C1ED00",
    x"31C1D4C4",
    x"31C1BC8B",
    x"31C1A455",
    x"31C18C22",
    x"31C173F2",
    x"31C15BC5",
    x"31C1439B",
    x"31C12B74",
    x"31C11350",
    x"31C0FB2F",
    x"31C0E311",
    x"31C0CAF7",
    x"31C0B2DF",
    x"31C09ACA",
    x"31C082B8",
    x"31C06AA9",
    x"31C0529D",
    x"31C03A94",
    x"31C0228F",
    x"31C00A8C",
    x"31BFF28C",
    x"31BFDA8F",
    x"31BFC295",
    x"31BFAA9F",
    x"31BF92AB",
    x"31BF7ABA",
    x"31BF62CC",
    x"31BF4AE1",
    x"31BF32F9",
    x"31BF1B14",
    x"31BF0333",
    x"31BEEB54",
    x"31BED378",
    x"31BEBB9F",
    x"31BEA3C9",
    x"31BE8BF6",
    x"31BE7426",
    x"31BE5C59",
    x"31BE448F",
    x"31BE2CC8",
    x"31BE1504",
    x"31BDFD42",
    x"31BDE584",
    x"31BDCDC9",
    x"31BDB611",
    x"31BD9E5C",
    x"31BD86A9",
    x"31BD6EFA",
    x"31BD574D",
    x"31BD3FA4",
    x"31BD27FE",
    x"31BD105A",
    x"31BCF8B9",
    x"31BCE11C",
    x"31BCC981",
    x"31BCB1E9",
    x"31BC9A55",
    x"31BC82C3",
    x"31BC6B34",
    x"31BC53A8",
    x"31BC3C1F",
    x"31BC2499",
    x"31BC0D16",
    x"31BBF596",
    x"31BBDE19",
    x"31BBC69E",
    x"31BBAF27",
    x"31BB97B2",
    x"31BB8041",
    x"31BB68D2",
    x"31BB5167",
    x"31BB39FE",
    x"31BB2298",
    x"31BB0B35",
    x"31BAF3D5",
    x"31BADC78",
    x"31BAC51E",
    x"31BAADC7",
    x"31BA9673",
    x"31BA7F22",
    x"31BA67D3",
    x"31BA5088",
    x"31BA393F",
    x"31BA21F9",
    x"31BA0AB6",
    x"31B9F377",
    x"31B9DC3A",
    x"31B9C500",
    x"31B9ADC8",
    x"31B99694",
    x"31B97F63",
    x"31B96834",
    x"31B95109",
    x"31B939E0",
    x"31B922BA",
    x"31B90B97",
    x"31B8F477",
    x"31B8DD5A",
    x"31B8C640",
    x"31B8AF29",
    x"31B89814",
    x"31B88103",
    x"31B869F4",
    x"31B852E8",
    x"31B83BDF",
    x"31B824D9",
    x"31B80DD6",
    x"31B7F6D6",
    x"31B7DFD8",
    x"31B7C8DE",
    x"31B7B1E6",
    x"31B79AF1",
    x"31B783FF",
    x"31B76D10",
    x"31B75624",
    x"31B73F3B",
    x"31B72854",
    x"31B71171",
    x"31B6FA90",
    x"31B6E3B2",
    x"31B6CCD7",
    x"31B6B5FF",
    x"31B69F29",
    x"31B68857",
    x"31B67187",
    x"31B65ABB",
    x"31B643F1",
    x"31B62D2A",
    x"31B61665",
    x"31B5FFA4",
    x"31B5E8E5",
    x"31B5D22A",
    x"31B5BB71",
    x"31B5A4BB",
    x"31B58E08",
    x"31B57757",
    x"31B560AA",
    x"31B549FF",
    x"31B53357",
    x"31B51CB2",
    x"31B50610",
    x"31B4EF71",
    x"31B4D8D4",
    x"31B4C23B",
    x"31B4ABA4",
    x"31B49510",
    x"31B47E7F",
    x"31B467F0",
    x"31B45165",
    x"31B43ADC",
    x"31B42456",
    x"31B40DD3",
    x"31B3F752",
    x"31B3E0D5",
    x"31B3CA5A",
    x"31B3B3E2",
    x"31B39D6D",
    x"31B386FB",
    x"31B3708B",
    x"31B35A1F",
    x"31B343B5",
    x"31B32D4E",
    x"31B316EA",
    x"31B30088",
    x"31B2EA29",
    x"31B2D3CE",
    x"31B2BD75",
    x"31B2A71E",
    x"31B290CB",
    x"31B27A7A",
    x"31B2642C",
    x"31B24DE1",
    x"31B23799",
    x"31B22153",
    x"31B20B10",
    x"31B1F4D0",
    x"31B1DE93",
    x"31B1C859",
    x"31B1B221",
    x"31B19BEC",
    x"31B185BA",
    x"31B16F8B",
    x"31B1595E",
    x"31B14334",
    x"31B12D0D",
    x"31B116E9",
    x"31B100C8",
    x"31B0EAA9",
    x"31B0D48D",
    x"31B0BE74",
    x"31B0A85D",
    x"31B0924A",
    x"31B07C39",
    x"31B0662B",
    x"31B0501F",
    x"31B03A17",
    x"31B02411",
    x"31B00E0E",
    x"31AFF80D",
    x"31AFE210",
    x"31AFCC15",
    x"31AFB61D",
    x"31AFA027",
    x"31AF8A35",
    x"31AF7445",
    x"31AF5E57",
    x"31AF486D",
    x"31AF3285",
    x"31AF1CA0",
    x"31AF06BE",
    x"31AEF0DF",
    x"31AEDB02",
    x"31AEC528",
    x"31AEAF51",
    x"31AE997C",
    x"31AE83AA",
    x"31AE6DDB",
    x"31AE580F",
    x"31AE4245",
    x"31AE2C7E",
    x"31AE16BA",
    x"31AE00F9",
    x"31ADEB3A",
    x"31ADD57E",
    x"31ADBFC4",
    x"31ADAA0E",
    x"31AD945A",
    x"31AD7EA9",
    x"31AD68FA",
    x"31AD534F",
    x"31AD3DA5",
    x"31AD27FF",
    x"31AD125B",
    x"31ACFCBB",
    x"31ACE71C",
    x"31ACD181",
    x"31ACBBE8",
    x"31ACA652",
    x"31AC90BE",
    x"31AC7B2E",
    x"31AC65A0",
    x"31AC5014",
    x"31AC3A8C",
    x"31AC2506",
    x"31AC0F82",
    x"31ABFA02",
    x"31ABE484",
    x"31ABCF09",
    x"31ABB990",
    x"31ABA41A",
    x"31AB8EA7",
    x"31AB7936",
    x"31AB63C9",
    x"31AB4E5E",
    x"31AB38F5",
    x"31AB238F",
    x"31AB0E2C",
    x"31AAF8CC",
    x"31AAE36E",
    x"31AACE13",
    x"31AAB8BA",
    x"31AAA365",
    x"31AA8E12",
    x"31AA78C1",
    x"31AA6373",
    x"31AA4E28",
    x"31AA38E0",
    x"31AA239A",
    x"31AA0E57",
    x"31A9F917",
    x"31A9E3D9",
    x"31A9CE9E",
    x"31A9B965",
    x"31A9A42F",
    x"31A98EFC",
    x"31A979CB",
    x"31A9649E",
    x"31A94F72",
    x"31A93A4A",
    x"31A92524",
    x"31A91000",
    x"31A8FAE0",
    x"31A8E5C2",
    x"31A8D0A6",
    x"31A8BB8E",
    x"31A8A677",
    x"31A89164",
    x"31A87C53",
    x"31A86745",
    x"31A85239",
    x"31A83D30",
    x"31A8282A",
    x"31A81326",
    x"31A7FE25",
    x"31A7E927",
    x"31A7D42B",
    x"31A7BF32",
    x"31A7AA3B",
    x"31A79547",
    x"31A78056",
    x"31A76B67",
    x"31A7567B",
    x"31A74191",
    x"31A72CAB",
    x"31A717C6",
    x"31A702E5",
    x"31A6EE06",
    x"31A6D929",
    x"31A6C44F",
    x"31A6AF78",
    x"31A69AA3",
    x"31A685D1",
    x"31A67102",
    x"31A65C35",
    x"31A6476B",
    x"31A632A3",
    x"31A61DDE",
    x"31A6091C",
    x"31A5F45C",
    x"31A5DF9F",
    x"31A5CAE4",
    x"31A5B62C",
    x"31A5A176",
    x"31A58CC4",
    x"31A57813",
    x"31A56366",
    x"31A54EBA",
    x"31A53A12",
    x"31A5256C",
    x"31A510C9",
    x"31A4FC28",
    x"31A4E789",
    x"31A4D2EE",
    x"31A4BE55",
    x"31A4A9BE",
    x"31A4952A",
    x"31A48099",
    x"31A46C0A",
    x"31A4577E",
    x"31A442F4",
    x"31A42E6D",
    x"31A419E9",
    x"31A40567",
    x"31A3F0E7",
    x"31A3DC6A",
    x"31A3C7F0",
    x"31A3B379",
    x"31A39F03",
    x"31A38A91",
    x"31A37621",
    x"31A361B3",
    x"31A34D48",
    x"31A338E0",
    x"31A3247A",
    x"31A31017",
    x"31A2FBB6",
    x"31A2E758",
    x"31A2D2FC",
    x"31A2BEA3",
    x"31A2AA4D",
    x"31A295F9",
    x"31A281A7",
    x"31A26D58",
    x"31A2590C",
    x"31A244C2",
    x"31A2307B",
    x"31A21C36",
    x"31A207F3",
    x"31A1F3B4",
    x"31A1DF77",
    x"31A1CB3C",
    x"31A1B704",
    x"31A1A2CE",
    x"31A18E9B",
    x"31A17A6A",
    x"31A1663C",
    x"31A15211",
    x"31A13DE8",
    x"31A129C1",
    x"31A1159D",
    x"31A1017C",
    x"31A0ED5D",
    x"31A0D941",
    x"31A0C527",
    x"31A0B10F",
    x"31A09CFB",
    x"31A088E8",
    x"31A074D8",
    x"31A060CB",
    x"31A04CC0",
    x"31A038B8",
    x"31A024B2",
    x"31A010AF",
    x"319FFCAE",
    x"319FE8AF",
    x"319FD4B4",
    x"319FC0BA",
    x"319FACC3",
    x"319F98CF",
    x"319F84DD",
    x"319F70EE",
    x"319F5D01",
    x"319F4917",
    x"319F352F",
    x"319F2149",
    x"319F0D66",
    x"319EF986",
    x"319EE5A8",
    x"319ED1CD",
    x"319EBDF4",
    x"319EAA1D",
    x"319E9649",
    x"319E8277",
    x"319E6EA8",
    x"319E5ADC",
    x"319E4712",
    x"319E334A",
    x"319E1F85",
    x"319E0BC2",
    x"319DF802",
    x"319DE444",
    x"319DD089",
    x"319DBCD0",
    x"319DA91A",
    x"319D9566",
    x"319D81B4",
    x"319D6E05",
    x"319D5A59",
    x"319D46AF",
    x"319D3307",
    x"319D1F62",
    x"319D0BBF",
    x"319CF81F",
    x"319CE481",
    x"319CD0E6",
    x"319CBD4D",
    x"319CA9B7",
    x"319C9623",
    x"319C8291",
    x"319C6F02",
    x"319C5B75",
    x"319C47EB",
    x"319C3463",
    x"319C20DE",
    x"319C0D5B",
    x"319BF9DB",
    x"319BE65D",
    x"319BD2E1",
    x"319BBF68",
    x"319BABF1",
    x"319B987D",
    x"319B850B",
    x"319B719C",
    x"319B5E2F",
    x"319B4AC4",
    x"319B375C",
    x"319B23F6",
    x"319B1093",
    x"319AFD32",
    x"319AE9D4",
    x"319AD678",
    x"319AC31E",
    x"319AAFC7",
    x"319A9C72",
    x"319A8920",
    x"319A75D0",
    x"319A6282",
    x"319A4F37",
    x"319A3BEF",
    x"319A28A8",
    x"319A1564",
    x"319A0223",
    x"3199EEE4",
    x"3199DBA7",
    x"3199C86D",
    x"3199B535",
    x"3199A200",
    x"31998ECD",
    x"31997B9C",
    x"3199686E",
    x"31995542",
    x"31994218",
    x"31992EF1",
    x"31991BCD",
    x"319908AA",
    x"3198F58A",
    x"3198E26D",
    x"3198CF52",
    x"3198BC39",
    x"3198A923",
    x"3198960F",
    x"319882FD",
    x"31986FEE",
    x"31985CE1",
    x"319849D7",
    x"319836CF",
    x"319823C9",
    x"319810C6",
    x"3197FDC5",
    x"3197EAC6",
    x"3197D7CA",
    x"3197C4D0",
    x"3197B1D9",
    x"31979EE4",
    x"31978BF1",
    x"31977901",
    x"31976613",
    x"31975328",
    x"3197403E",
    x"31972D57",
    x"31971A73",
    x"31970791",
    x"3196F4B1",
    x"3196E1D4",
    x"3196CEF9",
    x"3196BC20",
    x"3196A94A",
    x"31969676",
    x"319683A4",
    x"319670D5",
    x"31965E08",
    x"31964B3D",
    x"31963875",
    x"319625AF",
    x"319612EC",
    x"3196002A",
    x"3195ED6B",
    x"3195DAAF",
    x"3195C7F5",
    x"3195B53D",
    x"3195A288",
    x"31958FD4",
    x"31957D24",
    x"31956A75",
    x"319557C9",
    x"3195451F",
    x"31953278",
    x"31951FD3",
    x"31950D30",
    x"3194FA8F",
    x"3194E7F1",
    x"3194D555",
    x"3194C2BC",
    x"3194B025",
    x"31949D90",
    x"31948AFD",
    x"3194786D",
    x"319465DF",
    x"31945353",
    x"319440CA",
    x"31942E43",
    x"31941BBF",
    x"3194093C",
    x"3193F6BC",
    x"3193E43F",
    x"3193D1C3",
    x"3193BF4A",
    x"3193ACD3",
    x"31939A5F",
    x"319387ED",
    x"3193757D",
    x"3193630F",
    x"319350A4",
    x"31933E3B",
    x"31932BD5",
    x"31931970",
    x"3193070E",
    x"3192F4AF",
    x"3192E251",
    x"3192CFF6",
    x"3192BD9D",
    x"3192AB47",
    x"319298F2",
    x"319286A0",
    x"31927451",
    x"31926203",
    x"31924FB8",
    x"31923D6F",
    x"31922B29",
    x"319218E5",
    x"319206A3",
    x"3191F463",
    x"3191E226",
    x"3191CFEA",
    x"3191BDB2",
    x"3191AB7B",
    x"31919947",
    x"31918715",
    x"319174E5",
    x"319162B7",
    x"3191508C",
    x"31913E63",
    x"31912C3D",
    x"31911A18",
    x"319107F6",
    x"3190F5D6",
    x"3190E3B9",
    x"3190D19D",
    x"3190BF84",
    x"3190AD6D",
    x"31909B59",
    x"31908947",
    x"31907737",
    x"31906529",
    x"3190531D",
    x"31904114",
    x"31902F0D",
    x"31901D08",
    x"31900B06",
    x"318FF905",
    x"318FE707",
    x"318FD50C",
    x"318FC312",
    x"318FB11B",
    x"318F9F26",
    x"318F8D33",
    x"318F7B43",
    x"318F6954",
    x"318F5768",
    x"318F457F",
    x"318F3397",
    x"318F21B2",
    x"318F0FCF",
    x"318EFDEE",
    x"318EEC0F",
    x"318EDA33",
    x"318EC858",
    x"318EB681",
    x"318EA4AB",
    x"318E92D7",
    x"318E8106",
    x"318E6F37",
    x"318E5D6A",
    x"318E4BA0",
    x"318E39D7",
    x"318E2811",
    x"318E164D",
    x"318E048C",
    x"318DF2CC",
    x"318DE10F",
    x"318DCF54",
    x"318DBD9B",
    x"318DABE5",
    x"318D9A30",
    x"318D887E",
    x"318D76CE",
    x"318D6520",
    x"318D5375",
    x"318D41CB",
    x"318D3024",
    x"318D1E7F",
    x"318D0CDD",
    x"318CFB3C",
    x"318CE99E",
    x"318CD802",
    x"318CC668",
    x"318CB4D0",
    x"318CA33B",
    x"318C91A7",
    x"318C8016",
    x"318C6E87",
    x"318C5CFB",
    x"318C4B70",
    x"318C39E8",
    x"318C2862",
    x"318C16DE",
    x"318C055C",
    x"318BF3DC",
    x"318BE25F",
    x"318BD0E4",
    x"318BBF6B",
    x"318BADF4",
    x"318B9C7F",
    x"318B8B0D",
    x"318B799D",
    x"318B682E",
    x"318B56C2",
    x"318B4559",
    x"318B33F1",
    x"318B228C",
    x"318B1129",
    x"318AFFC7",
    x"318AEE69",
    x"318ADD0C",
    x"318ACBB1",
    x"318ABA59",
    x"318AA903",
    x"318A97AF",
    x"318A865D",
    x"318A750D",
    x"318A63C0",
    x"318A5274",
    x"318A412B",
    x"318A2FE4",
    x"318A1E9F",
    x"318A0D5C",
    x"3189FC1C",
    x"3189EADD",
    x"3189D9A1",
    x"3189C867",
    x"3189B72F",
    x"3189A5F9",
    x"318994C5",
    x"31898394",
    x"31897264",
    x"31896137",
    x"3189500C",
    x"31893EE3",
    x"31892DBC",
    x"31891C98",
    x"31890B75",
    x"3188FA55",
    x"3188E937",
    x"3188D81B",
    x"3188C701",
    x"3188B5E9",
    x"3188A4D3",
    x"318893C0",
    x"318882AE",
    x"3188719F",
    x"31886092",
    x"31884F87",
    x"31883E7E",
    x"31882D77",
    x"31881C73",
    x"31880B70",
    x"3187FA70",
    x"3187E971",
    x"3187D875",
    x"3187C77B",
    x"3187B683",
    x"3187A58E",
    x"3187949A",
    x"318783A9",
    x"318772B9",
    x"318761CC",
    x"318750E1",
    x"31873FF8",
    x"31872F11",
    x"31871E2C",
    x"31870D49",
    x"3186FC69",
    x"3186EB8A",
    x"3186DAAE",
    x"3186C9D3",
    x"3186B8FB",
    x"3186A825",
    x"31869751",
    x"3186867F",
    x"318675B0",
    x"318664E2",
    x"31865416",
    x"3186434D",
    x"31863286",
    x"318621C0",
    x"318610FD",
    x"3186003C",
    x"3185EF7D",
    x"3185DEC0",
    x"3185CE05",
    x"3185BD4D",
    x"3185AC96",
    x"31859BE1",
    x"31858B2F",
    x"31857A7F",
    x"318569D0",
    x"31855924",
    x"3185487A",
    x"318537D2",
    x"3185272C",
    x"31851688",
    x"318505E7",
    x"3184F547",
    x"3184E4A9",
    x"3184D40E",
    x"3184C374",
    x"3184B2DD",
    x"3184A247",
    x"318491B4",
    x"31848123",
    x"31847094",
    x"31846007",
    x"31844F7C",
    x"31843EF3",
    x"31842E6C",
    x"31841DE7",
    x"31840D65",
    x"3183FCE4",
    x"3183EC66",
    x"3183DBE9",
    x"3183CB6F",
    x"3183BAF6",
    x"3183AA80",
    x"31839A0C",
    x"31838999",
    x"31837929",
    x"318368BB",
    x"3183584F",
    x"318347E5",
    x"3183377D",
    x"31832717",
    x"318316B3",
    x"31830651",
    x"3182F5F2",
    x"3182E594",
    x"3182D538",
    x"3182C4DF",
    x"3182B487",
    x"3182A431",
    x"318293DE",
    x"3182838C",
    x"3182733D",
    x"318262F0",
    x"318252A4",
    x"3182425B",
    x"31823214",
    x"318221CE",
    x"3182118B",
    x"3182014A",
    x"3181F10B",
    x"3181E0CE",
    x"3181D093",
    x"3181C05A",
    x"3181B023",
    x"31819FEE",
    x"31818FBB",
    x"31817F8A",
    x"31816F5B",
    x"31815F2E",
    x"31814F03",
    x"31813EDA",
    x"31812EB3",
    x"31811E8E",
    x"31810E6C",
    x"3180FE4B",
    x"3180EE2C",
    x"3180DE0F",
    x"3180CDF5",
    x"3180BDDC",
    x"3180ADC5",
    x"31809DB0",
    x"31808D9E",
    x"31807D8D",
    x"31806D7E",
    x"31805D72",
    x"31804D67",
    x"31803D5E",
    x"31802D58",
    x"31801D53",
    x"31800D50",
    x"317FFA9F",
    x"317FDAA2",
    x"317FBAA9",
    x"317F9AB3",
    x"317F7AC2",
    x"317F5AD4",
    x"317F3AEB",
    x"317F1B06",
    x"317EFB24",
    x"317EDB47",
    x"317EBB6E",
    x"317E9B98",
    x"317E7BC7",
    x"317E5BF9",
    x"317E3C30",
    x"317E1C6A",
    x"317DFCA9",
    x"317DDCEB",
    x"317DBD31",
    x"317D9D7C",
    x"317D7DCA",
    x"317D5E1C",
    x"317D3E72",
    x"317D1ECD",
    x"317CFF2B",
    x"317CDF8D",
    x"317CBFF3",
    x"317CA05D",
    x"317C80CB",
    x"317C613D",
    x"317C41B2",
    x"317C222C",
    x"317C02AA",
    x"317BE32C",
    x"317BC3B1",
    x"317BA43B",
    x"317B84C8",
    x"317B6559",
    x"317B45EF",
    x"317B2688",
    x"317B0725",
    x"317AE7C6",
    x"317AC86B",
    x"317AA914",
    x"317A89C1",
    x"317A6A72",
    x"317A4B26",
    x"317A2BDF",
    x"317A0C9B",
    x"3179ED5C",
    x"3179CE20",
    x"3179AEE8",
    x"31798FB4",
    x"31797084",
    x"31795158",
    x"31793230",
    x"3179130C",
    x"3178F3EB",
    x"3178D4CF",
    x"3178B5B6",
    x"317896A1",
    x"31787790",
    x"31785883",
    x"3178397A",
    x"31781A75",
    x"3177FB73",
    x"3177DC76",
    x"3177BD7C",
    x"31779E87",
    x"31777F95",
    x"317760A7",
    x"317741BD",
    x"317722D6",
    x"317703F4",
    x"3176E515",
    x"3176C63B",
    x"3176A764",
    x"31768891",
    x"317669C2",
    x"31764AF6",
    x"31762C2F",
    x"31760D6B",
    x"3175EEAC",
    x"3175CFF0",
    x"3175B138",
    x"31759283",
    x"317573D3",
    x"31755526",
    x"3175367E",
    x"317517D9",
    x"3174F938",
    x"3174DA9A",
    x"3174BC01",
    x"31749D6B",
    x"31747EDA",
    x"3174604C",
    x"317441C2",
    x"3174233B",
    x"317404B9",
    x"3173E63A",
    x"3173C7BF",
    x"3173A948",
    x"31738AD5",
    x"31736C65",
    x"31734DFA",
    x"31732F92",
    x"3173112E",
    x"3172F2CE",
    x"3172D471",
    x"3172B619",
    x"317297C4",
    x"31727973",
    x"31725B25",
    x"31723CDC",
    x"31721E96",
    x"31720054",
    x"3171E216",
    x"3171C3DC",
    x"3171A5A5",
    x"31718772",
    x"31716943",
    x"31714B18",
    x"31712CF0",
    x"31710ECD",
    x"3170F0AD",
    x"3170D290",
    x"3170B478",
    x"31709663",
    x"31707852",
    x"31705A45",
    x"31703C3C",
    x"31701E36",
    x"31700034",
    x"316FE236",
    x"316FC43C",
    x"316FA645",
    x"316F8852",
    x"316F6A63",
    x"316F4C78",
    x"316F2E90",
    x"316F10AC",
    x"316EF2CC",
    x"316ED4EF",
    x"316EB717",
    x"316E9941",
    x"316E7B70",
    x"316E5DA3",
    x"316E3FD9",
    x"316E2213",
    x"316E0450",
    x"316DE692",
    x"316DC8D7",
    x"316DAB1F",
    x"316D8D6C",
    x"316D6FBC",
    x"316D5210",
    x"316D3468",
    x"316D16C3",
    x"316CF922",
    x"316CDB85",
    x"316CBDEB",
    x"316CA055",
    x"316C82C3",
    x"316C6534",
    x"316C47AA",
    x"316C2A22",
    x"316C0C9F",
    x"316BEF1F",
    x"316BD1A3",
    x"316BB42B",
    x"316B96B6",
    x"316B7945",
    x"316B5BD8",
    x"316B3E6E",
    x"316B2108",
    x"316B03A6",
    x"316AE647",
    x"316AC8EC",
    x"316AAB95",
    x"316A8E42",
    x"316A70F2",
    x"316A53A5",
    x"316A365D",
    x"316A1918",
    x"3169FBD6",
    x"3169DE99",
    x"3169C15F",
    x"3169A428",
    x"316986F6",
    x"316969C7",
    x"31694C9B",
    x"31692F73",
    x"3169124F",
    x"3168F52F",
    x"3168D812",
    x"3168BAF9",
    x"31689DE3",
    x"316880D1",
    x"316863C3",
    x"316846B8",
    x"316829B1",
    x"31680CAE",
    x"3167EFAE",
    x"3167D2B2",
    x"3167B5BA",
    x"316798C5",
    x"31677BD3",
    x"31675EE6",
    x"316741FC",
    x"31672515",
    x"31670832",
    x"3166EB53",
    x"3166CE78",
    x"3166B1A0",
    x"316694CB",
    x"316677FA",
    x"31665B2D",
    x"31663E64",
    x"3166219E",
    x"316604DB",
    x"3165E81C",
    x"3165CB61",
    x"3165AEAA",
    x"316591F5",
    x"31657545",
    x"31655898",
    x"31653BEF",
    x"31651F49",
    x"316502A7",
    x"3164E609",
    x"3164C96E",
    x"3164ACD6",
    x"31649042",
    x"316473B2",
    x"31645725",
    x"31643A9C",
    x"31641E17",
    x"31640195",
    x"3163E516",
    x"3163C89C",
    x"3163AC24",
    x"31638FB0",
    x"31637340",
    x"316356D4",
    x"31633A6B",
    x"31631E05",
    x"316301A3",
    x"3162E545",
    x"3162C8EA",
    x"3162AC92",
    x"3162903F",
    x"316273EE",
    x"316257A2",
    x"31623B58",
    x"31621F13",
    x"316202D1",
    x"3161E692",
    x"3161CA57",
    x"3161AE20",
    x"316191EC",
    x"316175BB",
    x"3161598E",
    x"31613D65",
    x"3161213F",
    x"3161051C",
    x"3160E8FD",
    x"3160CCE2",
    x"3160B0CA",
    x"316094B6",
    x"316078A5",
    x"31605C98",
    x"3160408E",
    x"31602488",
    x"31600885",
    x"315FEC85",
    x"315FD08A",
    x"315FB491",
    x"315F989C",
    x"315F7CAB",
    x"315F60BD",
    x"315F44D3",
    x"315F28EC",
    x"315F0D09",
    x"315EF129",
    x"315ED54C",
    x"315EB974",
    x"315E9D9E",
    x"315E81CC",
    x"315E65FE",
    x"315E4A33",
    x"315E2E6B",
    x"315E12A7",
    x"315DF6E6",
    x"315DDB29",
    x"315DBF70",
    x"315DA3B9",
    x"315D8807",
    x"315D6C57",
    x"315D50AC",
    x"315D3503",
    x"315D195E",
    x"315CFDBD",
    x"315CE21F",
    x"315CC684",
    x"315CAAED",
    x"315C8F5A",
    x"315C73C9",
    x"315C583D",
    x"315C3CB3",
    x"315C212E",
    x"315C05AB",
    x"315BEA2C",
    x"315BCEB1",
    x"315BB338",
    x"315B97C4",
    x"315B7C53",
    x"315B60E5",
    x"315B457A",
    x"315B2A13",
    x"315B0EB0",
    x"315AF350",
    x"315AD7F3",
    x"315ABC9A",
    x"315AA144",
    x"315A85F1",
    x"315A6AA2",
    x"315A4F57",
    x"315A340E",
    x"315A18CA",
    x"3159FD88",
    x"3159E24A",
    x"3159C710",
    x"3159ABD9",
    x"315990A5",
    x"31597574",
    x"31595A47",
    x"31593F1E",
    x"315923F8",
    x"315908D5",
    x"3158EDB5",
    x"3158D299",
    x"3158B781",
    x"31589C6B",
    x"3158815A",
    x"3158664B",
    x"31584B40",
    x"31583038",
    x"31581534",
    x"3157FA33",
    x"3157DF35",
    x"3157C43B",
    x"3157A944",
    x"31578E51",
    x"31577361",
    x"31575874",
    x"31573D8B",
    x"315722A5",
    x"315707C2",
    x"3156ECE3",
    x"3156D207",
    x"3156B72E",
    x"31569C59",
    x"31568187",
    x"315666B9",
    x"31564BED",
    x"31563126",
    x"31561661",
    x"3155FBA0",
    x"3155E0E2",
    x"3155C628",
    x"3155AB71",
    x"315590BD",
    x"3155760D",
    x"31555B5F",
    x"315540B6",
    x"3155260F",
    x"31550B6C",
    x"3154F0CC",
    x"3154D630",
    x"3154BB97",
    x"3154A101",
    x"3154866F",
    x"31546BDF",
    x"31545154",
    x"315436CB",
    x"31541C46",
    x"315401C4",
    x"3153E746",
    x"3153CCCA",
    x"3153B252",
    x"315397DE",
    x"31537D6C",
    x"315362FE",
    x"31534894",
    x"31532E2C",
    x"315313C8",
    x"3152F967",
    x"3152DF0A",
    x"3152C4AF",
    x"3152AA59",
    x"31529005",
    x"315275B5",
    x"31525B67",
    x"3152411E",
    x"315226D7",
    x"31520C94",
    x"3151F254",
    x"3151D817",
    x"3151BDDE",
    x"3151A3A8",
    x"31518975",
    x"31516F46",
    x"31515519",
    x"31513AF0",
    x"315120CB",
    x"315106A8",
    x"3150EC89",
    x"3150D26D",
    x"3150B854",
    x"31509E3F",
    x"3150842D",
    x"31506A1E",
    x"31505012",
    x"3150360A",
    x"31501C05",
    x"31500203",
    x"314FE804",
    x"314FCE09",
    x"314FB411",
    x"314F9A1C",
    x"314F802A",
    x"314F663C",
    x"314F4C51",
    x"314F3269",
    x"314F1884",
    x"314EFEA3",
    x"314EE4C4",
    x"314ECAE9",
    x"314EB112",
    x"314E973D",
    x"314E7D6C",
    x"314E639E",
    x"314E49D3",
    x"314E300B",
    x"314E1647",
    x"314DFC86",
    x"314DE2C8",
    x"314DC90D",
    x"314DAF55",
    x"314D95A1",
    x"314D7BF0",
    x"314D6242",
    x"314D4897",
    x"314D2EF0",
    x"314D154C",
    x"314CFBAB",
    x"314CE20D",
    x"314CC872",
    x"314CAEDB",
    x"314C9546",
    x"314C7BB5",
    x"314C6228",
    x"314C489D",
    x"314C2F15",
    x"314C1591",
    x"314BFC10",
    x"314BE292",
    x"314BC917",
    x"314BAFA0",
    x"314B962B",
    x"314B7CBA",
    x"314B634C",
    x"314B49E1",
    x"314B307A",
    x"314B1715",
    x"314AFDB4",
    x"314AE456",
    x"314ACAFB",
    x"314AB1A3",
    x"314A984F",
    x"314A7EFD",
    x"314A65AF",
    x"314A4C64",
    x"314A331C",
    x"314A19D7",
    x"314A0095",
    x"3149E757",
    x"3149CE1B",
    x"3149B4E3",
    x"31499BAE",
    x"3149827C",
    x"3149694E",
    x"31495022",
    x"314936FA",
    x"31491DD4",
    x"314904B2",
    x"3148EB93",
    x"3148D277",
    x"3148B95E",
    x"3148A049",
    x"31488736",
    x"31486E27",
    x"3148551B",
    x"31483C12",
    x"3148230C",
    x"31480A09",
    x"3147F109",
    x"3147D80D",
    x"3147BF13",
    x"3147A61D",
    x"31478D2A",
    x"3147743A",
    x"31475B4D",
    x"31474263",
    x"3147297C",
    x"31471098",
    x"3146F7B8",
    x"3146DEDB",
    x"3146C600",
    x"3146AD29",
    x"31469455",
    x"31467B84",
    x"314662B6",
    x"314649EB",
    x"31463124",
    x"3146185F",
    x"3145FF9D",
    x"3145E6DF",
    x"3145CE24",
    x"3145B56C",
    x"31459CB6",
    x"31458404",
    x"31456B55",
    x"314552AA",
    x"31453A01",
    x"3145215B",
    x"314508B8",
    x"3144F019",
    x"3144D77C",
    x"3144BEE3",
    x"3144A64D",
    x"31448DB9",
    x"31447529",
    x"31445C9C",
    x"31444412",
    x"31442B8B",
    x"31441307",
    x"3143FA86",
    x"3143E209",
    x"3143C98E",
    x"3143B116",
    x"314398A2",
    x"31438030",
    x"314367C1",
    x"31434F56",
    x"314336EE",
    x"31431E88",
    x"31430626",
    x"3142EDC7",
    x"3142D56B",
    x"3142BD11",
    x"3142A4BB",
    x"31428C68",
    x"31427418",
    x"31425BCB",
    x"31424381",
    x"31422B3A",
    x"314212F6",
    x"3141FAB6",
    x"3141E278",
    x"3141CA3D",
    x"3141B205",
    x"314199D0",
    x"3141819F",
    x"31416970",
    x"31415144",
    x"3141391C",
    x"314120F6",
    x"314108D4",
    x"3140F0B4",
    x"3140D897",
    x"3140C07E",
    x"3140A867",
    x"31409054",
    x"31407843",
    x"31406036",
    x"3140482B",
    x"31403024",
    x"3140181F",
    x"3140001E",
    x"313FE81F",
    x"313FD023",
    x"313FB82B",
    x"313FA035",
    x"313F8843",
    x"313F7053",
    x"313F5867",
    x"313F407D",
    x"313F2897",
    x"313F10B3",
    x"313EF8D3",
    x"313EE0F5",
    x"313EC91A",
    x"313EB143",
    x"313E996E",
    x"313E819C",
    x"313E69CE",
    x"313E5202",
    x"313E3A39",
    x"313E2273",
    x"313E0AB0",
    x"313DF2F1",
    x"313DDB34",
    x"313DC37A",
    x"313DABC3",
    x"313D940F",
    x"313D7C5E",
    x"313D64B0",
    x"313D4D05",
    x"313D355D",
    x"313D1DB7",
    x"313D0615",
    x"313CEE76",
    x"313CD6D9",
    x"313CBF40",
    x"313CA7AA",
    x"313C9016",
    x"313C7886",
    x"313C60F8",
    x"313C496D",
    x"313C31E6",
    x"313C1A61",
    x"313C02DF",
    x"313BEB60",
    x"313BD3E4",
    x"313BBC6B",
    x"313BA4F5",
    x"313B8D82",
    x"313B7612",
    x"313B5EA4",
    x"313B473A",
    x"313B2FD3",
    x"313B186E",
    x"313B010D",
    x"313AE9AE",
    x"313AD252",
    x"313ABAF9",
    x"313AA3A3",
    x"313A8C50",
    x"313A7500",
    x"313A5DB3",
    x"313A4669",
    x"313A2F22",
    x"313A17DD",
    x"313A009C",
    x"3139E95D",
    x"3139D221",
    x"3139BAE8",
    x"3139A3B3",
    x"31398C80",
    x"3139754F",
    x"31395E22",
    x"313946F8",
    x"31392FD0",
    x"313918AC",
    x"3139018A",
    x"3138EA6C",
    x"3138D350",
    x"3138BC37",
    x"3138A521",
    x"31388E0D",
    x"313876FD",
    x"31385FF0",
    x"313848E5",
    x"313831DD",
    x"31381AD9",
    x"313803D7",
    x"3137ECD8",
    x"3137D5DC",
    x"3137BEE2",
    x"3137A7EC",
    x"313790F8",
    x"31377A08",
    x"3137631A",
    x"31374C2F",
    x"31373547",
    x"31371E61",
    x"3137077F",
    x"3136F0A0",
    x"3136D9C3",
    x"3136C2E9",
    x"3136AC12",
    x"3136953E",
    x"31367E6D",
    x"3136679F",
    x"313650D3",
    x"31363A0A",
    x"31362344",
    x"31360C81",
    x"3135F5C1",
    x"3135DF04",
    x"3135C84A",
    x"3135B192",
    x"31359ADD",
    x"3135842B",
    x"31356D7C",
    x"313556D0",
    x"31354026",
    x"31352980",
    x"313512DC",
    x"3134FC3B",
    x"3134E59D",
    x"3134CF02",
    x"3134B869",
    x"3134A1D4",
    x"31348B41",
    x"313474B1",
    x"31345E24",
    x"31344799",
    x"31343112",
    x"31341A8D",
    x"3134040B",
    x"3133ED8C",
    x"3133D710",
    x"3133C096",
    x"3133AA20",
    x"313393AC",
    x"31337D3B",
    x"313366CC",
    x"31335061",
    x"313339F8",
    x"31332392",
    x"31330D2F",
    x"3132F6CF",
    x"3132E072",
    x"3132CA17",
    x"3132B3BF",
    x"31329D6A",
    x"31328718",
    x"313270C8",
    x"31325A7C",
    x"31324432",
    x"31322DEB",
    x"313217A6",
    x"31320165",
    x"3131EB26",
    x"3131D4EA",
    x"3131BEB1",
    x"3131A87A",
    x"31319247",
    x"31317C16",
    x"313165E8",
    x"31314FBC",
    x"31313994",
    x"3131236E",
    x"31310D4B",
    x"3130F72A",
    x"3130E10D",
    x"3130CAF2",
    x"3130B4DA",
    x"31309EC5",
    x"313088B3",
    x"313072A3",
    x"31305C96",
    x"3130468C",
    x"31303084",
    x"31301A80",
    x"3130047E",
    x"312FEE7E",
    x"312FD882",
    x"312FC288",
    x"312FAC91",
    x"312F969D",
    x"312F80AC",
    x"312F6ABD",
    x"312F54D1",
    x"312F3EE8",
    x"312F2901",
    x"312F131E",
    x"312EFD3C",
    x"312EE75E",
    x"312ED183",
    x"312EBBAA",
    x"312EA5D4",
    x"312E9000",
    x"312E7A30",
    x"312E6462",
    x"312E4E97",
    x"312E38CE",
    x"312E2308",
    x"312E0D45",
    x"312DF785",
    x"312DE1C8",
    x"312DCC0D",
    x"312DB655",
    x"312DA09F",
    x"312D8AEC",
    x"312D753C",
    x"312D5F8F",
    x"312D49E4",
    x"312D343D",
    x"312D1E97",
    x"312D08F5",
    x"312CF355",
    x"312CDDB8",
    x"312CC81E",
    x"312CB286",
    x"312C9CF1",
    x"312C875F",
    x"312C71CF",
    x"312C5C42",
    x"312C46B8",
    x"312C3131",
    x"312C1BAC",
    x"312C062A",
    x"312BF0AA",
    x"312BDB2E",
    x"312BC5B4",
    x"312BB03C",
    x"312B9AC7",
    x"312B8555",
    x"312B6FE6",
    x"312B5A7A",
    x"312B4510",
    x"312B2FA8",
    x"312B1A44",
    x"312B04E2",
    x"312AEF82",
    x"312ADA26",
    x"312AC4CC",
    x"312AAF75",
    x"312A9A20",
    x"312A84CE",
    x"312A6F7F",
    x"312A5A32",
    x"312A44E8",
    x"312A2FA1",
    x"312A1A5C",
    x"312A051A",
    x"3129EFDB",
    x"3129DA9E",
    x"3129C564",
    x"3129B02D",
    x"31299AF8",
    x"312985C6",
    x"31297097",
    x"31295B6A",
    x"31294640",
    x"31293119",
    x"31291BF4",
    x"312906D2",
    x"3128F1B2",
    x"3128DC95",
    x"3128C77B",
    x"3128B263",
    x"31289D4E",
    x"3128883C",
    x"3128732C",
    x"31285E1F",
    x"31284915",
    x"3128340D",
    x"31281F08",
    x"31280A05",
    x"3127F505",
    x"3127E008",
    x"3127CB0D",
    x"3127B615",
    x"3127A120",
    x"31278C2D",
    x"3127773D",
    x"3127624F",
    x"31274D64",
    x"3127387C",
    x"31272396",
    x"31270EB3",
    x"3126F9D2",
    x"3126E4F4",
    x"3126D019",
    x"3126BB40",
    x"3126A66A",
    x"31269197",
    x"31267CC6",
    x"312667F8",
    x"3126532C",
    x"31263E63",
    x"3126299C",
    x"312614D8",
    x"31260017",
    x"3125EB58",
    x"3125D69C",
    x"3125C1E3",
    x"3125AD2C",
    x"31259877",
    x"312583C6",
    x"31256F16",
    x"31255A6A",
    x"312545C0",
    x"31253118",
    x"31251C74",
    x"312507D1",
    x"3124F332",
    x"3124DE94",
    x"3124C9FA",
    x"3124B562",
    x"3124A0CD",
    x"31248C3A",
    x"312477AA",
    x"3124631C",
    x"31244E91",
    x"31243A08",
    x"31242582",
    x"312410FF",
    x"3123FC7E",
    x"3123E800",
    x"3123D384",
    x"3123BF0B",
    x"3123AA94",
    x"31239620",
    x"312381AF",
    x"31236D40",
    x"312358D3",
    x"3123446A",
    x"31233002",
    x"31231B9E",
    x"3123073B",
    x"3122F2DC",
    x"3122DE7F",
    x"3122CA24",
    x"3122B5CC",
    x"3122A177",
    x"31228D24",
    x"312278D3",
    x"31226486",
    x"3122503A",
    x"31223BF2",
    x"312227AB",
    x"31221368",
    x"3121FF26",
    x"3121EAE8",
    x"3121D6AC",
    x"3121C272",
    x"3121AE3B",
    x"31219A07",
    x"312185D5",
    x"312171A5",
    x"31215D78",
    x"3121494E",
    x"31213526",
    x"31212100",
    x"31210CDE",
    x"3120F8BD",
    x"3120E49F",
    x"3120D084",
    x"3120BC6B",
    x"3120A855",
    x"31209441",
    x"31208030",
    x"31206C21",
    x"31205815",
    x"3120440B",
    x"31203004",
    x"31201BFF",
    x"312007FD",
    x"311FF3FD",
    x"311FE000",
    x"311FCC05",
    x"311FB80D",
    x"311FA417",
    x"311F9024",
    x"311F7C33",
    x"311F6845",
    x"311F5459",
    x"311F4070",
    x"311F2C89",
    x"311F18A5",
    x"311F04C3",
    x"311EF0E3",
    x"311EDD07",
    x"311EC92C",
    x"311EB554",
    x"311EA17F",
    x"311E8DAC",
    x"311E79DB",
    x"311E660D",
    x"311E5242",
    x"311E3E79",
    x"311E2AB2",
    x"311E16EE",
    x"311E032D",
    x"311DEF6D",
    x"311DDBB1",
    x"311DC7F6",
    x"311DB43F",
    x"311DA089",
    x"311D8CD7",
    x"311D7926",
    x"311D6578",
    x"311D51CD",
    x"311D3E24",
    x"311D2A7D",
    x"311D16D9",
    x"311D0338",
    x"311CEF98",
    x"311CDBFC",
    x"311CC861",
    x"311CB4CA",
    x"311CA134",
    x"311C8DA1",
    x"311C7A11",
    x"311C6683",
    x"311C52F7",
    x"311C3F6E",
    x"311C2BE7",
    x"311C1863",
    x"311C04E1",
    x"311BF162",
    x"311BDDE5",
    x"311BCA6A",
    x"311BB6F2",
    x"311BA37D",
    x"311B9009",
    x"311B7C99",
    x"311B692A",
    x"311B55BE",
    x"311B4255",
    x"311B2EEE",
    x"311B1B89",
    x"311B0827",
    x"311AF4C7",
    x"311AE16A",
    x"311ACE0F",
    x"311ABAB6",
    x"311AA760",
    x"311A940C",
    x"311A80BB",
    x"311A6D6C",
    x"311A5A20",
    x"311A46D6",
    x"311A338E",
    x"311A2049",
    x"311A0D06",
    x"3119F9C5",
    x"3119E687",
    x"3119D34C",
    x"3119C013",
    x"3119ACDC",
    x"311999A7",
    x"31198675",
    x"31197346",
    x"31196019",
    x"31194CEE",
    x"311939C5",
    x"3119269F",
    x"3119137C",
    x"3119005A",
    x"3118ED3C",
    x"3118DA1F",
    x"3118C705",
    x"3118B3ED",
    x"3118A0D8",
    x"31188DC5",
    x"31187AB5",
    x"311867A6",
    x"3118549B",
    x"31184191",
    x"31182E8A",
    x"31181B86",
    x"31180883",
    x"3117F584",
    x"3117E286",
    x"3117CF8B",
    x"3117BC92",
    x"3117A99C",
    x"311796A8",
    x"311783B6",
    x"311770C7",
    x"31175DDA",
    x"31174AEF",
    x"31173807",
    x"31172521",
    x"3117123E",
    x"3116FF5D",
    x"3116EC7E",
    x"3116D9A2",
    x"3116C6C8",
    x"3116B3F0",
    x"3116A11B",
    x"31168E48",
    x"31167B77",
    x"311668A9",
    x"311655DD",
    x"31164313",
    x"3116304C",
    x"31161D87",
    x"31160AC5",
    x"3115F805",
    x"3115E547",
    x"3115D28B",
    x"3115BFD2",
    x"3115AD1B",
    x"31159A67",
    x"311587B5",
    x"31157505",
    x"31156257",
    x"31154FAC",
    x"31153D04",
    x"31152A5D",
    x"311517B9",
    x"31150517",
    x"3114F278",
    x"3114DFDB",
    x"3114CD40",
    x"3114BAA7",
    x"3114A811",
    x"3114957D",
    x"311482EC",
    x"3114705C",
    x"31145DD0",
    x"31144B45",
    x"311438BD",
    x"31142637",
    x"311413B3",
    x"31140132",
    x"3113EEB3",
    x"3113DC36",
    x"3113C9BC",
    x"3113B744",
    x"3113A4CE",
    x"3113925B",
    x"31137FE9",
    x"31136D7B",
    x"31135B0E",
    x"311348A4",
    x"3113363C",
    x"311323D6",
    x"31131173",
    x"3112FF12",
    x"3112ECB3",
    x"3112DA57",
    x"3112C7FD",
    x"3112B5A5",
    x"3112A34F",
    x"311290FC",
    x"31127EAB",
    x"31126C5C",
    x"31125A10",
    x"311247C6",
    x"3112357E",
    x"31122338",
    x"311210F5",
    x"3111FEB4",
    x"3111EC75",
    x"3111DA39",
    x"3111C7FF",
    x"3111B5C7",
    x"3111A391",
    x"3111915E",
    x"31117F2D",
    x"31116CFE",
    x"31115AD2",
    x"311148A8",
    x"31113680",
    x"3111245A",
    x"31111237",
    x"31110015",
    x"3110EDF7",
    x"3110DBDA",
    x"3110C9C0",
    x"3110B7A8",
    x"3110A592",
    x"3110937E",
    x"3110816D",
    x"31106F5E",
    x"31105D51",
    x"31104B46",
    x"3110393E",
    x"31102738",
    x"31101534",
    x"31100333",
    x"310FF134",
    x"310FDF37",
    x"310FCD3C",
    x"310FBB43",
    x"310FA94D",
    x"310F9759",
    x"310F8567",
    x"310F7378",
    x"310F618A",
    x"310F4F9F",
    x"310F3DB6",
    x"310F2BD0",
    x"310F19EB",
    x"310F0809",
    x"310EF629",
    x"310EE44C",
    x"310ED270",
    x"310EC097",
    x"310EAEC0",
    x"310E9CEB",
    x"310E8B19",
    x"310E7949",
    x"310E677B",
    x"310E55AF",
    x"310E43E5",
    x"310E321E",
    x"310E2059",
    x"310E0E96",
    x"310DFCD5",
    x"310DEB17",
    x"310DD95A",
    x"310DC7A0",
    x"310DB5E8",
    x"310DA433",
    x"310D927F",
    x"310D80CE",
    x"310D6F1F",
    x"310D5D72",
    x"310D4BC8",
    x"310D3A1F",
    x"310D2879",
    x"310D16D5",
    x"310D0533",
    x"310CF394",
    x"310CE1F7",
    x"310CD05B",
    x"310CBEC2",
    x"310CAD2C",
    x"310C9B97",
    x"310C8A05",
    x"310C7875",
    x"310C66E7",
    x"310C555B",
    x"310C43D1",
    x"310C324A",
    x"310C20C5",
    x"310C0F42",
    x"310BFDC1",
    x"310BEC42",
    x"310BDAC6",
    x"310BC94C",
    x"310BB7D4",
    x"310BA65E",
    x"310B94EA",
    x"310B8378",
    x"310B7209",
    x"310B609C",
    x"310B4F31",
    x"310B3DC8",
    x"310B2C62",
    x"310B1AFD",
    x"310B099B",
    x"310AF83B",
    x"310AE6DD",
    x"310AD581",
    x"310AC427",
    x"310AB2D0",
    x"310AA17B",
    x"310A9028",
    x"310A7ED7",
    x"310A6D88",
    x"310A5C3B",
    x"310A4AF1",
    x"310A39A9",
    x"310A2862",
    x"310A171E",
    x"310A05DD",
    x"3109F49D",
    x"3109E35F",
    x"3109D224",
    x"3109C0EB",
    x"3109AFB4",
    x"31099E7F",
    x"31098D4C",
    x"31097C1C",
    x"31096AED",
    x"310959C1",
    x"31094897",
    x"3109376F",
    x"31092649",
    x"31091525",
    x"31090404",
    x"3108F2E4",
    x"3108E1C7",
    x"3108D0AC",
    x"3108BF93",
    x"3108AE7C",
    x"31089D67",
    x"31088C55",
    x"31087B44",
    x"31086A36",
    x"31085929",
    x"3108481F",
    x"31083717",
    x"31082612",
    x"3108150E",
    x"3108040C",
    x"3107F30D",
    x"3107E210",
    x"3107D114",
    x"3107C01B",
    x"3107AF24",
    x"31079E30",
    x"31078D3D",
    x"31077C4C",
    x"31076B5E",
    x"31075A71",
    x"31074987",
    x"3107389F",
    x"310727B9",
    x"310716D5",
    x"310705F3",
    x"3106F514",
    x"3106E436",
    x"3106D35B",
    x"3106C281",
    x"3106B1AA",
    x"3106A0D5",
    x"31069002",
    x"31067F31",
    x"31066E62",
    x"31065D95",
    x"31064CCB",
    x"31063C02",
    x"31062B3C",
    x"31061A77",
    x"310609B5",
    x"3105F8F5",
    x"3105E837",
    x"3105D77B",
    x"3105C6C1",
    x"3105B609",
    x"3105A553",
    x"310594A0",
    x"310583EE",
    x"3105733F",
    x"31056291",
    x"310551E6",
    x"3105413D",
    x"31053096",
    x"31051FF1",
    x"31050F4E",
    x"3104FEAD",
    x"3104EE0E",
    x"3104DD71",
    x"3104CCD7",
    x"3104BC3E",
    x"3104ABA8",
    x"31049B13",
    x"31048A81",
    x"310479F1",
    x"31046962",
    x"310458D6",
    x"3104484C",
    x"310437C4",
    x"3104273E",
    x"310416BA",
    x"31040639",
    x"3103F5B9",
    x"3103E53B",
    x"3103D4C0",
    x"3103C446",
    x"3103B3CE",
    x"3103A359",
    x"310392E6",
    x"31038274",
    x"31037205",
    x"31036198",
    x"3103512D",
    x"310340C3",
    x"3103305C",
    x"31031FF7",
    x"31030F94",
    x"3102FF33",
    x"3102EED5",
    x"3102DE78",
    x"3102CE1D",
    x"3102BDC4",
    x"3102AD6E",
    x"31029D19",
    x"31028CC6",
    x"31027C76",
    x"31026C27",
    x"31025BDB",
    x"31024B90",
    x"31023B48",
    x"31022B01",
    x"31021ABD",
    x"31020A7B",
    x"3101FA3A",
    x"3101E9FC",
    x"3101D9C0",
    x"3101C986",
    x"3101B94E",
    x"3101A917",
    x"310198E3",
    x"310188B1",
    x"31017881",
    x"31016853",
    x"31015827",
    x"310147FD",
    x"310137D5",
    x"310127AF",
    x"3101178B",
    x"31010769",
    x"3100F749",
    x"3100E72B",
    x"3100D70F",
    x"3100C6F6",
    x"3100B6DE",
    x"3100A6C8",
    x"310096B4",
    x"310086A2",
    x"31007692",
    x"31006685",
    x"31005679",
    x"3100466F",
    x"31003667",
    x"31002661",
    x"3100165D",
    x"3100065C",
    x"30FFECB8",
    x"30FFCCBC",
    x"30FFACC5",
    x"30FF8CD1",
    x"30FF6CE1",
    x"30FF4CF6",
    x"30FF2D0E",
    x"30FF0D2B",
    x"30FEED4B",
    x"30FECD6F",
    x"30FEAD98",
    x"30FE8DC4",
    x"30FE6DF4",
    x"30FE4E28",
    x"30FE2E61",
    x"30FE0E9D",
    x"30FDEEDD",
    x"30FDCF21",
    x"30FDAF69",
    x"30FD8FB5",
    x"30FD7005",
    x"30FD5059",
    x"30FD30B1",
    x"30FD110D",
    x"30FCF16D",
    x"30FCD1D1",
    x"30FCB238",
    x"30FC92A4",
    x"30FC7314",
    x"30FC5387",
    x"30FC33FF",
    x"30FC147A",
    x"30FBF4FA",
    x"30FBD57D",
    x"30FBB604",
    x"30FB9690",
    x"30FB771F",
    x"30FB57B2",
    x"30FB3849",
    x"30FB18E4",
    x"30FAF983",
    x"30FADA25",
    x"30FABACC",
    x"30FA9B77",
    x"30FA7C25",
    x"30FA5CD8",
    x"30FA3D8E",
    x"30FA1E48",
    x"30F9FF06",
    x"30F9DFC8",
    x"30F9C08E",
    x"30F9A158",
    x"30F98226",
    x"30F962F8",
    x"30F943CD",
    x"30F924A7",
    x"30F90584",
    x"30F8E665",
    x"30F8C74B",
    x"30F8A834",
    x"30F88921",
    x"30F86A11",
    x"30F84B06",
    x"30F82BFF",
    x"30F80CFB",
    x"30F7EDFB",
    x"30F7CF00",
    x"30F7B008",
    x"30F79113",
    x"30F77223",
    x"30F75337",
    x"30F7344E",
    x"30F7156A",
    x"30F6F689",
    x"30F6D7AC",
    x"30F6B8D3",
    x"30F699FE",
    x"30F67B2D",
    x"30F65C5F",
    x"30F63D96",
    x"30F61ED0",
    x"30F6000E",
    x"30F5E150",
    x"30F5C296",
    x"30F5A3DF",
    x"30F5852D",
    x"30F5667E",
    x"30F547D3",
    x"30F5292C",
    x"30F50A89",
    x"30F4EBE9",
    x"30F4CD4E",
    x"30F4AEB6",
    x"30F49022",
    x"30F47192",
    x"30F45306",
    x"30F4347D",
    x"30F415F9",
    x"30F3F778",
    x"30F3D8FB",
    x"30F3BA81",
    x"30F39C0C",
    x"30F37D9A",
    x"30F35F2D",
    x"30F340C3",
    x"30F3225C",
    x"30F303FA",
    x"30F2E59B",
    x"30F2C741",
    x"30F2A8EA",
    x"30F28A96",
    x"30F26C47",
    x"30F24DFB",
    x"30F22FB3",
    x"30F2116F",
    x"30F1F32F",
    x"30F1D4F3",
    x"30F1B6BA",
    x"30F19885",
    x"30F17A54",
    x"30F15C26",
    x"30F13DFD",
    x"30F11FD7",
    x"30F101B5",
    x"30F0E396",
    x"30F0C57C",
    x"30F0A765",
    x"30F08952",
    x"30F06B43",
    x"30F04D37",
    x"30F02F2F",
    x"30F0112B",
    x"30EFF32B",
    x"30EFD52F",
    x"30EFB736",
    x"30EF9941",
    x"30EF7B50",
    x"30EF5D62",
    x"30EF3F78",
    x"30EF2192",
    x"30EF03B0",
    x"30EEE5D1",
    x"30EEC7F6",
    x"30EEAA1F",
    x"30EE8C4C",
    x"30EE6E7C",
    x"30EE50B0",
    x"30EE32E8",
    x"30EE1523",
    x"30EDF763",
    x"30EDD9A6",
    x"30EDBBEC",
    x"30ED9E37",
    x"30ED8085",
    x"30ED62D6",
    x"30ED452C",
    x"30ED2785",
    x"30ED09E2",
    x"30ECEC43",
    x"30ECCEA7",
    x"30ECB10F",
    x"30EC937B",
    x"30EC75EA",
    x"30EC585D",
    x"30EC3AD4",
    x"30EC1D4F",
    x"30EBFFCD",
    x"30EBE24F",
    x"30EBC4D4",
    x"30EBA75D",
    x"30EB89EA",
    x"30EB6C7B",
    x"30EB4F0F",
    x"30EB31A7",
    x"30EB1443",
    x"30EAF6E2",
    x"30EAD985",
    x"30EABC2C",
    x"30EA9ED6",
    x"30EA8184",
    x"30EA6436",
    x"30EA46EB",
    x"30EA29A4",
    x"30EA0C61",
    x"30E9EF21",
    x"30E9D1E5",
    x"30E9B4AC",
    x"30E99778",
    x"30E97A47",
    x"30E95D19",
    x"30E93FEF",
    x"30E922C9",
    x"30E905A7",
    x"30E8E888",
    x"30E8CB6C",
    x"30E8AE55",
    x"30E89141",
    x"30E87430",
    x"30E85724",
    x"30E83A1B",
    x"30E81D15",
    x"30E80013",
    x"30E7E315",
    x"30E7C61B",
    x"30E7A924",
    x"30E78C30",
    x"30E76F41",
    x"30E75255",
    x"30E7356C",
    x"30E71887",
    x"30E6FBA6",
    x"30E6DEC8",
    x"30E6C1EE",
    x"30E6A518",
    x"30E68845",
    x"30E66B76",
    x"30E64EAA",
    x"30E631E2",
    x"30E6151E",
    x"30E5F85D",
    x"30E5DBA0",
    x"30E5BEE6",
    x"30E5A230",
    x"30E5857D",
    x"30E568CE",
    x"30E54C23",
    x"30E52F7B",
    x"30E512D7",
    x"30E4F637",
    x"30E4D99A",
    x"30E4BD00",
    x"30E4A06A",
    x"30E483D8",
    x"30E46749",
    x"30E44ABE",
    x"30E42E37",
    x"30E411B3",
    x"30E3F532",
    x"30E3D8B6",
    x"30E3BC3C",
    x"30E39FC6",
    x"30E38354",
    x"30E366E6",
    x"30E34A7B",
    x"30E32E13",
    x"30E311AF",
    x"30E2F54F",
    x"30E2D8F2",
    x"30E2BC98",
    x"30E2A043",
    x"30E283F0",
    x"30E267A2",
    x"30E24B56",
    x"30E22F0F",
    x"30E212CB",
    x"30E1F68A",
    x"30E1DA4D",
    x"30E1BE13",
    x"30E1A1DD",
    x"30E185AB",
    x"30E1697C",
    x"30E14D51",
    x"30E13129",
    x"30E11504",
    x"30E0F8E3",
    x"30E0DCC6",
    x"30E0C0AC",
    x"30E0A496",
    x"30E08883",
    x"30E06C74",
    x"30E05068",
    x"30E03460",
    x"30E0185B",
    x"30DFFC5A",
    x"30DFE05C",
    x"30DFC462",
    x"30DFA86B",
    x"30DF8C77",
    x"30DF7088",
    x"30DF549B",
    x"30DF38B2",
    x"30DF1CCD",
    x"30DF00EB",
    x"30DEE50D",
    x"30DEC932",
    x"30DEAD5B",
    x"30DE9187",
    x"30DE75B6",
    x"30DE59E9",
    x"30DE3E20",
    x"30DE225A",
    x"30DE0697",
    x"30DDEAD8",
    x"30DDCF1C",
    x"30DDB364",
    x"30DD97B0",
    x"30DD7BFE",
    x"30DD6051",
    x"30DD44A6",
    x"30DD28FF",
    x"30DD0D5C",
    x"30DCF1BC",
    x"30DCD620",
    x"30DCBA87",
    x"30DC9EF1",
    x"30DC835F",
    x"30DC67D0",
    x"30DC4C45",
    x"30DC30BD",
    x"30DC1539",
    x"30DBF9B8",
    x"30DBDE3A",
    x"30DBC2C0",
    x"30DBA74A",
    x"30DB8BD6",
    x"30DB7067",
    x"30DB54FA",
    x"30DB3991",
    x"30DB1E2C",
    x"30DB02CA",
    x"30DAE76B",
    x"30DACC10",
    x"30DAB0B8",
    x"30DA9564",
    x"30DA7A13",
    x"30DA5EC5",
    x"30DA437B",
    x"30DA2834",
    x"30DA0CF1",
    x"30D9F1B1",
    x"30D9D675",
    x"30D9BB3C",
    x"30D9A006",
    x"30D984D4",
    x"30D969A5",
    x"30D94E79",
    x"30D93351",
    x"30D9182C",
    x"30D8FD0B",
    x"30D8E1ED",
    x"30D8C6D2",
    x"30D8ABBB",
    x"30D890A8",
    x"30D87597",
    x"30D85A8A",
    x"30D83F81",
    x"30D8247A",
    x"30D80977",
    x"30D7EE78",
    x"30D7D37C",
    x"30D7B883",
    x"30D79D8E",
    x"30D7829C",
    x"30D767AD",
    x"30D74CC2",
    x"30D731DA",
    x"30D716F5",
    x"30D6FC14",
    x"30D6E136",
    x"30D6C65C",
    x"30D6AB85",
    x"30D690B1",
    x"30D675E0",
    x"30D65B13",
    x"30D6404A",
    x"30D62583",
    x"30D60AC0",
    x"30D5F001",
    x"30D5D544",
    x"30D5BA8B",
    x"30D59FD6",
    x"30D58523",
    x"30D56A74",
    x"30D54FC9",
    x"30D53520",
    x"30D51A7B",
    x"30D4FFDA",
    x"30D4E53C",
    x"30D4CAA1",
    x"30D4B009",
    x"30D49575",
    x"30D47AE3",
    x"30D46056",
    x"30D445CB",
    x"30D42B44",
    x"30D410C1",
    x"30D3F640",
    x"30D3DBC3",
    x"30D3C149",
    x"30D3A6D3",
    x"30D38C5F",
    x"30D371F0",
    x"30D35783",
    x"30D33D1A",
    x"30D322B4",
    x"30D30851",
    x"30D2EDF2",
    x"30D2D396",
    x"30D2B93D",
    x"30D29EE7",
    x"30D28495",
    x"30D26A46",
    x"30D24FFA",
    x"30D235B2",
    x"30D21B6D",
    x"30D2012B",
    x"30D1E6ED",
    x"30D1CCB2",
    x"30D1B27A",
    x"30D19845",
    x"30D17E14",
    x"30D163E5",
    x"30D149BB",
    x"30D12F93",
    x"30D1156F",
    x"30D0FB4E",
    x"30D0E130",
    x"30D0C715",
    x"30D0ACFE",
    x"30D092EA",
    x"30D078D9",
    x"30D05ECC",
    x"30D044C2",
    x"30D02ABB",
    x"30D010B7",
    x"30CFF6B6",
    x"30CFDCB9",
    x"30CFC2BF",
    x"30CFA8C9",
    x"30CF8ED5",
    x"30CF74E5",
    x"30CF5AF8",
    x"30CF410E",
    x"30CF2728",
    x"30CF0D44",
    x"30CEF364",
    x"30CED987",
    x"30CEBFAE",
    x"30CEA5D8",
    x"30CE8C04",
    x"30CE7235",
    x"30CE5868",
    x"30CE3E9E",
    x"30CE24D8",
    x"30CE0B15",
    x"30CDF155",
    x"30CDD799",
    x"30CDBDE0",
    x"30CDA429",
    x"30CD8A77",
    x"30CD70C7",
    x"30CD571A",
    x"30CD3D71",
    x"30CD23CB",
    x"30CD0A28",
    x"30CCF088",
    x"30CCD6EC",
    x"30CCBD53",
    x"30CCA3BD",
    x"30CC8A2A",
    x"30CC709A",
    x"30CC570E",
    x"30CC3D84",
    x"30CC23FE",
    x"30CC0A7B",
    x"30CBF0FC",
    x"30CBD77F",
    x"30CBBE06",
    x"30CBA490",
    x"30CB8B1D",
    x"30CB71AD",
    x"30CB5840",
    x"30CB3ED7",
    x"30CB2570",
    x"30CB0C0D",
    x"30CAF2AD",
    x"30CAD951",
    x"30CABFF7",
    x"30CAA6A1",
    x"30CA8D4D",
    x"30CA73FD",
    x"30CA5AB0",
    x"30CA4167",
    x"30CA2820",
    x"30CA0EDD",
    x"30C9F59C",
    x"30C9DC5F",
    x"30C9C325",
    x"30C9A9EE",
    x"30C990BB",
    x"30C9778A",
    x"30C95E5D",
    x"30C94533",
    x"30C92C0C",
    x"30C912E8",
    x"30C8F9C7",
    x"30C8E0A9",
    x"30C8C78F",
    x"30C8AE77",
    x"30C89563",
    x"30C87C52",
    x"30C86344",
    x"30C84A39",
    x"30C83131",
    x"30C8182D",
    x"30C7FF2B",
    x"30C7E62D",
    x"30C7CD32",
    x"30C7B43A",
    x"30C79B45",
    x"30C78253",
    x"30C76964",
    x"30C75079",
    x"30C73790",
    x"30C71EAB",
    x"30C705C8",
    x"30C6ECE9",
    x"30C6D40D",
    x"30C6BB34",
    x"30C6A25E",
    x"30C6898C",
    x"30C670BC",
    x"30C657F0",
    x"30C63F26",
    x"30C62660",
    x"30C60D9C",
    x"30C5F4DC",
    x"30C5DC1F",
    x"30C5C365",
    x"30C5AAAE",
    x"30C591FB",
    x"30C5794A",
    x"30C5609C",
    x"30C547F2",
    x"30C52F4A",
    x"30C516A6",
    x"30C4FE05",
    x"30C4E566",
    x"30C4CCCB",
    x"30C4B433",
    x"30C49B9E",
    x"30C4830C",
    x"30C46A7D",
    x"30C451F2",
    x"30C43969",
    x"30C420E3",
    x"30C40861",
    x"30C3EFE1",
    x"30C3D765",
    x"30C3BEEB",
    x"30C3A675",
    x"30C38E02",
    x"30C37592",
    x"30C35D24",
    x"30C344BA",
    x"30C32C53",
    x"30C313EF",
    x"30C2FB8E",
    x"30C2E330",
    x"30C2CAD5",
    x"30C2B27E",
    x"30C29A29",
    x"30C281D7",
    x"30C26988",
    x"30C2513D",
    x"30C238F4",
    x"30C220AE",
    x"30C2086C",
    x"30C1F02C",
    x"30C1D7F0",
    x"30C1BFB6",
    x"30C1A780",
    x"30C18F4C",
    x"30C1771C",
    x"30C15EEF",
    x"30C146C4",
    x"30C12E9D",
    x"30C11679",
    x"30C0FE57",
    x"30C0E639",
    x"30C0CE1E",
    x"30C0B606",
    x"30C09DF0",
    x"30C085DE",
    x"30C06DCF",
    x"30C055C3",
    x"30C03DB9",
    x"30C025B3",
    x"30C00DB0",
    x"30BFF5B0",
    x"30BFDDB3",
    x"30BFC5B8",
    x"30BFADC1",
    x"30BF95CD",
    x"30BF7DDC",
    x"30BF65ED",
    x"30BF4E02",
    x"30BF361A",
    x"30BF1E35",
    x"30BF0652",
    x"30BEEE73",
    x"30BED697",
    x"30BEBEBD",
    x"30BEA6E7",
    x"30BE8F14",
    x"30BE7743",
    x"30BE5F76",
    x"30BE47AB",
    x"30BE2FE4",
    x"30BE181F",
    x"30BE005E",
    x"30BDE89F",
    x"30BDD0E4",
    x"30BDB92B",
    x"30BDA176",
    x"30BD89C3",
    x"30BD7213",
    x"30BD5A66",
    x"30BD42BC",
    x"30BD2B16",
    x"30BD1372",
    x"30BCFBD1",
    x"30BCE433",
    x"30BCCC98",
    x"30BCB500",
    x"30BC9D6A",
    x"30BC85D8",
    x"30BC6E49",
    x"30BC56BD",
    x"30BC3F33",
    x"30BC27AD",
    x"30BC1029",
    x"30BBF8A9",
    x"30BBE12B",
    x"30BBC9B1",
    x"30BBB239",
    x"30BB9AC4",
    x"30BB8352",
    x"30BB6BE3",
    x"30BB5477",
    x"30BB3D0E",
    x"30BB25A8",
    x"30BB0E45",
    x"30BAF6E4",
    x"30BADF87",
    x"30BAC82C",
    x"30BAB0D5",
    x"30BA9980",
    x"30BA822E",
    x"30BA6AE0",
    x"30BA5394",
    x"30BA3C4B",
    x"30BA2505",
    x"30BA0DC2",
    x"30B9F681",
    x"30B9DF44",
    x"30B9C809",
    x"30B9B0D2",
    x"30B9999D",
    x"30B9826B",
    x"30B96B3D",
    x"30B95411",
    x"30B93CE8",
    x"30B925C1",
    x"30B90E9E",
    x"30B8F77E",
    x"30B8E060",
    x"30B8C946",
    x"30B8B22E",
    x"30B89B19",
    x"30B88407",
    x"30B86CF8",
    x"30B855EC",
    x"30B83EE3",
    x"30B827DC",
    x"30B810D9",
    x"30B7F9D8",
    x"30B7E2DA",
    x"30B7CBDF",
    x"30B7B4E7",
    x"30B79DF2",
    x"30B78700",
    x"30B77010",
    x"30B75924",
    x"30B7423A",
    x"30B72B53",
    x"30B7146F",
    x"30B6FD8E",
    x"30B6E6B0",
    x"30B6CFD4",
    x"30B6B8FC",
    x"30B6A226",
    x"30B68B53",
    x"30B67483",
    x"30B65DB6",
    x"30B646EC",
    x"30B63024",
    x"30B61960",
    x"30B6029E",
    x"30B5EBDF",
    x"30B5D523",
    x"30B5BE6A",
    x"30B5A7B4",
    x"30B59100",
    x"30B57A4F",
    x"30B563A1",
    x"30B54CF6",
    x"30B5364E",
    x"30B51FA9",
    x"30B50906",
    x"30B4F267",
    x"30B4DBCA",
    x"30B4C530",
    x"30B4AE98",
    x"30B49804",
    x"30B48172",
    x"30B46AE4",
    x"30B45458",
    x"30B43DCF",
    x"30B42748",
    x"30B410C5",
    x"30B3FA44",
    x"30B3E3C6",
    x"30B3CD4B",
    x"30B3B6D3",
    x"30B3A05D",
    x"30B389EB",
    x"30B3737B",
    x"30B35D0E",
    x"30B346A4",
    x"30B3303C",
    x"30B319D8",
    x"30B30376",
    x"30B2ED17",
    x"30B2D6BA",
    x"30B2C061",
    x"30B2AA0A",
    x"30B293B6",
    x"30B27D65",
    x"30B26717",
    x"30B250CC",
    x"30B23A83",
    x"30B2243D",
    x"30B20DFA",
    x"30B1F7BA",
    x"30B1E17C",
    x"30B1CB41",
    x"30B1B509",
    x"30B19ED4",
    x"30B188A1",
    x"30B17272",
    x"30B15C45",
    x"30B1461B",
    x"30B12FF3",
    x"30B119CF",
    x"30B103AD",
    x"30B0ED8E",
    x"30B0D771",
    x"30B0C158",
    x"30B0AB41",
    x"30B0952D",
    x"30B07F1C",
    x"30B0690D",
    x"30B05302",
    x"30B03CF9",
    x"30B026F2",
    x"30B010EF",
    x"30AFFAEE",
    x"30AFE4F0",
    x"30AFCEF5",
    x"30AFB8FC",
    x"30AFA307",
    x"30AF8D14",
    x"30AF7723",
    x"30AF6136",
    x"30AF4B4B",
    x"30AF3563",
    x"30AF1F7E",
    x"30AF099B",
    x"30AEF3BB",
    x"30AEDDDE",
    x"30AEC804",
    x"30AEB22C",
    x"30AE9C57",
    x"30AE8685",
    x"30AE70B6",
    x"30AE5AE9",
    x"30AE451F",
    x"30AE2F58",
    x"30AE1993",
    x"30AE03D1",
    x"30ADEE12",
    x"30ADD856",
    x"30ADC29C",
    x"30ADACE5",
    x"30AD9731",
    x"30AD817F",
    x"30AD6BD0",
    x"30AD5624",
    x"30AD407B",
    x"30AD2AD4",
    x"30AD1530",
    x"30ACFF8F",
    x"30ACE9F0",
    x"30ACD454",
    x"30ACBEBB",
    x"30ACA925",
    x"30AC9391",
    x"30AC7E00",
    x"30AC6871",
    x"30AC52E6",
    x"30AC3D5D",
    x"30AC27D6",
    x"30AC1253",
    x"30ABFCD2",
    x"30ABE754",
    x"30ABD1D8",
    x"30ABBC5F",
    x"30ABA6E9",
    x"30AB9175",
    x"30AB7C05",
    x"30AB6696",
    x"30AB512B",
    x"30AB3BC2",
    x"30AB265C",
    x"30AB10F8",
    x"30AAFB98",
    x"30AAE63A",
    x"30AAD0DE",
    x"30AABB85",
    x"30AAA62F",
    x"30AA90DC",
    x"30AA7B8B",
    x"30AA663D",
    x"30AA50F1",
    x"30AA3BA9",
    x"30AA2663",
    x"30AA111F",
    x"30A9FBDE",
    x"30A9E6A0",
    x"30A9D165",
    x"30A9BC2C",
    x"30A9A6F6",
    x"30A991C2",
    x"30A97C91",
    x"30A96763",
    x"30A95237",
    x"30A93D0E",
    x"30A927E8",
    x"30A912C4",
    x"30A8FDA3",
    x"30A8E885",
    x"30A8D369",
    x"30A8BE50",
    x"30A8A93A",
    x"30A89426",
    x"30A87F15",
    x"30A86A06",
    x"30A854FA",
    x"30A83FF1",
    x"30A82AEA",
    x"30A815E6",
    x"30A800E5",
    x"30A7EBE6",
    x"30A7D6EA",
    x"30A7C1F0",
    x"30A7ACF9",
    x"30A79805",
    x"30A78313",
    x"30A76E24",
    x"30A75938",
    x"30A7444E",
    x"30A72F67",
    x"30A71A82",
    x"30A705A0",
    x"30A6F0C1",
    x"30A6DBE4",
    x"30A6C70A",
    x"30A6B232",
    x"30A69D5D",
    x"30A6888B",
    x"30A673BB",
    x"30A65EEE",
    x"30A64A23",
    x"30A6355B",
    x"30A62096",
    x"30A60BD3",
    x"30A5F713",
    x"30A5E255",
    x"30A5CD9A",
    x"30A5B8E2",
    x"30A5A42C",
    x"30A58F79",
    x"30A57AC8",
    x"30A5661A",
    x"30A5516F",
    x"30A53CC6",
    x"30A5281F",
    x"30A5137C",
    x"30A4FEDB",
    x"30A4EA3C",
    x"30A4D5A0",
    x"30A4C107",
    x"30A4AC70",
    x"30A497DB",
    x"30A4834A",
    x"30A46EBB",
    x"30A45A2E",
    x"30A445A4",
    x"30A4311D",
    x"30A41C98",
    x"30A40816",
    x"30A3F396",
    x"30A3DF19",
    x"30A3CA9E",
    x"30A3B626",
    x"30A3A1B0",
    x"30A38D3E",
    x"30A378CD",
    x"30A3645F",
    x"30A34FF4",
    x"30A33B8B",
    x"30A32725",
    x"30A312C2",
    x"30A2FE61",
    x"30A2EA02",
    x"30A2D5A6",
    x"30A2C14D",
    x"30A2ACF6",
    x"30A298A1",
    x"30A28450",
    x"30A27000",
    x"30A25BB4",
    x"30A24769",
    x"30A23322",
    x"30A21EDD",
    x"30A20A9A",
    x"30A1F65A",
    x"30A1E21C",
    x"30A1CDE1",
    x"30A1B9A9",
    x"30A1A573",
    x"30A19140",
    x"30A17D0F",
    x"30A168E0",
    x"30A154B4",
    x"30A1408B",
    x"30A12C64",
    x"30A11840",
    x"30A1041E",
    x"30A0EFFF",
    x"30A0DBE2",
    x"30A0C7C8",
    x"30A0B3B0",
    x"30A09F9B",
    x"30A08B88",
    x"30A07778",
    x"30A0636B",
    x"30A04F5F",
    x"30A03B57",
    x"30A02751",
    x"30A0134D",
    x"309FFF4C",
    x"309FEB4D",
    x"309FD751",
    x"309FC357",
    x"309FAF60",
    x"309F9B6B",
    x"309F8779",
    x"309F7389",
    x"309F5F9C",
    x"309F4BB2",
    x"309F37C9",
    x"309F23E4",
    x"309F1000",
    x"309EFC20",
    x"309EE841",
    x"309ED466",
    x"309EC08C",
    x"309EACB5",
    x"309E98E1",
    x"309E850F",
    x"309E7140",
    x"309E5D73",
    x"309E49A8",
    x"309E35E0",
    x"309E221B",
    x"309E0E58",
    x"309DFA97",
    x"309DE6D9",
    x"309DD31E",
    x"309DBF65",
    x"309DABAE",
    x"309D97FA",
    x"309D8448",
    x"309D7099",
    x"309D5CEC",
    x"309D4941",
    x"309D3599",
    x"309D21F4",
    x"309D0E51",
    x"309CFAB0",
    x"309CE712",
    x"309CD377",
    x"309CBFDD",
    x"309CAC47",
    x"309C98B2",
    x"309C8520",
    x"309C7191",
    x"309C5E04",
    x"309C4A79",
    x"309C36F1",
    x"309C236C",
    x"309C0FE9",
    x"309BFC68",
    x"309BE8E9",
    x"309BD56E",
    x"309BC1F4",
    x"309BAE7D",
    x"309B9B08",
    x"309B8796",
    x"309B7427",
    x"309B60B9",
    x"309B4D4E",
    x"309B39E6",
    x"309B2680",
    x"309B131C",
    x"309AFFBB",
    x"309AEC5C",
    x"309AD900",
    x"309AC5A6",
    x"309AB24F",
    x"309A9EFA",
    x"309A8BA7",
    x"309A7857",
    x"309A6509",
    x"309A51BD",
    x"309A3E74",
    x"309A2B2E",
    x"309A17EA",
    x"309A04A8",
    x"3099F168",
    x"3099DE2B",
    x"3099CAF1",
    x"3099B7B9",
    x"3099A483",
    x"30999150",
    x"30997E1F",
    x"30996AF0",
    x"309957C4",
    x"3099449A",
    x"30993173",
    x"30991E4E",
    x"30990B2B",
    x"3098F80B",
    x"3098E4ED",
    x"3098D1D2",
    x"3098BEB9",
    x"3098ABA2",
    x"3098988E",
    x"3098857C",
    x"3098726C",
    x"30985F5F",
    x"30984C55",
    x"3098394C",
    x"30982646",
    x"30981343",
    x"30980041",
    x"3097ED43",
    x"3097DA46",
    x"3097C74C",
    x"3097B454",
    x"3097A15F",
    x"30978E6C",
    x"30977B7B",
    x"3097688D",
    x"309755A1",
    x"309742B8",
    x"30972FD0",
    x"30971CEC",
    x"30970A09",
    x"3096F729",
    x"3096E44B",
    x"3096D170",
    x"3096BE97",
    x"3096ABC0",
    x"309698EC",
    x"3096861A",
    x"3096734B",
    x"3096607D",
    x"30964DB3",
    x"30963AEA",
    x"30962824",
    x"30961560",
    x"3096029E",
    x"3095EFDF",
    x"3095DD22",
    x"3095CA68",
    x"3095B7B0",
    x"3095A4FA",
    x"30959247",
    x"30957F96",
    x"30956CE7",
    x"30955A3A",
    x"30954790",
    x"309534E8",
    x"30952243",
    x"30950FA0",
    x"3094FCFF",
    x"3094EA61",
    x"3094D7C4",
    x"3094C52B",
    x"3094B293",
    x"30949FFE",
    x"30948D6B",
    x"30947ADB",
    x"3094684C",
    x"309455C1",
    x"30944337",
    x"309430B0",
    x"30941E2B",
    x"30940BA8",
    x"3093F928",
    x"3093E6AA",
    x"3093D42E",
    x"3093C1B5",
    x"3093AF3E",
    x"30939CC9",
    x"30938A57",
    x"309377E6",
    x"30936579",
    x"3093530D",
    x"309340A4",
    x"30932E3D",
    x"30931BD8",
    x"30930976",
    x"3092F716",
    x"3092E4B8",
    x"3092D25D",
    x"3092C004",
    x"3092ADAD",
    x"30929B58",
    x"30928906",
    x"309276B6",
    x"30926468",
    x"3092521D",
    x"30923FD4",
    x"30922D8D",
    x"30921B48",
    x"30920906",
    x"3091F6C6",
    x"3091E488",
    x"3091D24D",
    x"3091C014",
    x"3091ADDD",
    x"30919BA8",
    x"30918976",
    x"30917746",
    x"30916518",
    x"309152ED",
    x"309140C3",
    x"30912E9D",
    x"30911C78",
    x"30910A55",
    x"3090F835",
    x"3090E617",
    x"3090D3FC",
    x"3090C1E2",
    x"3090AFCB",
    x"30909DB6",
    x"30908BA4",
    x"30907993",
    x"30906785",
    x"3090557A",
    x"30904370",
    x"30903169",
    x"30901F64",
    x"30900D61",
    x"308FFB60",
    x"308FE962",
    x"308FD766",
    x"308FC56C",
    x"308FB375",
    x"308FA17F",
    x"308F8F8C",
    x"308F7D9B",
    x"308F6BAD",
    x"308F59C1",
    x"308F47D6",
    x"308F35EF",
    x"308F2409",
    x"308F1226",
    x"308F0044",
    x"308EEE66",
    x"308EDC89",
    x"308ECAAE",
    x"308EB8D6",
    x"308EA700",
    x"308E952C",
    x"308E835B",
    x"308E718C",
    x"308E5FBE",
    x"308E4DF4",
    x"308E3C2B",
    x"308E2A65",
    x"308E18A0",
    x"308E06DE",
    x"308DF51F",
    x"308DE361",
    x"308DD1A6",
    x"308DBFED",
    x"308DAE36",
    x"308D9C81",
    x"308D8ACF",
    x"308D791E",
    x"308D6770",
    x"308D55C5",
    x"308D441B",
    x"308D3274",
    x"308D20CE",
    x"308D0F2B",
    x"308CFD8B",
    x"308CEBEC",
    x"308CDA50",
    x"308CC8B5",
    x"308CB71D",
    x"308CA588",
    x"308C93F4",
    x"308C8263",
    x"308C70D3",
    x"308C5F46",
    x"308C4DBC",
    x"308C3C33",
    x"308C2AAD",
    x"308C1928",
    x"308C07A6",
    x"308BF626",
    x"308BE4A9",
    x"308BD32D",
    x"308BC1B4",
    x"308BB03D",
    x"308B9EC8",
    x"308B8D55",
    x"308B7BE5",
    x"308B6A76",
    x"308B590A",
    x"308B47A0",
    x"308B3638",
    x"308B24D2",
    x"308B136F",
    x"308B020D",
    x"308AF0AE",
    x"308ADF51",
    x"308ACDF6",
    x"308ABC9E",
    x"308AAB47",
    x"308A99F3",
    x"308A88A1",
    x"308A7751",
    x"308A6603",
    x"308A54B7",
    x"308A436E",
    x"308A3226",
    x"308A20E1",
    x"308A0F9E",
    x"3089FE5D",
    x"3089ED1F",
    x"3089DBE2",
    x"3089CAA8",
    x"3089B96F",
    x"3089A839",
    x"30899705",
    x"308985D4",
    x"308974A4",
    x"30896376",
    x"3089524B",
    x"30894122",
    x"30892FFB",
    x"30891ED6",
    x"30890DB3",
    x"3088FC92",
    x"3088EB74",
    x"3088DA58",
    x"3088C93D",
    x"3088B825",
    x"3088A70F",
    x"308895FC",
    x"308884EA",
    x"308873DA",
    x"308862CD",
    x"308851C2",
    x"308840B8",
    x"30882FB1",
    x"30881EAC",
    x"30880DAA",
    x"3087FCA9",
    x"3087EBAB",
    x"3087DAAE",
    x"3087C9B4",
    x"3087B8BC",
    x"3087A7C6",
    x"308796D2",
    x"308785E0",
    x"308774F0",
    x"30876403",
    x"30875317",
    x"3087422E",
    x"30873147",
    x"30872062",
    x"30870F7F",
    x"3086FE9E",
    x"3086EDBF",
    x"3086DCE2",
    x"3086CC08",
    x"3086BB2F",
    x"3086AA59",
    x"30869985",
    x"308688B3",
    x"308677E3",
    x"30866715",
    x"30865649",
    x"3086457F",
    x"308634B7",
    x"308623F2",
    x"3086132E",
    x"3086026D",
    x"3085F1AE",
    x"3085E0F1",
    x"3085D036",
    x"3085BF7D",
    x"3085AEC6",
    x"30859E11",
    x"30858D5E",
    x"30857CAE",
    x"30856BFF",
    x"30855B53",
    x"30854AA8",
    x"30853A00",
    x"3085295A",
    x"308518B6",
    x"30850814",
    x"3084F774",
    x"3084E6D6",
    x"3084D63A",
    x"3084C5A0",
    x"3084B508",
    x"3084A473",
    x"308493DF",
    x"3084834E",
    x"308472BF",
    x"30846231",
    x"308451A6",
    x"3084411D",
    x"30843096",
    x"30842011",
    x"30840F8E",
    x"3083FF0D",
    x"3083EE8E",
    x"3083DE11",
    x"3083CD96",
    x"3083BD1E",
    x"3083ACA7",
    x"30839C33",
    x"30838BC0",
    x"30837B50",
    x"30836AE1",
    x"30835A75",
    x"30834A0B",
    x"308339A2",
    x"3083293C",
    x"308318D8",
    x"30830876",
    x"3082F816",
    x"3082E7B8",
    x"3082D75C",
    x"3082C702",
    x"3082B6AA",
    x"3082A654",
    x"30829601",
    x"308285AF",
    x"3082755F",
    x"30826512",
    x"308254C6",
    x"3082447C",
    x"30823435",
    x"308223EF",
    x"308213AC",
    x"3082036A",
    x"3081F32B",
    x"3081E2EE",
    x"3081D2B2",
    x"3081C279",
    x"3081B242",
    x"3081A20C",
    x"308191D9",
    x"308181A8",
    x"30817179",
    x"3081614C",
    x"30815120",
    x"308140F7",
    x"308130D0",
    x"308120AB",
    x"30811088",
    x"30810067",
    x"3080F048",
    x"3080E02B",
    x"3080D010",
    x"3080BFF7",
    x"3080AFE0",
    x"30809FCB",
    x"30808FB8",
    x"30807FA7",
    x"30806F98",
    x"30805F8B",
    x"30804F80",
    x"30803F77",
    x"30802F70",
    x"30801F6B",
    x"30800F68",
    x"307FFECF",
    x"307FDED1",
    x"307FBED7",
    x"307F9EE1",
    x"307F7EF0",
    x"307F5F02",
    x"307F3F18",
    x"307F1F32",
    x"307EFF50",
    x"307EDF72",
    x"307EBF98",
    x"307E9FC2",
    x"307E7FF0",
    x"307E6022",
    x"307E4058",
    x"307E2092",
    x"307E00D0",
    x"307DE112",
    x"307DC158",
    x"307DA1A2",
    x"307D81EF",
    x"307D6241",
    x"307D4297",
    x"307D22F1",
    x"307D034E",
    x"307CE3B0",
    x"307CC415",
    x"307CA47F",
    x"307C84EC",
    x"307C655D",
    x"307C45D3",
    x"307C264C",
    x"307C06C9",
    x"307BE74A",
    x"307BC7CF",
    x"307BA858",
    x"307B88E5",
    x"307B6976",
    x"307B4A0B",
    x"307B2AA4",
    x"307B0B40",
    x"307AEBE1",
    x"307ACC85",
    x"307AAD2E",
    x"307A8DDA",
    x"307A6E8A",
    x"307A4F3E",
    x"307A2FF6",
    x"307A10B2",
    x"3079F172",
    x"3079D236",
    x"3079B2FE",
    x"307993C9",
    x"30797499",
    x"3079556C",
    x"30793643",
    x"3079171E",
    x"3078F7FE",
    x"3078D8E0",
    x"3078B9C7",
    x"30789AB2",
    x"30787BA1",
    x"30785C93",
    x"30783D8A",
    x"30781E84",
    x"3077FF82",
    x"3077E084",
    x"3077C18A",
    x"3077A293",
    x"307783A1",
    x"307764B3",
    x"307745C8",
    x"307726E1",
    x"307707FE",
    x"3076E91F",
    x"3076CA44",
    x"3076AB6D",
    x"30768C99",
    x"30766DC9",
    x"30764EFE",
    x"30763036",
    x"30761172",
    x"3075F2B1",
    x"3075D3F5",
    x"3075B53C",
    x"30759688",
    x"307577D7",
    x"3075592A",
    x"30753A80",
    x"30751BDB",
    x"3074FD39",
    x"3074DE9C",
    x"3074C002",
    x"3074A16C",
    x"307482D9",
    x"3074644B",
    x"307445C0",
    x"3074273A",
    x"307408B7",
    x"3073EA37",
    x"3073CBBC",
    x"3073AD44",
    x"30738ED1",
    x"30737061",
    x"307351F5",
    x"3073338C",
    x"30731528",
    x"3072F6C7",
    x"3072D86A",
    x"3072BA11",
    x"30729BBB",
    x"30727D6A",
    x"30725F1C",
    x"307240D2",
    x"3072228C",
    x"30720449",
    x"3071E60B",
    x"3071C7D0",
    x"3071A999",
    x"30718B66",
    x"30716D36",
    x"30714F0A",
    x"307130E2",
    x"307112BE",
    x"3070F49E",
    x"3070D681",
    x"3070B868",
    x"30709A53",
    x"30707C41",
    x"30705E34",
    x"3070402A",
    x"30702224",
    x"30700421",
    x"306FE623",
    x"306FC828",
    x"306FAA31",
    x"306F8C3D",
    x"306F6E4E",
    x"306F5062",
    x"306F3279",
    x"306F1495",
    x"306EF6B4",
    x"306ED8D7",
    x"306EBAFE",
    x"306E9D29",
    x"306E7F57",
    x"306E6189",
    x"306E43BE",
    x"306E25F8",
    x"306E0835",
    x"306DEA76",
    x"306DCCBA",
    x"306DAF03",
    x"306D914F",
    x"306D739E",
    x"306D55F2",
    x"306D3849",
    x"306D1AA4",
    x"306CFD02",
    x"306CDF64",
    x"306CC1CA",
    x"306CA434",
    x"306C86A1",
    x"306C6912",
    x"306C4B87",
    x"306C2DFF",
    x"306C107B",
    x"306BF2FB",
    x"306BD57F",
    x"306BB806",
    x"306B9A91",
    x"306B7D1F",
    x"306B5FB1",
    x"306B4247",
    x"306B24E1",
    x"306B077E",
    x"306AEA1F",
    x"306ACCC4",
    x"306AAF6C",
    x"306A9218",
    x"306A74C7",
    x"306A577A",
    x"306A3A31",
    x"306A1CEC",
    x"3069FFAA",
    x"3069E26C",
    x"3069C532",
    x"3069A7FB",
    x"30698AC8",
    x"30696D98",
    x"3069506C",
    x"30693344",
    x"3069161F",
    x"3068F8FE",
    x"3068DBE1",
    x"3068BEC7",
    x"3068A1B1",
    x"3068849F",
    x"30686790",
    x"30684A85",
    x"30682D7E",
    x"3068107A",
    x"3067F379",
    x"3067D67D",
    x"3067B984",
    x"30679C8E",
    x"30677F9D",
    x"306762AF",
    x"306745C4",
    x"306728DD",
    x"30670BFA",
    x"3066EF1A",
    x"3066D23E",
    x"3066B566",
    x"30669891",
    x"30667BBF",
    x"30665EF2",
    x"30664228",
    x"30662561",
    x"3066089E",
    x"3065EBDF",
    x"3065CF23",
    x"3065B26B",
    x"306595B7",
    x"30657906",
    x"30655C59",
    x"30653FAF",
    x"30652309",
    x"30650666",
    x"3064E9C7",
    x"3064CD2C",
    x"3064B094",
    x"306493FF",
    x"3064776F",
    x"30645AE2",
    x"30643E58",
    x"306421D2",
    x"30640550",
    x"3063E8D1",
    x"3063CC55",
    x"3063AFDE",
    x"30639369",
    x"306376F9",
    x"30635A8C",
    x"30633E22",
    x"306321BC",
    x"3063055A",
    x"3062E8FB",
    x"3062CC9F",
    x"3062B048",
    x"306293F3",
    x"306277A3",
    x"30625B55",
    x"30623F0C",
    x"306222C6",
    x"30620683",
    x"3061EA44",
    x"3061CE09",
    x"3061B1D1",
    x"3061959C",
    x"3061796B",
    x"30615D3E",
    x"30614114",
    x"306124ED",
    x"306108CB",
    x"3060ECAB",
    x"3060D08F",
    x"3060B477",
    x"30609862",
    x"30607C51",
    x"30606043",
    x"30604439",
    x"30602832",
    x"30600C2F",
    x"305FF02F",
    x"305FD433",
    x"305FB83A",
    x"305F9C45",
    x"305F8053",
    x"305F6465",
    x"305F487A",
    x"305F2C93",
    x"305F10AF",
    x"305EF4CE",
    x"305ED8F2",
    x"305EBD18",
    x"305EA142",
    x"305E8570",
    x"305E69A1",
    x"305E4DD5",
    x"305E320D",
    x"305E1649",
    x"305DFA88",
    x"305DDECA",
    x"305DC310",
    x"305DA75A",
    x"305D8BA6",
    x"305D6FF7",
    x"305D544A",
    x"305D38A2",
    x"305D1CFC",
    x"305D015A",
    x"305CE5BC",
    x"305CCA21",
    x"305CAE89",
    x"305C92F5",
    x"305C7765",
    x"305C5BD7",
    x"305C404E",
    x"305C24C7",
    x"305C0944",
    x"305BEDC5",
    x"305BD249",
    x"305BB6D0",
    x"305B9B5B",
    x"305B7FEA",
    x"305B647B",
    x"305B4910",
    x"305B2DA9",
    x"305B1245",
    x"305AF6E4",
    x"305ADB87",
    x"305AC02E",
    x"305AA4D7",
    x"305A8984",
    x"305A6E35",
    x"305A52E9",
    x"305A37A0",
    x"305A1C5B",
    x"305A0119",
    x"3059E5DB",
    x"3059CAA0",
    x"3059AF68",
    x"30599434",
    x"30597903",
    x"30595DD6",
    x"305942AB",
    x"30592785",
    x"30590C62",
    x"3058F142",
    x"3058D625",
    x"3058BB0C",
    x"30589FF7",
    x"305884E4",
    x"305869D5",
    x"30584ECA",
    x"305833C2",
    x"305818BD",
    x"3057FDBB",
    x"3057E2BD",
    x"3057C7C3",
    x"3057ACCB",
    x"305791D8",
    x"305776E7",
    x"30575BFA",
    x"30574110",
    x"3057262A",
    x"30570B46",
    x"3056F067",
    x"3056D58A",
    x"3056BAB1",
    x"30569FDC",
    x"30568509",
    x"30566A3A",
    x"30564F6F",
    x"305634A7",
    x"305619E2",
    x"3055FF20",
    x"3055E462",
    x"3055C9A7",
    x"3055AEEF",
    x"3055943B",
    x"3055798A",
    x"30555EDD",
    x"30554433",
    x"3055298C",
    x"30550EE8",
    x"3054F448",
    x"3054D9AB",
    x"3054BF12",
    x"3054A47B",
    x"305489E9",
    x"30546F59",
    x"305454CD",
    x"30543A44",
    x"30541FBE",
    x"3054053C",
    x"3053EABD",
    x"3053D041",
    x"3053B5C9",
    x"30539B54",
    x"305380E2",
    x"30536673",
    x"30534C08",
    x"305331A0",
    x"3053173C",
    x"3052FCDB",
    x"3052E27D",
    x"3052C822",
    x"3052ADCB",
    x"30529377",
    x"30527926",
    x"30525ED8",
    x"3052448E",
    x"30522A47",
    x"30521004",
    x"3051F5C3",
    x"3051DB86",
    x"3051C14C",
    x"3051A716",
    x"30518CE3",
    x"305172B3",
    x"30515886",
    x"30513E5C",
    x"30512436",
    x"30510A13",
    x"3050EFF4",
    x"3050D5D7",
    x"3050BBBE",
    x"3050A1A8",
    x"30508796",
    x"30506D87",
    x"3050537A",
    x"30503972",
    x"30501F6C",
    x"3050056A",
    x"304FEB6B",
    x"304FD16F",
    x"304FB776",
    x"304F9D81",
    x"304F838F",
    x"304F69A0",
    x"304F4FB5",
    x"304F35CC",
    x"304F1BE7",
    x"304F0205",
    x"304EE827",
    x"304ECE4B",
    x"304EB473",
    x"304E9A9E",
    x"304E80CC",
    x"304E66FE",
    x"304E4D33",
    x"304E336B",
    x"304E19A6",
    x"304DFFE4",
    x"304DE626",
    x"304DCC6B",
    x"304DB2B3",
    x"304D98FE",
    x"304D7F4C",
    x"304D659E",
    x"304D4BF3",
    x"304D324B",
    x"304D18A7",
    x"304CFF05",
    x"304CE567",
    x"304CCBCC",
    x"304CB234",
    x"304C989F",
    x"304C7F0E",
    x"304C657F",
    x"304C4BF4",
    x"304C326C",
    x"304C18E8",
    x"304BFF66",
    x"304BE5E8",
    x"304BCC6D",
    x"304BB2F5",
    x"304B9980",
    x"304B800E",
    x"304B66A0",
    x"304B4D35",
    x"304B33CD",
    x"304B1A68",
    x"304B0106",
    x"304AE7A7",
    x"304ACE4C",
    x"304AB4F4",
    x"304A9B9F",
    x"304A824D",
    x"304A68FE",
    x"304A4FB3",
    x"304A366A",
    x"304A1D25",
    x"304A03E3",
    x"3049EAA4",
    x"3049D168",
    x"3049B830",
    x"30499EFA",
    x"304985C8",
    x"30496C99",
    x"3049536D",
    x"30493A44",
    x"3049211E",
    x"304907FC",
    x"3048EEDC",
    x"3048D5C0",
    x"3048BCA7",
    x"3048A391",
    x"30488A7E",
    x"3048716E",
    x"30485862",
    x"30483F58",
    x"30482652",
    x"30480D4F",
    x"3047F44F",
    x"3047DB52",
    x"3047C258",
    x"3047A961",
    x"3047906D",
    x"3047777D",
    x"30475E8F",
    x"304745A5",
    x"30472CBE",
    x"304713DA",
    x"3046FAF9",
    x"3046E21B",
    x"3046C941",
    x"3046B069",
    x"30469794",
    x"30467EC3",
    x"304665F5",
    x"30464D2A",
    x"30463461",
    x"30461B9C",
    x"304602DB",
    x"3045EA1C",
    x"3045D160",
    x"3045B8A7",
    x"30459FF2",
    x"3045873F",
    x"30456E90",
    x"304555E4",
    x"30453D3B",
    x"30452494",
    x"30450BF1",
    x"3044F351",
    x"3044DAB5",
    x"3044C21B",
    x"3044A984",
    x"304490F0",
    x"30447860",
    x"30445FD2",
    x"30444748",
    x"30442EC1",
    x"3044163C",
    x"3043FDBB",
    x"3043E53D",
    x"3043CCC2",
    x"3043B44A",
    x"30439BD5",
    x"30438363",
    x"30436AF4",
    x"30435288",
    x"30433A1F",
    x"304321B9",
    x"30430957",
    x"3042F0F7",
    x"3042D89A",
    x"3042C041",
    x"3042A7EA",
    x"30428F97",
    x"30427746",
    x"30425EF9",
    x"304246AF",
    x"30422E67",
    x"30421623",
    x"3041FDE2",
    x"3041E5A4",
    x"3041CD68",
    x"3041B530",
    x"30419CFB",
    x"304184C9",
    x"30416C9A",
    x"3041546E",
    x"30413C45",
    x"3041241F",
    x"30410BFC",
    x"3040F3DC",
    x"3040DBBF",
    x"3040C3A5",
    x"3040AB8E",
    x"3040937A",
    x"30407B69",
    x"3040635B",
    x"30404B50",
    x"30403348",
    x"30401B43",
    x"30400342",
    x"303FEB43",
    x"303FD347",
    x"303FBB4E",
    x"303FA358",
    x"303F8B65",
    x"303F7375",
    x"303F5B88",
    x"303F439E",
    x"303F2BB7",
    x"303F13D3",
    x"303EFBF2",
    x"303EE414",
    x"303ECC39",
    x"303EB461",
    x"303E9C8C",
    x"303E84BA",
    x"303E6CEB",
    x"303E551F",
    x"303E3D56",
    x"303E258F",
    x"303E0DCC",
    x"303DF60C",
    x"303DDE4F",
    x"303DC694",
    x"303DAEDD",
    x"303D9729",
    x"303D7F77",
    x"303D67C9",
    x"303D501D",
    x"303D3875",
    x"303D20CF",
    x"303D092D",
    x"303CF18D",
    x"303CD9F0",
    x"303CC256",
    x"303CAAC0",
    x"303C932C",
    x"303C7B9B",
    x"303C640D",
    x"303C4C82",
    x"303C34FA",
    x"303C1D75",
    x"303C05F2",
    x"303BEE73",
    x"303BD6F7",
    x"303BBF7D",
    x"303BA807",
    x"303B9093",
    x"303B7923",
    x"303B61B5",
    x"303B4A4A",
    x"303B32E3",
    x"303B1B7E",
    x"303B041C",
    x"303AECBD",
    x"303AD560",
    x"303ABE07",
    x"303AA6B1",
    x"303A8F5E",
    x"303A780D",
    x"303A60C0",
    x"303A4975",
    x"303A322D",
    x"303A1AE8",
    x"303A03A6",
    x"3039EC67",
    x"3039D52B",
    x"3039BDF2",
    x"3039A6BC",
    x"30398F88",
    x"30397858",
    x"3039612A",
    x"30394A00",
    x"303932D8",
    x"30391BB3",
    x"30390491",
    x"3038ED72",
    x"3038D656",
    x"3038BF3C",
    x"3038A826",
    x"30389112",
    x"30387A02",
    x"303862F4",
    x"30384BE9",
    x"303834E1",
    x"30381DDC",
    x"303806D9",
    x"3037EFDA",
    x"3037D8DD",
    x"3037C1E4",
    x"3037AAED",
    x"303793F9",
    x"30377D08",
    x"3037661A",
    x"30374F2E",
    x"30373846",
    x"30372160",
    x"30370A7E",
    x"3036F39E",
    x"3036DCC1",
    x"3036C5E6",
    x"3036AF0F",
    x"3036983B",
    x"30368169",
    x"30366A9A",
    x"303653CE",
    x"30363D05",
    x"3036263F",
    x"30360F7C",
    x"3035F8BB",
    x"3035E1FE",
    x"3035CB43",
    x"3035B48B",
    x"30359DD6",
    x"30358723",
    x"30357074",
    x"303559C7",
    x"3035431D",
    x"30352C76",
    x"303515D2",
    x"3034FF31",
    x"3034E893",
    x"3034D1F7",
    x"3034BB5E",
    x"3034A4C8",
    x"30348E35",
    x"303477A4",
    x"30346117",
    x"30344A8C",
    x"30343404",
    x"30341D7F",
    x"303406FD",
    x"3033F07D",
    x"3033DA01",
    x"3033C387",
    x"3033AD10",
    x"3033969C",
    x"3033802A",
    x"303369BC",
    x"30335350",
    x"30333CE7",
    x"30332681",
    x"3033101D",
    x"3032F9BD",
    x"3032E35F",
    x"3032CD04",
    x"3032B6AB",
    x"3032A056",
    x"30328A03",
    x"303273B4",
    x"30325D66",
    x"3032471C",
    x"303230D5",
    x"30321A90",
    x"3032044E",
    x"3031EE0F",
    x"3031D7D3",
    x"3031C199",
    x"3031AB62",
    x"3031952E",
    x"30317EFD",
    x"303168CE",
    x"303152A3",
    x"30313C7A",
    x"30312654",
    x"30311030",
    x"3030FA0F",
    x"3030E3F2",
    x"3030CDD6",
    x"3030B7BE",
    x"3030A1A9",
    x"30308B96",
    x"30307586",
    x"30305F78",
    x"3030496E",
    x"30303366",
    x"30301D61",
    x"3030075F",
    x"302FF15F",
    x"302FDB62",
    x"302FC568",
    x"302FAF71",
    x"302F997C",
    x"302F838B",
    x"302F6D9B",
    x"302F57AF",
    x"302F41C6",
    x"302F2BDF",
    x"302F15FB",
    x"302F0019",
    x"302EEA3B",
    x"302ED45F",
    x"302EBE85",
    x"302EA8AF",
    x"302E92DB",
    x"302E7D0A",
    x"302E673C",
    x"302E5171",
    x"302E3BA8",
    x"302E25E2",
    x"302E101E",
    x"302DFA5E",
    x"302DE4A0",
    x"302DCEE4",
    x"302DB92C",
    x"302DA376",
    x"302D8DC3",
    x"302D7813",
    x"302D6265",
    x"302D4CBA",
    x"302D3712",
    x"302D216C",
    x"302D0BC9",
    x"302CF629",
    x"302CE08C",
    x"302CCAF1",
    x"302CB559",
    x"302C9FC4",
    x"302C8A31",
    x"302C74A1",
    x"302C5F14",
    x"302C498A",
    x"302C3402",
    x"302C1E7D",
    x"302C08FA",
    x"302BF37A",
    x"302BDDFD",
    x"302BC883",
    x"302BB30B",
    x"302B9D96",
    x"302B8824",
    x"302B72B4",
    x"302B5D47",
    x"302B47DD",
    x"302B3275",
    x"302B1D10",
    x"302B07AE",
    x"302AF24E",
    x"302ADCF1",
    x"302AC797",
    x"302AB23F",
    x"302A9CEA",
    x"302A8798",
    x"302A7248",
    x"302A5CFC",
    x"302A47B1",
    x"302A326A",
    x"302A1D25",
    x"302A07E2",
    x"3029F2A3",
    x"3029DD66",
    x"3029C82B",
    x"3029B2F4",
    x"30299DBF",
    x"3029888C",
    x"3029735C",
    x"30295E2F",
    x"30294905",
    x"302933DD",
    x"30291EB8",
    x"30290995",
    x"3028F476",
    x"3028DF58",
    x"3028CA3E",
    x"3028B526",
    x"3028A010",
    x"30288AFE",
    x"302875EE",
    x"302860E0",
    x"30284BD5",
    x"302836CD",
    x"302821C8",
    x"30280CC5",
    x"3027F7C5",
    x"3027E2C7",
    x"3027CDCC",
    x"3027B8D3",
    x"3027A3DE",
    x"30278EEA",
    x"302779FA",
    x"3027650C",
    x"30275021",
    x"30273B38",
    x"30272652",
    x"3027116E",
    x"3026FC8D",
    x"3026E7AF",
    x"3026D2D4",
    x"3026BDFB",
    x"3026A924",
    x"30269450",
    x"30267F7F",
    x"30266AB0",
    x"302655E4",
    x"3026411B",
    x"30262C54",
    x"30261790",
    x"302602CE",
    x"3025EE0F",
    x"3025D953",
    x"3025C499",
    x"3025AFE1",
    x"30259B2D",
    x"3025867B",
    x"302571CB",
    x"30255D1E",
    x"30254874",
    x"302533CC",
    x"30251F27",
    x"30250A84",
    x"3024F5E4",
    x"3024E147",
    x"3024CCAC",
    x"3024B814",
    x"3024A37E",
    x"30248EEB",
    x"30247A5A",
    x"302465CC",
    x"30245141",
    x"30243CB8",
    x"30242832",
    x"302413AE",
    x"3023FF2D",
    x"3023EAAE",
    x"3023D632",
    x"3023C1B9",
    x"3023AD42",
    x"302398CD",
    x"3023845B",
    x"30236FEC",
    x"30235B7F",
    x"30234715",
    x"302332AE",
    x"30231E49",
    x"302309E6",
    x"3022F586",
    x"3022E129",
    x"3022CCCE",
    x"3022B875",
    x"3022A420",
    x"30228FCC",
    x"30227B7C",
    x"3022672E",
    x"302252E2",
    x"30223E99",
    x"30222A52",
    x"3022160E",
    x"302201CD",
    x"3021ED8E",
    x"3021D951",
    x"3021C518",
    x"3021B0E0",
    x"30219CAB",
    x"30218879",
    x"30217449",
    x"3021601C",
    x"30214BF1",
    x"302137C9",
    x"302123A3",
    x"30210F80",
    x"3020FB5F",
    x"3020E741",
    x"3020D326",
    x"3020BF0C",
    x"3020AAF6",
    x"302096E2",
    x"302082D0",
    x"30206EC1",
    x"30205AB4",
    x"302046AA",
    x"302032A3",
    x"30201E9E",
    x"30200A9B",
    x"301FF69B",
    x"301FE29D",
    x"301FCEA2",
    x"301FBAAA",
    x"301FA6B4",
    x"301F92C0",
    x"301F7ECF",
    x"301F6AE0",
    x"301F56F4",
    x"301F430B",
    x"301F2F23",
    x"301F1B3F",
    x"301F075D",
    x"301EF37D",
    x"301EDFA0",
    x"301ECBC5",
    x"301EB7ED",
    x"301EA417",
    x"301E9044",
    x"301E7C73",
    x"301E68A5",
    x"301E54D9",
    x"301E410F",
    x"301E2D49",
    x"301E1984",
    x"301E05C2",
    x"301DF203",
    x"301DDE46",
    x"301DCA8B",
    x"301DB6D3",
    x"301DA31D",
    x"301D8F6A",
    x"301D7BBA",
    x"301D680B",
    x"301D5460",
    x"301D40B6",
    x"301D2D0F",
    x"301D196B",
    x"301D05C9",
    x"301CF22A",
    x"301CDE8C",
    x"301CCAF2",
    x"301CB75A",
    x"301CA3C4",
    x"301C9031",
    x"301C7CA0",
    x"301C6912",
    x"301C5586",
    x"301C41FC",
    x"301C2E75",
    x"301C1AF1",
    x"301C076F",
    x"301BF3EF",
    x"301BE072",
    x"301BCCF7",
    x"301BB97E",
    x"301BA608",
    x"301B9295",
    x"301B7F24",
    x"301B6BB5",
    x"301B5849",
    x"301B44DF",
    x"301B3178",
    x"301B1E13",
    x"301B0AB0",
    x"301AF750",
    x"301AE3F2",
    x"301AD097",
    x"301ABD3E",
    x"301AA9E8",
    x"301A9694",
    x"301A8342",
    x"301A6FF3",
    x"301A5CA6",
    x"301A495C",
    x"301A3614",
    x"301A22CE",
    x"301A0F8B",
    x"3019FC4A",
    x"3019E90C",
    x"3019D5D0",
    x"3019C296",
    x"3019AF5F",
    x"30199C2B",
    x"301988F8",
    x"301975C8",
    x"3019629B",
    x"30194F70",
    x"30193C47",
    x"30192921",
    x"301915FD",
    x"301902DB",
    x"3018EFBC",
    x"3018DC9F",
    x"3018C985",
    x"3018B66D",
    x"3018A357",
    x"30189044",
    x"30187D33",
    x"30186A25",
    x"30185719",
    x"3018440F",
    x"30183108",
    x"30181E03",
    x"30180B00",
    x"3017F800",
    x"3017E502",
    x"3017D207",
    x"3017BF0E",
    x"3017AC17",
    x"30179923",
    x"30178631",
    x"30177341",
    x"30176054",
    x"30174D69",
    x"30173A80",
    x"3017279A",
    x"301714B6",
    x"301701D5",
    x"3016EEF6",
    x"3016DC19",
    x"3016C93F",
    x"3016B667",
    x"3016A391",
    x"301690BE",
    x"30167DED",
    x"30166B1F",
    x"30165852",
    x"30164589",
    x"301632C1",
    x"30161FFC",
    x"30160D39",
    x"3015FA79",
    x"3015E7BA",
    x"3015D4FF",
    x"3015C245",
    x"3015AF8E",
    x"30159CD9",
    x"30158A27",
    x"30157777",
    x"301564C9",
    x"3015521E",
    x"30153F74",
    x"30152CCE",
    x"30151A29",
    x"30150787",
    x"3014F4E7",
    x"3014E24A",
    x"3014CFAF",
    x"3014BD16",
    x"3014AA80",
    x"301497EB",
    x"3014855A",
    x"301472CA",
    x"3014603D",
    x"30144DB2",
    x"30143B29",
    x"301428A3",
    x"3014161F",
    x"3014039E",
    x"3013F11E",
    x"3013DEA1",
    x"3013CC27",
    x"3013B9AE",
    x"3013A738",
    x"301394C5",
    x"30138253",
    x"30136FE4",
    x"30135D77",
    x"30134B0D",
    x"301338A4",
    x"3013263E",
    x"301313DB",
    x"30130179",
    x"3012EF1A",
    x"3012DCBE",
    x"3012CA63",
    x"3012B80B",
    x"3012A5B5",
    x"30129362",
    x"30128110",
    x"30126EC1",
    x"30125C75",
    x"30124A2A",
    x"301237E2",
    x"3012259C",
    x"30121359",
    x"30120117",
    x"3011EED8",
    x"3011DC9C",
    x"3011CA61",
    x"3011B829",
    x"3011A5F3",
    x"301193C0",
    x"3011818E",
    x"30116F5F",
    x"30115D33",
    x"30114B08",
    x"301138E0",
    x"301126BA",
    x"30111496",
    x"30110275",
    x"3010F055",
    x"3010DE39",
    x"3010CC1E",
    x"3010BA06",
    x"3010A7EF",
    x"301095DC",
    x"301083CA",
    x"301071BB",
    x"30105FAD",
    x"30104DA3",
    x"30103B9A",
    x"30102994",
    x"30101790",
    x"3010058E",
    x"300FF38E",
    x"300FE191",
    x"300FCF96",
    x"300FBD9D",
    x"300FABA7",
    x"300F99B2",
    x"300F87C0",
    x"300F75D0",
    x"300F63E3",
    x"300F51F7",
    x"300F400E",
    x"300F2E27",
    x"300F1C43",
    x"300F0A60",
    x"300EF880",
    x"300EE6A2",
    x"300ED4C6",
    x"300EC2ED",
    x"300EB116",
    x"300E9F41",
    x"300E8D6E",
    x"300E7B9D",
    x"300E69CF",
    x"300E5803",
    x"300E4639",
    x"300E3471",
    x"300E22AC",
    x"300E10E9",
    x"300DFF28",
    x"300DED69",
    x"300DDBAC",
    x"300DC9F2",
    x"300DB83A",
    x"300DA684",
    x"300D94D0",
    x"300D831F",
    x"300D716F",
    x"300D5FC2",
    x"300D4E17",
    x"300D3C6F",
    x"300D2AC8",
    x"300D1924",
    x"300D0782",
    x"300CF5E2",
    x"300CE444",
    x"300CD2A9",
    x"300CC110",
    x"300CAF79",
    x"300C9DE4",
    x"300C8C51",
    x"300C7AC1",
    x"300C6933",
    x"300C57A7",
    x"300C461D",
    x"300C3495",
    x"300C2310",
    x"300C118C",
    x"300C000B",
    x"300BEE8C",
    x"300BDD10",
    x"300BCB95",
    x"300BBA1D",
    x"300BA8A6",
    x"300B9732",
    x"300B85C1",
    x"300B7451",
    x"300B62E4",
    x"300B5178",
    x"300B400F",
    x"300B2EA8",
    x"300B1D44",
    x"300B0BE1",
    x"300AFA81",
    x"300AE922",
    x"300AD7C6",
    x"300AC66C",
    x"300AB515",
    x"300AA3BF",
    x"300A926C",
    x"300A811B",
    x"300A6FCC",
    x"300A5E7F",
    x"300A4D34",
    x"300A3BEB",
    x"300A2AA5",
    x"300A1961",
    x"300A081F",
    x"3009F6DF",
    x"3009E5A1",
    x"3009D465",
    x"3009C32C",
    x"3009B1F4",
    x"3009A0BF",
    x"30098F8C",
    x"30097E5B",
    x"30096D2D",
    x"30095C00",
    x"30094AD6",
    x"300939AD",
    x"30092887",
    x"30091763",
    x"30090641",
    x"3008F522",
    x"3008E404",
    x"3008D2E9",
    x"3008C1CF",
    x"3008B0B8",
    x"30089FA3",
    x"30088E90",
    x"30087D80",
    x"30086C71",
    x"30085B64",
    x"30084A5A",
    x"30083952",
    x"3008284C",
    x"30081748",
    x"30080646",
    x"3007F546",
    x"3007E449",
    x"3007D34D",
    x"3007C254",
    x"3007B15D",
    x"3007A067",
    x"30078F74",
    x"30077E84",
    x"30076D95",
    x"30075CA8",
    x"30074BBE",
    x"30073AD5",
    x"300729EF",
    x"3007190B",
    x"30070829",
    x"3006F749",
    x"3006E66B",
    x"3006D58F",
    x"3006C4B5",
    x"3006B3DE",
    x"3006A309",
    x"30069235",
    x"30068164",
    x"30067095",
    x"30065FC8",
    x"30064EFD",
    x"30063E34",
    x"30062D6D",
    x"30061CA9",
    x"30060BE6",
    x"3005FB26",
    x"3005EA67",
    x"3005D9AB",
    x"3005C8F1",
    x"3005B839",
    x"3005A783",
    x"300596CF",
    x"3005861D",
    x"3005756D",
    x"300564C0",
    x"30055414",
    x"3005436B",
    x"300532C3",
    x"3005221E",
    x"3005117B",
    x"300500DA",
    x"3004F03B",
    x"3004DF9E",
    x"3004CF03",
    x"3004BE6A",
    x"3004ADD3",
    x"30049D3E",
    x"30048CAC",
    x"30047C1B",
    x"30046B8D",
    x"30045B00",
    x"30044A76",
    x"300439EE",
    x"30042968",
    x"300418E3",
    x"30040861",
    x"3003F7E1",
    x"3003E763",
    x"3003D6E8",
    x"3003C66E",
    x"3003B5F6",
    x"3003A580",
    x"3003950D",
    x"3003849B",
    x"3003742B",
    x"300363BE",
    x"30035352",
    x"300342E9",
    x"30033282",
    x"3003221C",
    x"300311B9",
    x"30030158",
    x"3002F0F9",
    x"3002E09C",
    x"3002D041",
    x"3002BFE8",
    x"3002AF91",
    x"30029F3C",
    x"30028EE9",
    x"30027E98",
    x"30026E49",
    x"30025DFD",
    x"30024DB2",
    x"30023D69",
    x"30022D22",
    x"30021CDE",
    x"30020C9B",
    x"3001FC5B",
    x"3001EC1C",
    x"3001DBE0",
    x"3001CBA5",
    x"3001BB6D",
    x"3001AB36",
    x"30019B02",
    x"30018AD0",
    x"30017A9F",
    x"30016A71",
    x"30015A45",
    x"30014A1A",
    x"300139F2",
    x"300129CC",
    x"300119A8",
    x"30010985",
    x"3000F965",
    x"3000E947",
    x"3000D92B",
    x"3000C911",
    x"3000B8F9",
    x"3000A8E3",
    x"300098CE",
    x"300088BC",
    x"300078AC",
    x"3000689E",
    x"30005892",
    x"30004888",
    x"30003880",
    x"3000287A",
    x"30001876",
    x"30000874",
    x"2FFFF0E7",
    x"2FFFD0EB",
    x"2FFFB0F3",
    x"2FFF90FF",
    x"2FFF710F",
    x"2FFF5123",
    x"2FFF313B",
    x"2FFF1157",
    x"2FFEF176",
    x"2FFED19A",
    x"2FFEB1C2",
    x"2FFE91EE",
    x"2FFE721D",
    x"2FFE5251",
    x"2FFE3289",
    x"2FFE12C5",
    x"2FFDF304",
    x"2FFDD348",
    x"2FFDB38F",
    x"2FFD93DB",
    x"2FFD742A",
    x"2FFD547E",
    x"2FFD34D5",
    x"2FFD1531",
    x"2FFCF590",
    x"2FFCD5F3",
    x"2FFCB65B",
    x"2FFC96C6",
    x"2FFC7735",
    x"2FFC57A8",
    x"2FFC381F",
    x"2FFC189A",
    x"2FFBF919",
    x"2FFBD99C",
    x"2FFBBA22",
    x"2FFB9AAD",
    x"2FFB7B3C",
    x"2FFB5BCE",
    x"2FFB3C65",
    x"2FFB1CFF",
    x"2FFAFD9D",
    x"2FFADE40",
    x"2FFABEE6",
    x"2FFA9F90",
    x"2FFA803E",
    x"2FFA60F0",
    x"2FFA41A6",
    x"2FFA2260",
    x"2FFA031D",
    x"2FF9E3DF",
    x"2FF9C4A4",
    x"2FF9A56E",
    x"2FF9863B",
    x"2FF9670C",
    x"2FF947E1",
    x"2FF928BA",
    x"2FF90997",
    x"2FF8EA78",
    x"2FF8CB5C",
    x"2FF8AC45",
    x"2FF88D31",
    x"2FF86E22",
    x"2FF84F16",
    x"2FF8300E",
    x"2FF8110A",
    x"2FF7F209",
    x"2FF7D30D",
    x"2FF7B415",
    x"2FF79520",
    x"2FF7762F",
    x"2FF75743",
    x"2FF7385A",
    x"2FF71975",
    x"2FF6FA93",
    x"2FF6DBB6",
    x"2FF6BCDC",
    x"2FF69E07",
    x"2FF67F35",
    x"2FF66067",
    x"2FF6419D",
    x"2FF622D6",
    x"2FF60414",
    x"2FF5E555",
    x"2FF5C69B",
    x"2FF5A7E4",
    x"2FF58931",
    x"2FF56A81",
    x"2FF54BD6",
    x"2FF52D2F",
    x"2FF50E8B",
    x"2FF4EFEB",
    x"2FF4D14F",
    x"2FF4B2B7",
    x"2FF49422",
    x"2FF47592",
    x"2FF45705",
    x"2FF4387C",
    x"2FF419F7",
    x"2FF3FB75",
    x"2FF3DCF8",
    x"2FF3BE7E",
    x"2FF3A008",
    x"2FF38196",
    x"2FF36328",
    x"2FF344BD",
    x"2FF32657",
    x"2FF307F4",
    x"2FF2E995",
    x"2FF2CB39",
    x"2FF2ACE2",
    x"2FF28E8E",
    x"2FF2703E",
    x"2FF251F2",
    x"2FF233AA",
    x"2FF21565",
    x"2FF1F724",
    x"2FF1D8E7",
    x"2FF1BAAE",
    x"2FF19C79",
    x"2FF17E47",
    x"2FF16019",
    x"2FF141EF",
    x"2FF123C9",
    x"2FF105A6",
    x"2FF0E787",
    x"2FF0C96C",
    x"2FF0AB55",
    x"2FF08D41",
    x"2FF06F31",
    x"2FF05125",
    x"2FF0331D",
    x"2FF01519",
    x"2FEFF718",
    x"2FEFD91B",
    x"2FEFBB22",
    x"2FEF9D2C",
    x"2FEF7F3A",
    x"2FEF614C",
    x"2FEF4362",
    x"2FEF257B",
    x"2FEF0799",
    x"2FEEE9BA",
    x"2FEECBDE",
    x"2FEEAE07",
    x"2FEE9033",
    x"2FEE7263",
    x"2FEE5496",
    x"2FEE36CD",
    x"2FEE1908",
    x"2FEDFB47",
    x"2FEDDD8A",
    x"2FEDBFD0",
    x"2FEDA21A",
    x"2FED8467",
    x"2FED66B9",
    x"2FED490E",
    x"2FED2B66",
    x"2FED0DC3",
    x"2FECF023",
    x"2FECD287",
    x"2FECB4EE",
    x"2FEC9759",
    x"2FEC79C8",
    x"2FEC5C3B",
    x"2FEC3EB1",
    x"2FEC212B",
    x"2FEC03A9",
    x"2FEBE62A",
    x"2FEBC8AF",
    x"2FEBAB38",
    x"2FEB8DC5",
    x"2FEB7055",
    x"2FEB52E9",
    x"2FEB3580",
    x"2FEB181B",
    x"2FEAFABA",
    x"2FEADD5D",
    x"2FEAC003",
    x"2FEAA2AD",
    x"2FEA855A",
    x"2FEA680B",
    x"2FEA4AC0",
    x"2FEA2D78",
    x"2FEA1035",
    x"2FE9F2F4",
    x"2FE9D5B8",
    x"2FE9B87F",
    x"2FE99B4A",
    x"2FE97E18",
    x"2FE960EA",
    x"2FE943C0",
    x"2FE92699",
    x"2FE90976",
    x"2FE8EC57",
    x"2FE8CF3B",
    x"2FE8B223",
    x"2FE8950F",
    x"2FE877FE",
    x"2FE85AF1",
    x"2FE83DE7",
    x"2FE820E1",
    x"2FE803DF",
    x"2FE7E6E0",
    x"2FE7C9E5",
    x"2FE7ACEE",
    x"2FE78FFA",
    x"2FE7730A",
    x"2FE7561D",
    x"2FE73934",
    x"2FE71C4F",
    x"2FE6FF6D",
    x"2FE6E28F",
    x"2FE6C5B5",
    x"2FE6A8DE",
    x"2FE68C0A",
    x"2FE66F3B",
    x"2FE6526E",
    x"2FE635A6",
    x"2FE618E1",
    x"2FE5FC20",
    x"2FE5DF62",
    x"2FE5C2A8",
    x"2FE5A5F1",
    x"2FE5893E",
    x"2FE56C8F",
    x"2FE54FE3",
    x"2FE5333B",
    x"2FE51696",
    x"2FE4F9F5",
    x"2FE4DD58",
    x"2FE4C0BE",
    x"2FE4A428",
    x"2FE48795",
    x"2FE46B06",
    x"2FE44E7A",
    x"2FE431F2",
    x"2FE4156E",
    x"2FE3F8ED",
    x"2FE3DC70",
    x"2FE3BFF6",
    x"2FE3A380",
    x"2FE3870D",
    x"2FE36A9E",
    x"2FE34E32",
    x"2FE331CA",
    x"2FE31566",
    x"2FE2F905",
    x"2FE2DCA8",
    x"2FE2C04E",
    x"2FE2A3F8",
    x"2FE287A5",
    x"2FE26B56",
    x"2FE24F0A",
    x"2FE232C2",
    x"2FE2167D",
    x"2FE1FA3C",
    x"2FE1DDFF",
    x"2FE1C1C5",
    x"2FE1A58E",
    x"2FE1895B",
    x"2FE16D2C",
    x"2FE15100",
    x"2FE134D8",
    x"2FE118B3",
    x"2FE0FC91",
    x"2FE0E074",
    x"2FE0C459",
    x"2FE0A843",
    x"2FE08C2F",
    x"2FE07020",
    x"2FE05413",
    x"2FE0380B",
    x"2FE01C05",
    x"2FE00004",
    x"2FDFE405",
    x"2FDFC80B",
    x"2FDFAC13",
    x"2FDF901F",
    x"2FDF742F",
    x"2FDF5842",
    x"2FDF3C59",
    x"2FDF2073",
    x"2FDF0491",
    x"2FDEE8B2",
    x"2FDECCD7",
    x"2FDEB0FF",
    x"2FDE952B",
    x"2FDE795A",
    x"2FDE5D8C",
    x"2FDE41C2",
    x"2FDE25FC",
    x"2FDE0A39",
    x"2FDDEE79",
    x"2FDDD2BD",
    x"2FDDB705",
    x"2FDD9B4F",
    x"2FDD7F9E",
    x"2FDD63F0",
    x"2FDD4845",
    x"2FDD2C9D",
    x"2FDD10FA",
    x"2FDCF559",
    x"2FDCD9BC",
    x"2FDCBE23",
    x"2FDCA28D",
    x"2FDC86FA",
    x"2FDC6B6B",
    x"2FDC4FDF",
    x"2FDC3457",
    x"2FDC18D2",
    x"2FDBFD51",
    x"2FDBE1D3",
    x"2FDBC658",
    x"2FDBAAE1",
    x"2FDB8F6E",
    x"2FDB73FD",
    x"2FDB5891",
    x"2FDB3D27",
    x"2FDB21C1",
    x"2FDB065F",
    x"2FDAEB00",
    x"2FDACFA4",
    x"2FDAB44C",
    x"2FDA98F7",
    x"2FDA7DA6",
    x"2FDA6258",
    x"2FDA470D",
    x"2FDA2BC6",
    x"2FDA1082",
    x"2FD9F542",
    x"2FD9DA05",
    x"2FD9BECB",
    x"2FD9A395",
    x"2FD98862",
    x"2FD96D33",
    x"2FD95207",
    x"2FD936DE",
    x"2FD91BB9",
    x"2FD90098",
    x"2FD8E579",
    x"2FD8CA5E",
    x"2FD8AF47",
    x"2FD89432",
    x"2FD87922",
    x"2FD85E14",
    x"2FD8430A",
    x"2FD82803",
    x"2FD80D00",
    x"2FD7F200",
    x"2FD7D704",
    x"2FD7BC0A",
    x"2FD7A115",
    x"2FD78622",
    x"2FD76B33",
    x"2FD75047",
    x"2FD7355F",
    x"2FD71A7A",
    x"2FD6FF98",
    x"2FD6E4BA",
    x"2FD6C9DF",
    x"2FD6AF08",
    x"2FD69433",
    x"2FD67962",
    x"2FD65E95",
    x"2FD643CB",
    x"2FD62904",
    x"2FD60E41",
    x"2FD5F380",
    x"2FD5D8C4",
    x"2FD5BE0A",
    x"2FD5A354",
    x"2FD588A1",
    x"2FD56DF2",
    x"2FD55346",
    x"2FD5389D",
    x"2FD51DF8",
    x"2FD50356",
    x"2FD4E8B7",
    x"2FD4CE1C",
    x"2FD4B383",
    x"2FD498EF",
    x"2FD47E5D",
    x"2FD463CF",
    x"2FD44944",
    x"2FD42EBD",
    x"2FD41439",
    x"2FD3F9B8",
    x"2FD3DF3A",
    x"2FD3C4C0",
    x"2FD3AA49",
    x"2FD38FD5",
    x"2FD37565",
    x"2FD35AF8",
    x"2FD3408E",
    x"2FD32628",
    x"2FD30BC5",
    x"2FD2F165",
    x"2FD2D708",
    x"2FD2BCAF",
    x"2FD2A259",
    x"2FD28807",
    x"2FD26DB7",
    x"2FD2536B",
    x"2FD23922",
    x"2FD21EDD",
    x"2FD2049B",
    x"2FD1EA5C",
    x"2FD1D020",
    x"2FD1B5E8",
    x"2FD19BB3",
    x"2FD18181",
    x"2FD16752",
    x"2FD14D27",
    x"2FD132FF",
    x"2FD118DA",
    x"2FD0FEB9",
    x"2FD0E49A",
    x"2FD0CA80",
    x"2FD0B068",
    x"2FD09653",
    x"2FD07C42",
    x"2FD06234",
    x"2FD0482A",
    x"2FD02E22",
    x"2FD0141E",
    x"2FCFFA1D",
    x"2FCFE020",
    x"2FCFC625",
    x"2FCFAC2E",
    x"2FCF923A",
    x"2FCF784A",
    x"2FCF5E5C",
    x"2FCF4472",
    x"2FCF2A8B",
    x"2FCF10A7",
    x"2FCEF6C7",
    x"2FCEDCEA",
    x"2FCEC310",
    x"2FCEA939",
    x"2FCE8F65",
    x"2FCE7595",
    x"2FCE5BC8",
    x"2FCE41FE",
    x"2FCE2837",
    x"2FCE0E74",
    x"2FCDF4B4",
    x"2FCDDAF7",
    x"2FCDC13D",
    x"2FCDA787",
    x"2FCD8DD3",
    x"2FCD7423",
    x"2FCD5A76",
    x"2FCD40CC",
    x"2FCD2726",
    x"2FCD0D83",
    x"2FCCF3E3",
    x"2FCCDA46",
    x"2FCCC0AC",
    x"2FCCA716",
    x"2FCC8D82",
    x"2FCC73F2",
    x"2FCC5A65",
    x"2FCC40DC",
    x"2FCC2755",
    x"2FCC0DD2",
    x"2FCBF452",
    x"2FCBDAD5",
    x"2FCBC15B",
    x"2FCBA7E4",
    x"2FCB8E71",
    x"2FCB7501",
    x"2FCB5B94",
    x"2FCB422A",
    x"2FCB28C3",
    x"2FCB0F60",
    x"2FCAF5FF",
    x"2FCADCA2",
    x"2FCAC348",
    x"2FCAA9F1",
    x"2FCA909E",
    x"2FCA774D",
    x"2FCA5E00",
    x"2FCA44B6",
    x"2FCA2B6F",
    x"2FCA122B",
    x"2FC9F8EA",
    x"2FC9DFAD",
    x"2FC9C672",
    x"2FC9AD3B",
    x"2FC99407",
    x"2FC97AD6",
    x"2FC961A8",
    x"2FC9487E",
    x"2FC92F56",
    x"2FC91632",
    x"2FC8FD10",
    x"2FC8E3F2",
    x"2FC8CAD7",
    x"2FC8B1C0",
    x"2FC898AB",
    x"2FC87F9A",
    x"2FC8668B",
    x"2FC84D80",
    x"2FC83478",
    x"2FC81B73",
    x"2FC80271",
    x"2FC7E972",
    x"2FC7D077",
    x"2FC7B77E",
    x"2FC79E89",
    x"2FC78596",
    x"2FC76CA7",
    x"2FC753BB",
    x"2FC73AD2",
    x"2FC721ED",
    x"2FC7090A",
    x"2FC6F02A",
    x"2FC6D74E",
    x"2FC6BE74",
    x"2FC6A59E",
    x"2FC68CCB",
    x"2FC673FB",
    x"2FC65B2E",
    x"2FC64264",
    x"2FC6299D",
    x"2FC610DA",
    x"2FC5F819",
    x"2FC5DF5C",
    x"2FC5C6A1",
    x"2FC5ADEA",
    x"2FC59536",
    x"2FC57C85",
    x"2FC563D7",
    x"2FC54B2C",
    x"2FC53284",
    x"2FC519DF",
    x"2FC5013E",
    x"2FC4E89F",
    x"2FC4D003",
    x"2FC4B76B",
    x"2FC49ED6",
    x"2FC48643",
    x"2FC46DB4",
    x"2FC45528",
    x"2FC43C9F",
    x"2FC42419",
    x"2FC40B96",
    x"2FC3F316",
    x"2FC3DA99",
    x"2FC3C21F",
    x"2FC3A9A8",
    x"2FC39135",
    x"2FC378C4",
    x"2FC36056",
    x"2FC347EC",
    x"2FC32F84",
    x"2FC31720",
    x"2FC2FEBF",
    x"2FC2E660",
    x"2FC2CE05",
    x"2FC2B5AD",
    x"2FC29D58",
    x"2FC28506",
    x"2FC26CB6",
    x"2FC2546A",
    x"2FC23C21",
    x"2FC223DB",
    x"2FC20B98",
    x"2FC1F358",
    x"2FC1DB1C",
    x"2FC1C2E2",
    x"2FC1AAAB",
    x"2FC19277",
    x"2FC17A46",
    x"2FC16218",
    x"2FC149EE",
    x"2FC131C6",
    x"2FC119A1",
    x"2FC10180",
    x"2FC0E961",
    x"2FC0D145",
    x"2FC0B92D",
    x"2FC0A117",
    x"2FC08904",
    x"2FC070F5",
    x"2FC058E8",
    x"2FC040DE",
    x"2FC028D8",
    x"2FC010D4",
    x"2FBFF8D4",
    x"2FBFE0D6",
    x"2FBFC8DB",
    x"2FBFB0E4",
    x"2FBF98EF",
    x"2FBF80FE",
    x"2FBF690F",
    x"2FBF5123",
    x"2FBF393B",
    x"2FBF2155",
    x"2FBF0972",
    x"2FBEF193",
    x"2FBED9B6",
    x"2FBEC1DC",
    x"2FBEAA05",
    x"2FBE9232",
    x"2FBE7A61",
    x"2FBE6293",
    x"2FBE4AC8",
    x"2FBE3300",
    x"2FBE1B3B",
    x"2FBE037A",
    x"2FBDEBBB",
    x"2FBDD3FF",
    x"2FBDBC46",
    x"2FBDA490",
    x"2FBD8CDC",
    x"2FBD752C",
    x"2FBD5D7F",
    x"2FBD45D5",
    x"2FBD2E2E",
    x"2FBD1689",
    x"2FBCFEE8",
    x"2FBCE74A",
    x"2FBCCFAE",
    x"2FBCB816",
    x"2FBCA080",
    x"2FBC88EE",
    x"2FBC715E",
    x"2FBC59D1",
    x"2FBC4248",
    x"2FBC2AC1",
    x"2FBC133D",
    x"2FBBFBBC",
    x"2FBBE43E",
    x"2FBBCCC3",
    x"2FBBB54B",
    x"2FBB9DD6",
    x"2FBB8663",
    x"2FBB6EF4",
    x"2FBB5788",
    x"2FBB401E",
    x"2FBB28B8",
    x"2FBB1154",
    x"2FBAF9F3",
    x"2FBAE295",
    x"2FBACB3B",
    x"2FBAB3E3",
    x"2FBA9C8E",
    x"2FBA853B",
    x"2FBA6DEC",
    x"2FBA56A0",
    x"2FBA3F57",
    x"2FBA2810",
    x"2FBA10CD",
    x"2FB9F98C",
    x"2FB9E24E",
    x"2FB9CB13",
    x"2FB9B3DB",
    x"2FB99CA6",
    x"2FB98574",
    x"2FB96E45",
    x"2FB95719",
    x"2FB93FEF",
    x"2FB928C9",
    x"2FB911A5",
    x"2FB8FA84",
    x"2FB8E366",
    x"2FB8CC4B",
    x"2FB8B533",
    x"2FB89E1E",
    x"2FB8870C",
    x"2FB86FFC",
    x"2FB858F0",
    x"2FB841E6",
    x"2FB82ADF",
    x"2FB813DB",
    x"2FB7FCDA",
    x"2FB7E5DC",
    x"2FB7CEE1",
    x"2FB7B7E9",
    x"2FB7A0F3",
    x"2FB78A00",
    x"2FB77310",
    x"2FB75C24",
    x"2FB74539",
    x"2FB72E52",
    x"2FB7176E",
    x"2FB7008C",
    x"2FB6E9AE",
    x"2FB6D2D2",
    x"2FB6BBF9",
    x"2FB6A523",
    x"2FB68E50",
    x"2FB6777F",
    x"2FB660B2",
    x"2FB649E7",
    x"2FB6331F",
    x"2FB61C5A",
    x"2FB60598",
    x"2FB5EED9",
    x"2FB5D81D",
    x"2FB5C163",
    x"2FB5AAAC",
    x"2FB593F8",
    x"2FB57D47",
    x"2FB56699",
    x"2FB54FEE",
    x"2FB53945",
    x"2FB5229F",
    x"2FB50BFC",
    x"2FB4F55C",
    x"2FB4DEBF",
    x"2FB4C825",
    x"2FB4B18D",
    x"2FB49AF8",
    x"2FB48466",
    x"2FB46DD7",
    x"2FB4574B",
    x"2FB440C1",
    x"2FB42A3B",
    x"2FB413B7",
    x"2FB3FD36",
    x"2FB3E6B7",
    x"2FB3D03C",
    x"2FB3B9C3",
    x"2FB3A34E",
    x"2FB38CDB",
    x"2FB3766A",
    x"2FB35FFD",
    x"2FB34992",
    x"2FB3332B",
    x"2FB31CC6",
    x"2FB30663",
    x"2FB2F004",
    x"2FB2D9A7",
    x"2FB2C34E",
    x"2FB2ACF6",
    x"2FB296A2",
    x"2FB28051",
    x"2FB26A02",
    x"2FB253B6",
    x"2FB23D6D",
    x"2FB22727",
    x"2FB210E3",
    x"2FB1FAA3",
    x"2FB1E465",
    x"2FB1CE2A",
    x"2FB1B7F1",
    x"2FB1A1BC",
    x"2FB18B89",
    x"2FB17559",
    x"2FB15F2B",
    x"2FB14901",
    x"2FB132D9",
    x"2FB11CB4",
    x"2FB10692",
    x"2FB0F073",
    x"2FB0DA56",
    x"2FB0C43C",
    x"2FB0AE25",
    x"2FB09811",
    x"2FB081FF",
    x"2FB06BF0",
    x"2FB055E4",
    x"2FB03FDB",
    x"2FB029D4",
    x"2FB013D0",
    x"2FAFFDCF",
    x"2FAFE7D1",
    x"2FAFD1D5",
    x"2FAFBBDC",
    x"2FAFA5E6",
    x"2FAF8FF3",
    x"2FAF7A02",
    x"2FAF6414",
    x"2FAF4E29",
    x"2FAF3841",
    x"2FAF225B",
    x"2FAF0C78",
    x"2FAEF698",
    x"2FAEE0BA",
    x"2FAECAE0",
    x"2FAEB508",
    x"2FAE9F32",
    x"2FAE8960",
    x"2FAE7390",
    x"2FAE5DC3",
    x"2FAE47F9",
    x"2FAE3231",
    x"2FAE1C6C",
    x"2FAE06AA",
    x"2FADF0EA",
    x"2FADDB2E",
    x"2FADC574",
    x"2FADAFBC",
    x"2FAD9A08",
    x"2FAD8456",
    x"2FAD6EA7",
    x"2FAD58FA",
    x"2FAD4350",
    x"2FAD2DA9",
    x"2FAD1805",
    x"2FAD0263",
    x"2FACECC4",
    x"2FACD728",
    x"2FACC18F",
    x"2FACABF8",
    x"2FAC9664",
    x"2FAC80D2",
    x"2FAC6B43",
    x"2FAC55B7",
    x"2FAC402E",
    x"2FAC2AA7",
    x"2FAC1523",
    x"2FABFFA2",
    x"2FABEA23",
    x"2FABD4A7",
    x"2FABBF2E",
    x"2FABA9B8",
    x"2FAB9444",
    x"2FAB7ED3",
    x"2FAB6964",
    x"2FAB53F8",
    x"2FAB3E8F",
    x"2FAB2929",
    x"2FAB13C5",
    x"2FAAFE64",
    x"2FAAE905",
    x"2FAAD3A9",
    x"2FAABE50",
    x"2FAAA8FA",
    x"2FAA93A6",
    x"2FAA7E55",
    x"2FAA6906",
    x"2FAA53BB",
    x"2FAA3E72",
    x"2FAA292B",
    x"2FAA13E7",
    x"2FA9FEA6",
    x"2FA9E968",
    x"2FA9D42C",
    x"2FA9BEF3",
    x"2FA9A9BC",
    x"2FA99488",
    x"2FA97F57",
    x"2FA96A28",
    x"2FA954FC",
    x"2FA93FD3",
    x"2FA92AAC",
    x"2FA91588",
    x"2FA90067",
    x"2FA8EB48",
    x"2FA8D62C",
    x"2FA8C113",
    x"2FA8ABFC",
    x"2FA896E8",
    x"2FA881D6",
    x"2FA86CC7",
    x"2FA857BB",
    x"2FA842B1",
    x"2FA82DAA",
    x"2FA818A6",
    x"2FA803A4",
    x"2FA7EEA5",
    x"2FA7D9A8",
    x"2FA7C4AF",
    x"2FA7AFB7",
    x"2FA79AC3",
    x"2FA785D1",
    x"2FA770E1",
    x"2FA75BF4",
    x"2FA7470A",
    x"2FA73223",
    x"2FA71D3E",
    x"2FA7085B",
    x"2FA6F37C",
    x"2FA6DE9E",
    x"2FA6C9C4",
    x"2FA6B4EC",
    x"2FA6A017",
    x"2FA68B44",
    x"2FA67674",
    x"2FA661A6",
    x"2FA64CDB",
    x"2FA63813",
    x"2FA6234D",
    x"2FA60E8A",
    x"2FA5F9CA",
    x"2FA5E50C",
    x"2FA5D051",
    x"2FA5BB98",
    x"2FA5A6E2",
    x"2FA5922E",
    x"2FA57D7D",
    x"2FA568CF",
    x"2FA55423",
    x"2FA53F7A",
    x"2FA52AD3",
    x"2FA5162F",
    x"2FA5018D",
    x"2FA4ECEF",
    x"2FA4D852",
    x"2FA4C3B8",
    x"2FA4AF21",
    x"2FA49A8D",
    x"2FA485FB",
    x"2FA4716B",
    x"2FA45CDE",
    x"2FA44854",
    x"2FA433CC",
    x"2FA41F47",
    x"2FA40AC4",
    x"2FA3F644",
    x"2FA3E1C7",
    x"2FA3CD4C",
    x"2FA3B8D4",
    x"2FA3A45E",
    x"2FA38FEA",
    x"2FA37B7A",
    x"2FA3670C",
    x"2FA352A0",
    x"2FA33E37",
    x"2FA329D0",
    x"2FA3156C",
    x"2FA3010B",
    x"2FA2ECAC",
    x"2FA2D850",
    x"2FA2C3F6",
    x"2FA2AF9F",
    x"2FA29B4A",
    x"2FA286F8",
    x"2FA272A8",
    x"2FA25E5B",
    x"2FA24A11",
    x"2FA235C9",
    x"2FA22183",
    x"2FA20D40",
    x"2FA1F900",
    x"2FA1E4C2",
    x"2FA1D087",
    x"2FA1BC4E",
    x"2FA1A818",
    x"2FA193E4",
    x"2FA17FB3",
    x"2FA16B84",
    x"2FA15758",
    x"2FA1432E",
    x"2FA12F07",
    x"2FA11AE3",
    x"2FA106C0",
    x"2FA0F2A1",
    x"2FA0DE84",
    x"2FA0CA69",
    x"2FA0B651",
    x"2FA0A23C",
    x"2FA08E29",
    x"2FA07A18",
    x"2FA0660A",
    x"2FA051FF",
    x"2FA03DF6",
    x"2FA029EF",
    x"2FA015EB",
    x"2FA001EA",
    x"2F9FEDEB",
    x"2F9FD9EE",
    x"2F9FC5F4",
    x"2F9FB1FD",
    x"2F9F9E08",
    x"2F9F8A15",
    x"2F9F7625",
    x"2F9F6238",
    x"2F9F4E4D",
    x"2F9F3A64",
    x"2F9F267E",
    x"2F9F129A",
    x"2F9EFEB9",
    x"2F9EEADB",
    x"2F9ED6FF",
    x"2F9EC325",
    x"2F9EAF4E",
    x"2F9E9B79",
    x"2F9E87A7",
    x"2F9E73D7",
    x"2F9E600A",
    x"2F9E4C3F",
    x"2F9E3877",
    x"2F9E24B1",
    x"2F9E10EE",
    x"2F9DFD2D",
    x"2F9DE96E",
    x"2F9DD5B3",
    x"2F9DC1F9",
    x"2F9DAE42",
    x"2F9D9A8E",
    x"2F9D86DB",
    x"2F9D732C",
    x"2F9D5F7F",
    x"2F9D4BD4",
    x"2F9D382C",
    x"2F9D2486",
    x"2F9D10E3",
    x"2F9CFD42",
    x"2F9CE9A3",
    x"2F9CD607",
    x"2F9CC26E",
    x"2F9CAED7",
    x"2F9C9B42",
    x"2F9C87B0",
    x"2F9C7420",
    x"2F9C6093",
    x"2F9C4D08",
    x"2F9C3980",
    x"2F9C25FA",
    x"2F9C1276",
    x"2F9BFEF5",
    x"2F9BEB76",
    x"2F9BD7FA",
    x"2F9BC480",
    x"2F9BB109",
    x"2F9B9D94",
    x"2F9B8A22",
    x"2F9B76B2",
    x"2F9B6344",
    x"2F9B4FD9",
    x"2F9B3C70",
    x"2F9B290A",
    x"2F9B15A6",
    x"2F9B0244",
    x"2F9AEEE5",
    x"2F9ADB88",
    x"2F9AC82E",
    x"2F9AB4D6",
    x"2F9AA181",
    x"2F9A8E2E",
    x"2F9A7ADD",
    x"2F9A678F",
    x"2F9A5444",
    x"2F9A40FA",
    x"2F9A2DB3",
    x"2F9A1A6F",
    x"2F9A072D",
    x"2F99F3ED",
    x"2F99E0B0",
    x"2F99CD75",
    x"2F99BA3C",
    x"2F99A706",
    x"2F9993D3",
    x"2F9980A1",
    x"2F996D72",
    x"2F995A46",
    x"2F99471C",
    x"2F9933F4",
    x"2F9920CF",
    x"2F990DAC",
    x"2F98FA8B",
    x"2F98E76D",
    x"2F98D452",
    x"2F98C138",
    x"2F98AE21",
    x"2F989B0D",
    x"2F9887FB",
    x"2F9874EB",
    x"2F9861DD",
    x"2F984ED2",
    x"2F983BCA",
    x"2F9828C3",
    x"2F9815BF",
    x"2F9802BE",
    x"2F97EFBF",
    x"2F97DCC2",
    x"2F97C9C8",
    x"2F97B6D0",
    x"2F97A3DA",
    x"2F9790E7",
    x"2F977DF6",
    x"2F976B07",
    x"2F97581B",
    x"2F974531",
    x"2F97324A",
    x"2F971F64",
    x"2F970C82",
    x"2F96F9A1",
    x"2F96E6C3",
    x"2F96D3E8",
    x"2F96C10E",
    x"2F96AE37",
    x"2F969B63",
    x"2F968891",
    x"2F9675C1",
    x"2F9662F3",
    x"2F965028",
    x"2F963D5F",
    x"2F962A99",
    x"2F9617D4",
    x"2F960513",
    x"2F95F253",
    x"2F95DF96",
    x"2F95CCDB",
    x"2F95BA23",
    x"2F95A76D",
    x"2F9594B9",
    x"2F958208",
    x"2F956F58",
    x"2F955CAC",
    x"2F954A01",
    x"2F953759",
    x"2F9524B3",
    x"2F951210",
    x"2F94FF6F",
    x"2F94ECD0",
    x"2F94DA34",
    x"2F94C79A",
    x"2F94B502",
    x"2F94A26C",
    x"2F948FD9",
    x"2F947D48",
    x"2F946ABA",
    x"2F94582E",
    x"2F9445A4",
    x"2F94331C",
    x"2F942097",
    x"2F940E14",
    x"2F93FB94",
    x"2F93E915",
    x"2F93D699",
    x"2F93C420",
    x"2F93B1A8",
    x"2F939F33",
    x"2F938CC0",
    x"2F937A50",
    x"2F9367E2",
    x"2F935576",
    x"2F93430C",
    x"2F9330A5",
    x"2F931E40",
    x"2F930BDE",
    x"2F92F97D",
    x"2F92E71F",
    x"2F92D4C4",
    x"2F92C26A",
    x"2F92B013",
    x"2F929DBE",
    x"2F928B6C",
    x"2F92791B",
    x"2F9266CD",
    x"2F925482",
    x"2F924238",
    x"2F922FF1",
    x"2F921DAC",
    x"2F920B6A",
    x"2F91F929",
    x"2F91E6EB",
    x"2F91D4B0",
    x"2F91C276",
    x"2F91B03F",
    x"2F919E0A",
    x"2F918BD7",
    x"2F9179A7",
    x"2F916779",
    x"2F91554D",
    x"2F914324",
    x"2F9130FC",
    x"2F911ED7",
    x"2F910CB5",
    x"2F90FA94",
    x"2F90E876",
    x"2F90D65A",
    x"2F90C441",
    x"2F90B229",
    x"2F90A014",
    x"2F908E01",
    x"2F907BF0",
    x"2F9069E2",
    x"2F9057D6",
    x"2F9045CC",
    x"2F9033C5",
    x"2F9021BF",
    x"2F900FBC",
    x"2F8FFDBB",
    x"2F8FEBBD",
    x"2F8FD9C0",
    x"2F8FC7C6",
    x"2F8FB5CE",
    x"2F8FA3D9",
    x"2F8F91E5",
    x"2F8F7FF4",
    x"2F8F6E05",
    x"2F8F5C19",
    x"2F8F4A2E",
    x"2F8F3846",
    x"2F8F2660",
    x"2F8F147D",
    x"2F8F029B",
    x"2F8EF0BC",
    x"2F8EDEDF",
    x"2F8ECD04",
    x"2F8EBB2C",
    x"2F8EA955",
    x"2F8E9781",
    x"2F8E85B0",
    x"2F8E73E0",
    x"2F8E6213",
    x"2F8E5048",
    x"2F8E3E7F",
    x"2F8E2CB8",
    x"2F8E1AF3",
    x"2F8E0931",
    x"2F8DF771",
    x"2F8DE5B3",
    x"2F8DD3F8",
    x"2F8DC23E",
    x"2F8DB087",
    x"2F8D9ED2",
    x"2F8D8D1F",
    x"2F8D7B6F",
    x"2F8D69C1",
    x"2F8D5814",
    x"2F8D466B",
    x"2F8D34C3",
    x"2F8D231D",
    x"2F8D117A",
    x"2F8CFFD9",
    x"2F8CEE3A",
    x"2F8CDC9D",
    x"2F8CCB03",
    x"2F8CB96B",
    x"2F8CA7D5",
    x"2F8C9641",
    x"2F8C84AF",
    x"2F8C7320",
    x"2F8C6192",
    x"2F8C5007",
    x"2F8C3E7E",
    x"2F8C2CF8",
    x"2F8C1B73",
    x"2F8C09F1",
    x"2F8BF871",
    x"2F8BE6F3",
    x"2F8BD577",
    x"2F8BC3FD",
    x"2F8BB286",
    x"2F8BA111",
    x"2F8B8F9E",
    x"2F8B7E2D",
    x"2F8B6CBE",
    x"2F8B5B51",
    x"2F8B49E7",
    x"2F8B387F",
    x"2F8B2719",
    x"2F8B15B5",
    x"2F8B0454",
    x"2F8AF2F4",
    x"2F8AE197",
    x"2F8AD03C",
    x"2F8ABEE3",
    x"2F8AAD8C",
    x"2F8A9C37",
    x"2F8A8AE5",
    x"2F8A7995",
    x"2F8A6847",
    x"2F8A56FB",
    x"2F8A45B1",
    x"2F8A3469",
    x"2F8A2324",
    x"2F8A11E0",
    x"2F8A009F",
    x"2F89EF60",
    x"2F89DE23",
    x"2F89CCE9",
    x"2F89BBB0",
    x"2F89AA7A",
    x"2F899946",
    x"2F898813",
    x"2F8976E4",
    x"2F8965B6",
    x"2F89548A",
    x"2F894361",
    x"2F893239",
    x"2F892114",
    x"2F890FF1",
    x"2F88FED0",
    x"2F88EDB1",
    x"2F88DC95",
    x"2F88CB7A",
    x"2F88BA62",
    x"2F88A94C",
    x"2F889837",
    x"2F888725",
    x"2F887616",
    x"2F886508",
    x"2F8853FC",
    x"2F8842F3",
    x"2F8831EC",
    x"2F8820E6",
    x"2F880FE3",
    x"2F87FEE3",
    x"2F87EDE4",
    x"2F87DCE7",
    x"2F87CBEC",
    x"2F87BAF4",
    x"2F87A9FE",
    x"2F87990A",
    x"2F878817",
    x"2F877728",
    x"2F87663A",
    x"2F87554E",
    x"2F874464",
    x"2F87337D",
    x"2F872298",
    x"2F8711B4",
    x"2F8700D3",
    x"2F86EFF4",
    x"2F86DF17",
    x"2F86CE3C",
    x"2F86BD64",
    x"2F86AC8D",
    x"2F869BB8",
    x"2F868AE6",
    x"2F867A16",
    x"2F866947",
    x"2F86587B",
    x"2F8647B1",
    x"2F8636E9",
    x"2F862624",
    x"2F861560",
    x"2F86049E",
    x"2F85F3DF",
    x"2F85E321",
    x"2F85D266",
    x"2F85C1AD",
    x"2F85B0F6",
    x"2F85A040",
    x"2F858F8D",
    x"2F857EDD",
    x"2F856E2E",
    x"2F855D81",
    x"2F854CD6",
    x"2F853C2E",
    x"2F852B87",
    x"2F851AE3",
    x"2F850A41",
    x"2F84F9A0",
    x"2F84E902",
    x"2F84D866",
    x"2F84C7CC",
    x"2F84B734",
    x"2F84A69E",
    x"2F84960B",
    x"2F848579",
    x"2F8474E9",
    x"2F84645C",
    x"2F8453D0",
    x"2F844347",
    x"2F8432BF",
    x"2F84223A",
    x"2F8411B7",
    x"2F840135",
    x"2F83F0B6",
    x"2F83E039",
    x"2F83CFBE",
    x"2F83BF45",
    x"2F83AECE",
    x"2F839E5A",
    x"2F838DE7",
    x"2F837D76",
    x"2F836D08",
    x"2F835C9B",
    x"2F834C30",
    x"2F833BC8",
    x"2F832B61",
    x"2F831AFD",
    x"2F830A9B",
    x"2F82FA3A",
    x"2F82E9DC",
    x"2F82D980",
    x"2F82C926",
    x"2F82B8CE",
    x"2F82A878",
    x"2F829824",
    x"2F8287D2",
    x"2F827782",
    x"2F826734",
    x"2F8256E8",
    x"2F82469E",
    x"2F823656",
    x"2F822610",
    x"2F8215CD",
    x"2F82058B",
    x"2F81F54B",
    x"2F81E50E",
    x"2F81D4D2",
    x"2F81C498",
    x"2F81B461",
    x"2F81A42B",
    x"2F8193F8",
    x"2F8183C6",
    x"2F817397",
    x"2F816369",
    x"2F81533E",
    x"2F814315",
    x"2F8132ED",
    x"2F8122C8",
    x"2F8112A4",
    x"2F810283",
    x"2F80F264",
    x"2F80E247",
    x"2F80D22B",
    x"2F80C212",
    x"2F80B1FB",
    x"2F80A1E6",
    x"2F8091D2",
    x"2F8081C1",
    x"2F8071B2",
    x"2F8061A5",
    x"2F805199",
    x"2F804190",
    x"2F803189",
    x"2F802184",
    x"2F801181",
    x"2F80017F",
    x"2F7FE301",
    x"2F7FC306",
    x"2F7FA310",
    x"2F7F831D",
    x"2F7F632F",
    x"2F7F4345",
    x"2F7F235E",
    x"2F7F037C",
    x"2F7EE39D",
    x"2F7EC3C3",
    x"2F7EA3EC",
    x"2F7E841A",
    x"2F7E644B",
    x"2F7E4481",
    x"2F7E24BA",
    x"2F7E04F8",
    x"2F7DE539",
    x"2F7DC57E",
    x"2F7DA5C8",
    x"2F7D8615",
    x"2F7D6666",
    x"2F7D46BB",
    x"2F7D2714",
    x"2F7D0772",
    x"2F7CE7D3",
    x"2F7CC838",
    x"2F7CA8A1",
    x"2F7C890D",
    x"2F7C697E",
    x"2F7C49F3",
    x"2F7C2A6C",
    x"2F7C0AE8",
    x"2F7BEB69",
    x"2F7BCBEE",
    x"2F7BAC76",
    x"2F7B8D03",
    x"2F7B6D93",
    x"2F7B4E27",
    x"2F7B2EBF",
    x"2F7B0F5B",
    x"2F7AEFFB",
    x"2F7AD09F",
    x"2F7AB147",
    x"2F7A91F3",
    x"2F7A72A3",
    x"2F7A5356",
    x"2F7A340E",
    x"2F7A14C9",
    x"2F79F589",
    x"2F79D64C",
    x"2F79B713",
    x"2F7997DE",
    x"2F7978AD",
    x"2F795980",
    x"2F793A57",
    x"2F791B32",
    x"2F78FC10",
    x"2F78DCF3",
    x"2F78BDD9",
    x"2F789EC3",
    x"2F787FB1",
    x"2F7860A3",
    x"2F784199",
    x"2F782293",
    x"2F780390",
    x"2F77E492",
    x"2F77C597",
    x"2F77A6A0",
    x"2F7787AE",
    x"2F7768BF",
    x"2F7749D3",
    x"2F772AEC",
    x"2F770C09",
    x"2F76ED29",
    x"2F76CE4D",
    x"2F76AF75",
    x"2F7690A1",
    x"2F7671D1",
    x"2F765305",
    x"2F76343D",
    x"2F761578",
    x"2F75F6B7",
    x"2F75D7FA",
    x"2F75B941",
    x"2F759A8C",
    x"2F757BDB",
    x"2F755D2D",
    x"2F753E83",
    x"2F751FDD",
    x"2F75013B",
    x"2F74E29D",
    x"2F74C403",
    x"2F74A56C",
    x"2F7486D9",
    x"2F74684A",
    x"2F7449BF",
    x"2F742B38",
    x"2F740CB4",
    x"2F73EE35",
    x"2F73CFB9",
    x"2F73B141",
    x"2F7392CD",
    x"2F73745C",
    x"2F7355EF",
    x"2F733787",
    x"2F731922",
    x"2F72FAC0",
    x"2F72DC63",
    x"2F72BE09",
    x"2F729FB3",
    x"2F728161",
    x"2F726313",
    x"2F7244C9",
    x"2F722682",
    x"2F72083F",
    x"2F71EA00",
    x"2F71CBC4",
    x"2F71AD8D",
    x"2F718F59",
    x"2F717129",
    x"2F7152FD",
    x"2F7134D4",
    x"2F7116B0",
    x"2F70F88F",
    x"2F70DA71",
    x"2F70BC58",
    x"2F709E42",
    x"2F708030",
    x"2F706222",
    x"2F704418",
    x"2F702611",
    x"2F70080E",
    x"2F6FEA0F",
    x"2F6FCC14",
    x"2F6FAE1C",
    x"2F6F9028",
    x"2F6F7238",
    x"2F6F544C",
    x"2F6F3663",
    x"2F6F187E",
    x"2F6EFA9D",
    x"2F6EDCBF",
    x"2F6EBEE6",
    x"2F6EA110",
    x"2F6E833D",
    x"2F6E656F",
    x"2F6E47A4",
    x"2F6E29DD",
    x"2F6E0C1A",
    x"2F6DEE5A",
    x"2F6DD09E",
    x"2F6DB2E6",
    x"2F6D9531",
    x"2F6D7781",
    x"2F6D59D3",
    x"2F6D3C2A",
    x"2F6D1E84",
    x"2F6D00E2",
    x"2F6CE344",
    x"2F6CC5AA",
    x"2F6CA813",
    x"2F6C8A80",
    x"2F6C6CF0",
    x"2F6C4F64",
    x"2F6C31DC",
    x"2F6C1458",
    x"2F6BF6D7",
    x"2F6BD95A",
    x"2F6BBBE1",
    x"2F6B9E6B",
    x"2F6B80F9",
    x"2F6B638B",
    x"2F6B4620",
    x"2F6B28B9",
    x"2F6B0B56",
    x"2F6AEDF7",
    x"2F6AD09B",
    x"2F6AB342",
    x"2F6A95EE",
    x"2F6A789D",
    x"2F6A5B50",
    x"2F6A3E06",
    x"2F6A20C0",
    x"2F6A037E",
    x"2F69E63F",
    x"2F69C904",
    x"2F69ABCD",
    x"2F698E99",
    x"2F697169",
    x"2F69543D",
    x"2F693714",
    x"2F6919EF",
    x"2F68FCCE",
    x"2F68DFB0",
    x"2F68C296",
    x"2F68A580",
    x"2F68886D",
    x"2F686B5D",
    x"2F684E52",
    x"2F68314A",
    x"2F681445",
    x"2F67F745",
    x"2F67DA48",
    x"2F67BD4E",
    x"2F67A058",
    x"2F678366",
    x"2F676677",
    x"2F67498C",
    x"2F672CA5",
    x"2F670FC1",
    x"2F66F2E1",
    x"2F66D605",
    x"2F66B92C",
    x"2F669C56",
    x"2F667F85",
    x"2F6662B6",
    x"2F6645EC",
    x"2F662925",
    x"2F660C62",
    x"2F65EFA2",
    x"2F65D2E6",
    x"2F65B62D",
    x"2F659978",
    x"2F657CC7",
    x"2F656019",
    x"2F65436F",
    x"2F6526C8",
    x"2F650A25",
    x"2F64ED86",
    x"2F64D0EA",
    x"2F64B451",
    x"2F6497BD",
    x"2F647B2B",
    x"2F645E9E",
    x"2F644214",
    x"2F64258D",
    x"2F64090A",
    x"2F63EC8B",
    x"2F63D00F",
    x"2F63B397",
    x"2F639722",
    x"2F637AB1",
    x"2F635E44",
    x"2F6341DA",
    x"2F632573",
    x"2F630910",
    x"2F62ECB1",
    x"2F62D055",
    x"2F62B3FD",
    x"2F6297A8",
    x"2F627B57",
    x"2F625F09",
    x"2F6242BF",
    x"2F622679",
    x"2F620A36",
    x"2F61EDF6",
    x"2F61D1BA",
    x"2F61B582",
    x"2F61994D",
    x"2F617D1B",
    x"2F6160ED",
    x"2F6144C3",
    x"2F61289C",
    x"2F610C79",
    x"2F60F059",
    x"2F60D43D",
    x"2F60B824",
    x"2F609C0F",
    x"2F607FFD",
    x"2F6063EF",
    x"2F6047E4",
    x"2F602BDD",
    x"2F600FD9",
    x"2F5FF3D9",
    x"2F5FD7DC",
    x"2F5FBBE3",
    x"2F5F9FED",
    x"2F5F83FB",
    x"2F5F680C",
    x"2F5F4C21",
    x"2F5F3039",
    x"2F5F1455",
    x"2F5EF874",
    x"2F5EDC97",
    x"2F5EC0BD",
    x"2F5EA4E7",
    x"2F5E8914",
    x"2F5E6D44",
    x"2F5E5178",
    x"2F5E35B0",
    x"2F5E19EB",
    x"2F5DFE29",
    x"2F5DE26B",
    x"2F5DC6B1",
    x"2F5DAAFA",
    x"2F5D8F46",
    x"2F5D7396",
    x"2F5D57E9",
    x"2F5D3C40",
    x"2F5D209A",
    x"2F5D04F8",
    x"2F5CE959",
    x"2F5CCDBD",
    x"2F5CB225",
    x"2F5C9691",
    x"2F5C7B00",
    x"2F5C5F72",
    x"2F5C43E8",
    x"2F5C2861",
    x"2F5C0CDE",
    x"2F5BF15E",
    x"2F5BD5E1",
    x"2F5BBA68",
    x"2F5B9EF3",
    x"2F5B8381",
    x"2F5B6812",
    x"2F5B4CA7",
    x"2F5B313F",
    x"2F5B15DA",
    x"2F5AFA79",
    x"2F5ADF1C",
    x"2F5AC3C2",
    x"2F5AA86B",
    x"2F5A8D17",
    x"2F5A71C8",
    x"2F5A567B",
    x"2F5A3B32",
    x"2F5A1FEC",
    x"2F5A04AA",
    x"2F59E96B",
    x"2F59CE30",
    x"2F59B2F8",
    x"2F5997C3",
    x"2F597C92",
    x"2F596164",
    x"2F594639",
    x"2F592B12",
    x"2F590FEE",
    x"2F58F4CE",
    x"2F58D9B1",
    x"2F58BE98",
    x"2F58A382",
    x"2F58886F",
    x"2F586D5F",
    x"2F585254",
    x"2F58374B",
    x"2F581C46",
    x"2F580144",
    x"2F57E645",
    x"2F57CB4A",
    x"2F57B053",
    x"2F57955E",
    x"2F577A6D",
    x"2F575F80",
    x"2F574495",
    x"2F5729AE",
    x"2F570ECB",
    x"2F56F3EB",
    x"2F56D90E",
    x"2F56BE34",
    x"2F56A35E",
    x"2F56888C",
    x"2F566DBC",
    x"2F5652F0",
    x"2F563828",
    x"2F561D62",
    x"2F5602A0",
    x"2F55E7E2",
    x"2F55CD26",
    x"2F55B26E",
    x"2F5597BA",
    x"2F557D08",
    x"2F55625A",
    x"2F5547B0",
    x"2F552D08",
    x"2F551264",
    x"2F54F7C4",
    x"2F54DD27",
    x"2F54C28D",
    x"2F54A7F6",
    x"2F548D63",
    x"2F5472D3",
    x"2F545846",
    x"2F543DBC",
    x"2F542336",
    x"2F5408B4",
    x"2F53EE34",
    x"2F53D3B8",
    x"2F53B93F",
    x"2F539ECA",
    x"2F538458",
    x"2F5369E9",
    x"2F534F7D",
    x"2F533515",
    x"2F531AB0",
    x"2F53004E",
    x"2F52E5F0",
    x"2F52CB95",
    x"2F52B13D",
    x"2F5296E8",
    x"2F527C97",
    x"2F526249",
    x"2F5247FF",
    x"2F522DB7",
    x"2F521373",
    x"2F51F932",
    x"2F51DEF5",
    x"2F51C4BB",
    x"2F51AA84",
    x"2F519050",
    x"2F517620",
    x"2F515BF2",
    x"2F5141C9",
    x"2F5127A2",
    x"2F510D7F",
    x"2F50F35F",
    x"2F50D942",
    x"2F50BF28",
    x"2F50A512",
    x"2F508AFF",
    x"2F5070EF",
    x"2F5056E3",
    x"2F503CDA",
    x"2F5022D4",
    x"2F5008D1",
    x"2F4FEED1",
    x"2F4FD4D5",
    x"2F4FBADC",
    x"2F4FA0E6",
    x"2F4F86F4",
    x"2F4F6D05",
    x"2F4F5319",
    x"2F4F3930",
    x"2F4F1F4A",
    x"2F4F0568",
    x"2F4EEB89",
    x"2F4ED1AD",
    x"2F4EB7D5",
    x"2F4E9DFF",
    x"2F4E842D",
    x"2F4E6A5E",
    x"2F4E5093",
    x"2F4E36CA",
    x"2F4E1D05",
    x"2F4E0343",
    x"2F4DE984",
    x"2F4DCFC8",
    x"2F4DB610",
    x"2F4D9C5B",
    x"2F4D82A9",
    x"2F4D68FA",
    x"2F4D4F4F",
    x"2F4D35A6",
    x"2F4D1C01",
    x"2F4D025F",
    x"2F4CE8C1",
    x"2F4CCF25",
    x"2F4CB58D",
    x"2F4C9BF8",
    x"2F4C8266",
    x"2F4C68D7",
    x"2F4C4F4C",
    x"2F4C35C3",
    x"2F4C1C3E",
    x"2F4C02BC",
    x"2F4BE93E",
    x"2F4BCFC2",
    x"2F4BB64A",
    x"2F4B9CD4",
    x"2F4B8362",
    x"2F4B69F4",
    x"2F4B5088",
    x"2F4B3720",
    x"2F4B1DBA",
    x"2F4B0458",
    x"2F4AEAF9",
    x"2F4AD19D",
    x"2F4AB845",
    x"2F4A9EEF",
    x"2F4A859D",
    x"2F4A6C4E",
    x"2F4A5302",
    x"2F4A39B9",
    x"2F4A2073",
    x"2F4A0731",
    x"2F49EDF2",
    x"2F49D4B6",
    x"2F49BB7C",
    x"2F49A247",
    x"2F498914",
    x"2F496FE4",
    x"2F4956B8",
    x"2F493D8F",
    x"2F492469",
    x"2F490B46",
    x"2F48F226",
    x"2F48D909",
    x"2F48BFEF",
    x"2F48A6D9",
    x"2F488DC6",
    x"2F4874B6",
    x"2F485BA9",
    x"2F48429F",
    x"2F482998",
    x"2F481094",
    x"2F47F794",
    x"2F47DE96",
    x"2F47C59C",
    x"2F47ACA5",
    x"2F4793B1",
    x"2F477AC0",
    x"2F4761D2",
    x"2F4748E8",
    x"2F473000",
    x"2F47171C",
    x"2F46FE3A",
    x"2F46E55C",
    x"2F46CC81",
    x"2F46B3A9",
    x"2F469AD4",
    x"2F468202",
    x"2F466934",
    x"2F465068",
    x"2F46379F",
    x"2F461EDA",
    x"2F460618",
    x"2F45ED59",
    x"2F45D49C",
    x"2F45BBE3",
    x"2F45A32D",
    x"2F458A7B",
    x"2F4571CB",
    x"2F45591E",
    x"2F454075",
    x"2F4527CE",
    x"2F450F2B",
    x"2F44F68A",
    x"2F44DDED",
    x"2F44C553",
    x"2F44ACBC",
    x"2F449428",
    x"2F447B97",
    x"2F446309",
    x"2F444A7E",
    x"2F4431F6",
    x"2F441971",
    x"2F4400F0",
    x"2F43E871",
    x"2F43CFF6",
    x"2F43B77D",
    x"2F439F08",
    x"2F438695",
    x"2F436E26",
    x"2F4355BA",
    x"2F433D51",
    x"2F4324EA",
    x"2F430C87",
    x"2F42F427",
    x"2F42DBCA",
    x"2F42C370",
    x"2F42AB19",
    x"2F4292C6",
    x"2F427A75",
    x"2F426227",
    x"2F4249DC",
    x"2F423195",
    x"2F421950",
    x"2F42010E",
    x"2F41E8D0",
    x"2F41D094",
    x"2F41B85B",
    x"2F41A026",
    x"2F4187F3",
    x"2F416FC4",
    x"2F415797",
    x"2F413F6E",
    x"2F412748",
    x"2F410F24",
    x"2F40F704",
    x"2F40DEE6",
    x"2F40C6CC",
    x"2F40AEB5",
    x"2F4096A0",
    x"2F407E8F",
    x"2F406681",
    x"2F404E75",
    x"2F40366D",
    x"2F401E68",
    x"2F400666",
    x"2F3FEE66",
    x"2F3FD66A",
    x"2F3FBE71",
    x"2F3FA67A",
    x"2F3F8E87",
    x"2F3F7697",
    x"2F3F5EA9",
    x"2F3F46BF",
    x"2F3F2ED8",
    x"2F3F16F3",
    x"2F3EFF12",
    x"2F3EE734",
    x"2F3ECF58",
    x"2F3EB780",
    x"2F3E9FAA",
    x"2F3E87D8",
    x"2F3E7008",
    x"2F3E583C",
    x"2F3E4072",
    x"2F3E28AC",
    x"2F3E10E8",
    x"2F3DF927",
    x"2F3DE16A",
    x"2F3DC9AF",
    x"2F3DB1F7",
    x"2F3D9A43",
    x"2F3D8291",
    x"2F3D6AE2",
    x"2F3D5336",
    x"2F3D3B8D",
    x"2F3D23E7",
    x"2F3D0C44",
    x"2F3CF4A4",
    x"2F3CDD07",
    x"2F3CC56D",
    x"2F3CADD6",
    x"2F3C9641",
    x"2F3C7EB0",
    x"2F3C6722",
    x"2F3C4F96",
    x"2F3C380E",
    x"2F3C2088",
    x"2F3C0906",
    x"2F3BF186",
    x"2F3BDA09",
    x"2F3BC290",
    x"2F3BAB19",
    x"2F3B93A5",
    x"2F3B7C34",
    x"2F3B64C6",
    x"2F3B4D5B",
    x"2F3B35F2",
    x"2F3B1E8D",
    x"2F3B072B",
    x"2F3AEFCB",
    x"2F3AD86F",
    x"2F3AC115",
    x"2F3AA9BF",
    x"2F3A926B",
    x"2F3A7B1A",
    x"2F3A63CC",
    x"2F3A4C81",
    x"2F3A3539",
    x"2F3A1DF4",
    x"2F3A06B1",
    x"2F39EF72",
    x"2F39D836",
    x"2F39C0FC",
    x"2F39A9C5",
    x"2F399291",
    x"2F397B61",
    x"2F396433",
    x"2F394D08",
    x"2F3935DF",
    x"2F391EBA",
    x"2F390798",
    x"2F38F078",
    x"2F38D95C",
    x"2F38C242",
    x"2F38AB2B",
    x"2F389417",
    x"2F387D06",
    x"2F3865F8",
    x"2F384EED",
    x"2F3837E4",
    x"2F3820DF",
    x"2F3809DC",
    x"2F37F2DC",
    x"2F37DBDF",
    x"2F37C4E5",
    x"2F37ADEE",
    x"2F3796FA",
    x"2F378008",
    x"2F37691A",
    x"2F37522E",
    x"2F373B45",
    x"2F37245F",
    x"2F370D7C",
    x"2F36F69C",
    x"2F36DFBE",
    x"2F36C8E4",
    x"2F36B20C",
    x"2F369B37",
    x"2F368465",
    x"2F366D96",
    x"2F3656CA",
    x"2F364000",
    x"2F36293A",
    x"2F361276",
    x"2F35FBB5",
    x"2F35E4F7",
    x"2F35CE3C",
    x"2F35B784",
    x"2F35A0CE",
    x"2F358A1B",
    x"2F35736C",
    x"2F355CBF",
    x"2F354614",
    x"2F352F6D",
    x"2F3518C9",
    x"2F350227",
    x"2F34EB88",
    x"2F34D4EC",
    x"2F34BE53",
    x"2F34A7BC",
    x"2F349129",
    x"2F347A98",
    x"2F34640A",
    x"2F344D7F",
    x"2F3436F7",
    x"2F342071",
    x"2F3409EF",
    x"2F33F36F",
    x"2F33DCF2",
    x"2F33C678",
    x"2F33B000",
    x"2F33998C",
    x"2F33831A",
    x"2F336CAB",
    x"2F33563F",
    x"2F333FD5",
    x"2F33296F",
    x"2F33130B",
    x"2F32FCAA",
    x"2F32E64C",
    x"2F32CFF0",
    x"2F32B998",
    x"2F32A342",
    x"2F328CEF",
    x"2F32769F",
    x"2F326051",
    x"2F324A07",
    x"2F3233BF",
    x"2F321D7A",
    x"2F320737",
    x"2F31F0F8",
    x"2F31DABB",
    x"2F31C481",
    x"2F31AE4A",
    x"2F319816",
    x"2F3181E4",
    x"2F316BB5",
    x"2F315589",
    x"2F313F60",
    x"2F312939",
    x"2F311316",
    x"2F30FCF5",
    x"2F30E6D6",
    x"2F30D0BB",
    x"2F30BAA2",
    x"2F30A48C",
    x"2F308E79",
    x"2F307869",
    x"2F30625B",
    x"2F304C50",
    x"2F303648",
    x"2F302042",
    x"2F300A40",
    x"2F2FF440",
    x"2F2FDE43",
    x"2F2FC848",
    x"2F2FB251",
    x"2F2F9C5C",
    x"2F2F866A",
    x"2F2F707A",
    x"2F2F5A8D",
    x"2F2F44A3",
    x"2F2F2EBC",
    x"2F2F18D8",
    x"2F2F02F6",
    x"2F2EED17",
    x"2F2ED73B",
    x"2F2EC161",
    x"2F2EAB8A",
    x"2F2E95B6",
    x"2F2E7FE5",
    x"2F2E6A16",
    x"2F2E544A",
    x"2F2E3E81",
    x"2F2E28BB",
    x"2F2E12F7",
    x"2F2DFD36",
    x"2F2DE778",
    x"2F2DD1BC",
    x"2F2DBC03",
    x"2F2DA64D",
    x"2F2D909A",
    x"2F2D7AE9",
    x"2F2D653B",
    x"2F2D4F90",
    x"2F2D39E7",
    x"2F2D2441",
    x"2F2D0E9E",
    x"2F2CF8FE",
    x"2F2CE360",
    x"2F2CCDC5",
    x"2F2CB82C",
    x"2F2CA297",
    x"2F2C8D04",
    x"2F2C7773",
    x"2F2C61E6",
    x"2F2C4C5B",
    x"2F2C36D3",
    x"2F2C214D",
    x"2F2C0BCA",
    x"2F2BF64A",
    x"2F2BE0CD",
    x"2F2BCB52",
    x"2F2BB5DA",
    x"2F2BA065",
    x"2F2B8AF2",
    x"2F2B7582",
    x"2F2B6015",
    x"2F2B4AAA",
    x"2F2B3542",
    x"2F2B1FDD",
    x"2F2B0A7A",
    x"2F2AF51A",
    x"2F2ADFBD",
    x"2F2ACA62",
    x"2F2AB50A",
    x"2F2A9FB5",
    x"2F2A8A62",
    x"2F2A7512",
    x"2F2A5FC5",
    x"2F2A4A7A",
    x"2F2A3532",
    x"2F2A1FED",
    x"2F2A0AAA",
    x"2F29F56A",
    x"2F29E02D",
    x"2F29CAF2",
    x"2F29B5BA",
    x"2F29A085",
    x"2F298B52",
    x"2F297622",
    x"2F2960F5",
    x"2F294BCA",
    x"2F2936A2",
    x"2F29217C",
    x"2F290C59",
    x"2F28F739",
    x"2F28E21B",
    x"2F28CD00",
    x"2F28B7E8",
    x"2F28A2D3",
    x"2F288DBF",
    x"2F2878AF",
    x"2F2863A1",
    x"2F284E96",
    x"2F28398E",
    x"2F282488",
    x"2F280F85",
    x"2F27FA84",
    x"2F27E586",
    x"2F27D08B",
    x"2F27BB92",
    x"2F27A69C",
    x"2F2791A8",
    x"2F277CB7",
    x"2F2767C9",
    x"2F2752DD",
    x"2F273DF4",
    x"2F27290E",
    x"2F27142A",
    x"2F26FF49",
    x"2F26EA6A",
    x"2F26D58E",
    x"2F26C0B5",
    x"2F26ABDE",
    x"2F26970A",
    x"2F268238",
    x"2F266D69",
    x"2F26589D",
    x"2F2643D3",
    x"2F262F0C",
    x"2F261A47",
    x"2F260585",
    x"2F25F0C6",
    x"2F25DC09",
    x"2F25C74F",
    x"2F25B297",
    x"2F259DE2",
    x"2F258930",
    x"2F257480",
    x"2F255FD3",
    x"2F254B28",
    x"2F253680",
    x"2F2521DA",
    x"2F250D37",
    x"2F24F897",
    x"2F24E3F9",
    x"2F24CF5E",
    x"2F24BAC5",
    x"2F24A62F",
    x"2F24919C",
    x"2F247D0B",
    x"2F24687D",
    x"2F2453F1",
    x"2F243F68",
    x"2F242AE1",
    x"2F24165D",
    x"2F2401DB",
    x"2F23ED5C",
    x"2F23D8E0",
    x"2F23C466",
    x"2F23AFEF",
    x"2F239B7A",
    x"2F238708",
    x"2F237299",
    x"2F235E2B",
    x"2F2349C1",
    x"2F233559",
    x"2F2320F4",
    x"2F230C91",
    x"2F22F830",
    x"2F22E3D3",
    x"2F22CF78",
    x"2F22BB1F",
    x"2F22A6C9",
    x"2F229275",
    x"2F227E24",
    x"2F2269D6",
    x"2F22558A",
    x"2F224140",
    x"2F222CF9",
    x"2F2218B5",
    x"2F220473",
    x"2F21F034",
    x"2F21DBF7",
    x"2F21C7BD",
    x"2F21B385",
    x"2F219F50",
    x"2F218B1D",
    x"2F2176ED",
    x"2F2162C0",
    x"2F214E95",
    x"2F213A6C",
    x"2F212646",
    x"2F211222",
    x"2F20FE01",
    x"2F20E9E3",
    x"2F20D5C7",
    x"2F20C1AD",
    x"2F20AD97",
    x"2F209982",
    x"2F208570",
    x"2F207161",
    x"2F205D54",
    x"2F204949",
    x"2F203541",
    x"2F20213C",
    x"2F200D39",
    x"2F1FF939",
    x"2F1FE53B",
    x"2F1FD13F",
    x"2F1FBD47",
    x"2F1FA950",
    x"2F1F955C",
    x"2F1F816B",
    x"2F1F6D7C",
    x"2F1F598F",
    x"2F1F45A5",
    x"2F1F31BE",
    x"2F1F1DD9",
    x"2F1F09F7",
    x"2F1EF617",
    x"2F1EE239",
    x"2F1ECE5E",
    x"2F1EBA85",
    x"2F1EA6AF",
    x"2F1E92DC",
    x"2F1E7F0B",
    x"2F1E6B3C",
    x"2F1E5770",
    x"2F1E43A6",
    x"2F1E2FDF",
    x"2F1E1C1A",
    x"2F1E0858",
    x"2F1DF498",
    x"2F1DE0DB",
    x"2F1DCD20",
    x"2F1DB967",
    x"2F1DA5B2",
    x"2F1D91FE",
    x"2F1D7E4D",
    x"2F1D6A9E",
    x"2F1D56F2",
    x"2F1D4349",
    x"2F1D2FA2",
    x"2F1D1BFD",
    x"2F1D085B",
    x"2F1CF4BB",
    x"2F1CE11D",
    x"2F1CCD82",
    x"2F1CB9EA",
    x"2F1CA654",
    x"2F1C92C0",
    x"2F1C7F2F",
    x"2F1C6BA1",
    x"2F1C5814",
    x"2F1C448B",
    x"2F1C3103",
    x"2F1C1D7E",
    x"2F1C09FC",
    x"2F1BF67C",
    x"2F1BE2FE",
    x"2F1BCF83",
    x"2F1BBC0A",
    x"2F1BA894",
    x"2F1B9520",
    x"2F1B81AF",
    x"2F1B6E40",
    x"2F1B5AD3",
    x"2F1B4769",
    x"2F1B3401",
    x"2F1B209C",
    x"2F1B0D39",
    x"2F1AF9D9",
    x"2F1AE67B",
    x"2F1AD31F",
    x"2F1ABFC6",
    x"2F1AAC6F",
    x"2F1A991B",
    x"2F1A85C9",
    x"2F1A7279",
    x"2F1A5F2C",
    x"2F1A4BE2",
    x"2F1A3899",
    x"2F1A2553",
    x"2F1A1210",
    x"2F19FECF",
    x"2F19EB90",
    x"2F19D854",
    x"2F19C51A",
    x"2F19B1E3",
    x"2F199EAE",
    x"2F198B7B",
    x"2F19784B",
    x"2F19651D",
    x"2F1951F2",
    x"2F193EC9",
    x"2F192BA2",
    x"2F19187E",
    x"2F19055C",
    x"2F18F23C",
    x"2F18DF1F",
    x"2F18CC05",
    x"2F18B8EC",
    x"2F18A5D6",
    x"2F1892C3",
    x"2F187FB2",
    x"2F186CA3",
    x"2F185996",
    x"2F18468C",
    x"2F183385",
    x"2F182080",
    x"2F180D7D",
    x"2F17FA7C",
    x"2F17E77E",
    x"2F17D482",
    x"2F17C189",
    x"2F17AE92",
    x"2F179B9D",
    x"2F1788AB",
    x"2F1775BB",
    x"2F1762CE",
    x"2F174FE2",
    x"2F173CFA",
    x"2F172A13",
    x"2F17172F",
    x"2F17044D",
    x"2F16F16E",
    x"2F16DE91",
    x"2F16CBB6",
    x"2F16B8DE",
    x"2F16A608",
    x"2F169335",
    x"2F168063",
    x"2F166D95",
    x"2F165AC8",
    x"2F1647FE",
    x"2F163536",
    x"2F162271",
    x"2F160FAD",
    x"2F15FCED",
    x"2F15EA2E",
    x"2F15D772",
    x"2F15C4B8",
    x"2F15B201",
    x"2F159F4C",
    x"2F158C99",
    x"2F1579E9",
    x"2F15673B",
    x"2F15548F",
    x"2F1541E5",
    x"2F152F3E",
    x"2F151C9A",
    x"2F1509F7",
    x"2F14F757",
    x"2F14E4B9",
    x"2F14D21E",
    x"2F14BF85",
    x"2F14ACEE",
    x"2F149A5A",
    x"2F1487C7",
    x"2F147538",
    x"2F1462AA",
    x"2F14501F",
    x"2F143D96",
    x"2F142B10",
    x"2F14188B",
    x"2F140609",
    x"2F13F38A",
    x"2F13E10D",
    x"2F13CE92",
    x"2F13BC19",
    x"2F13A9A3",
    x"2F13972F",
    x"2F1384BD",
    x"2F13724D",
    x"2F135FE0",
    x"2F134D75",
    x"2F133B0D",
    x"2F1328A7",
    x"2F131643",
    x"2F1303E1",
    x"2F12F182",
    x"2F12DF25",
    x"2F12CCCA",
    x"2F12BA71",
    x"2F12A81B",
    x"2F1295C7",
    x"2F128376",
    x"2F127127",
    x"2F125EDA",
    x"2F124C8F",
    x"2F123A46",
    x"2F122800",
    x"2F1215BC",
    x"2F12037B",
    x"2F11F13C",
    x"2F11DEFF",
    x"2F11CCC4",
    x"2F11BA8B",
    x"2F11A855",
    x"2F119621",
    x"2F1183F0",
    x"2F1171C0",
    x"2F115F93",
    x"2F114D68",
    x"2F113B40",
    x"2F11291A",
    x"2F1116F6",
    x"2F1104D4",
    x"2F10F2B4",
    x"2F10E097",
    x"2F10CE7C",
    x"2F10BC64",
    x"2F10AA4D",
    x"2F109839",
    x"2F108627",
    x"2F107417",
    x"2F10620A",
    x"2F104FFF",
    x"2F103DF6",
    x"2F102BEF",
    x"2F1019EB",
    x"2F1007E9",
    x"2F0FF5E9",
    x"2F0FE3EB",
    x"2F0FD1F0",
    x"2F0FBFF7",
    x"2F0FAE00",
    x"2F0F9C0B",
    x"2F0F8A19",
    x"2F0F7829",
    x"2F0F663B",
    x"2F0F544F",
    x"2F0F4266",
    x"2F0F307F",
    x"2F0F1E9A",
    x"2F0F0CB7",
    x"2F0EFAD7",
    x"2F0EE8F8",
    x"2F0ED71C",
    x"2F0EC543",
    x"2F0EB36B",
    x"2F0EA196",
    x"2F0E8FC3",
    x"2F0E7DF2",
    x"2F0E6C23",
    x"2F0E5A57",
    x"2F0E488D",
    x"2F0E36C5",
    x"2F0E24FF",
    x"2F0E133B",
    x"2F0E017A",
    x"2F0DEFBB",
    x"2F0DDDFE",
    x"2F0DCC44",
    x"2F0DBA8B",
    x"2F0DA8D5",
    x"2F0D9721",
    x"2F0D856F",
    x"2F0D73C0",
    x"2F0D6212",
    x"2F0D5067",
    x"2F0D3EBE",
    x"2F0D2D17",
    x"2F0D1B73",
    x"2F0D09D1",
    x"2F0CF830",
    x"2F0CE692",
    x"2F0CD4F7",
    x"2F0CC35D",
    x"2F0CB1C6",
    x"2F0CA031",
    x"2F0C8E9E",
    x"2F0C7D0D",
    x"2F0C6B7F",
    x"2F0C59F2",
    x"2F0C4868",
    x"2F0C36E0",
    x"2F0C255A",
    x"2F0C13D7",
    x"2F0C0255",
    x"2F0BF0D6",
    x"2F0BDF59",
    x"2F0BCDDE",
    x"2F0BBC66",
    x"2F0BAAEF",
    x"2F0B997B",
    x"2F0B8809",
    x"2F0B7699",
    x"2F0B652B",
    x"2F0B53C0",
    x"2F0B4256",
    x"2F0B30EF",
    x"2F0B1F8A",
    x"2F0B0E27",
    x"2F0AFCC7",
    x"2F0AEB68",
    x"2F0ADA0C",
    x"2F0AC8B2",
    x"2F0AB75A",
    x"2F0AA604",
    x"2F0A94B0",
    x"2F0A835F",
    x"2F0A720F",
    x"2F0A60C2",
    x"2F0A4F77",
    x"2F0A3E2E",
    x"2F0A2CE7",
    x"2F0A1BA3",
    x"2F0A0A61",
    x"2F09F920",
    x"2F09E7E2",
    x"2F09D6A6",
    x"2F09C56D",
    x"2F09B435",
    x"2F09A300",
    x"2F0991CC",
    x"2F09809B",
    x"2F096F6C",
    x"2F095E3F",
    x"2F094D15",
    x"2F093BEC",
    x"2F092AC6",
    x"2F0919A1",
    x"2F09087F",
    x"2F08F75F",
    x"2F08E641",
    x"2F08D526",
    x"2F08C40C",
    x"2F08B2F5",
    x"2F08A1DF",
    x"2F0890CC",
    x"2F087FBB",
    x"2F086EAC",
    x"2F085D9F",
    x"2F084C95",
    x"2F083B8C",
    x"2F082A86",
    x"2F081982",
    x"2F080880",
    x"2F07F780",
    x"2F07E682",
    x"2F07D586",
    x"2F07C48C",
    x"2F07B395",
    x"2F07A29F",
    x"2F0791AC",
    x"2F0780BB",
    x"2F076FCC",
    x"2F075EDF",
    x"2F074DF4",
    x"2F073D0B",
    x"2F072C25",
    x"2F071B40",
    x"2F070A5E",
    x"2F06F97E",
    x"2F06E8A0",
    x"2F06D7C4",
    x"2F06C6EA",
    x"2F06B612",
    x"2F06A53C",
    x"2F069469",
    x"2F068397",
    x"2F0672C8",
    x"2F0661FA",
    x"2F06512F",
    x"2F064066",
    x"2F062F9F",
    x"2F061EDA",
    x"2F060E17",
    x"2F05FD57",
    x"2F05EC98",
    x"2F05DBDC",
    x"2F05CB21",
    x"2F05BA69",
    x"2F05A9B3",
    x"2F0598FE",
    x"2F05884C",
    x"2F05779C",
    x"2F0566EE",
    x"2F055643",
    x"2F054599",
    x"2F0534F1",
    x"2F05244C",
    x"2F0513A8",
    x"2F050307",
    x"2F04F267",
    x"2F04E1CA",
    x"2F04D12F",
    x"2F04C096",
    x"2F04AFFF",
    x"2F049F6A",
    x"2F048ED7",
    x"2F047E46",
    x"2F046DB7",
    x"2F045D2B",
    x"2F044CA0",
    x"2F043C18",
    x"2F042B91",
    x"2F041B0D",
    x"2F040A8A",
    x"2F03FA0A",
    x"2F03E98C",
    x"2F03D910",
    x"2F03C895",
    x"2F03B81D",
    x"2F03A7A7",
    x"2F039734",
    x"2F0386C2",
    x"2F037652",
    x"2F0365E4",
    x"2F035578",
    x"2F03450F",
    x"2F0334A7",
    x"2F032442",
    x"2F0313DE",
    x"2F03037D",
    x"2F02F31D",
    x"2F02E2C0",
    x"2F02D264",
    x"2F02C20B",
    x"2F02B1B4",
    x"2F02A15F",
    x"2F02910C",
    x"2F0280BB",
    x"2F02706B",
    x"2F02601E",
    x"2F024FD3",
    x"2F023F8A",
    x"2F022F44",
    x"2F021EFF",
    x"2F020EBC",
    x"2F01FE7B",
    x"2F01EE3C",
    x"2F01DDFF",
    x"2F01CDC5",
    x"2F01BD8C",
    x"2F01AD55",
    x"2F019D21",
    x"2F018CEE",
    x"2F017CBD",
    x"2F016C8F",
    x"2F015C62",
    x"2F014C38",
    x"2F013C0F",
    x"2F012BE9",
    x"2F011BC4",
    x"2F010BA2",
    x"2F00FB81",
    x"2F00EB63",
    x"2F00DB46",
    x"2F00CB2C",
    x"2F00BB14",
    x"2F00AAFD",
    x"2F009AE9",
    x"2F008AD7",
    x"2F007AC6",
    x"2F006AB8",
    x"2F005AAC",
    x"2F004AA1",
    x"2F003A99",
    x"2F002A93",
    x"2F001A8E",
    x"2F000A8C",
    x"2EFFF517",
    x"2EFFD51B",
    x"2EFFB522",
    x"2EFF952D",
    x"2EFF753D",
    x"2EFF5550",
    x"2EFF3567",
    x"2EFF1583",
    x"2EFEF5A2",
    x"2EFED5C5",
    x"2EFEB5EC",
    x"2EFE9618",
    x"2EFE7647",
    x"2EFE567A",
    x"2EFE36B1",
    x"2EFE16EC",
    x"2EFDF72C",
    x"2EFDD76F",
    x"2EFDB7B6",
    x"2EFD9801",
    x"2EFD7850",
    x"2EFD58A3",
    x"2EFD38FA",
    x"2EFD1954",
    x"2EFCF9B3",
    x"2EFCDA16",
    x"2EFCBA7D",
    x"2EFC9AE7",
    x"2EFC7B56",
    x"2EFC5BC9",
    x"2EFC3C3F",
    x"2EFC1CB9",
    x"2EFBFD38",
    x"2EFBDDBA",
    x"2EFBBE40",
    x"2EFB9ECB",
    x"2EFB7F59",
    x"2EFB5FEB",
    x"2EFB4081",
    x"2EFB211B",
    x"2EFB01B8",
    x"2EFAE25A",
    x"2EFAC300",
    x"2EFAA3A9",
    x"2EFA8457",
    x"2EFA6508",
    x"2EFA45BE",
    x"2EFA2677",
    x"2EFA0734",
    x"2EF9E7F5",
    x"2EF9C8BA",
    x"2EF9A983",
    x"2EF98A50",
    x"2EF96B20",
    x"2EF94BF5",
    x"2EF92CCD",
    x"2EF90DAA",
    x"2EF8EE8A",
    x"2EF8CF6E",
    x"2EF8B056",
    x"2EF89142",
    x"2EF87232",
    x"2EF85325",
    x"2EF8341D",
    x"2EF81518",
    x"2EF7F618",
    x"2EF7D71B",
    x"2EF7B822",
    x"2EF7992D",
    x"2EF77A3C",
    x"2EF75B4E",
    x"2EF73C65",
    x"2EF71D7F",
    x"2EF6FE9D",
    x"2EF6DFC0",
    x"2EF6C0E6",
    x"2EF6A20F",
    x"2EF6833D",
    x"2EF6646F",
    x"2EF645A4",
    x"2EF626DD",
    x"2EF6081A",
    x"2EF5E95B",
    x"2EF5CAA0",
    x"2EF5ABE8",
    x"2EF58D35",
    x"2EF56E85",
    x"2EF54FD9",
    x"2EF53131",
    x"2EF5128D",
    x"2EF4F3ED",
    x"2EF4D550",
    x"2EF4B6B7",
    x"2EF49822",
    x"2EF47991",
    x"2EF45B04",
    x"2EF43C7A",
    x"2EF41DF5",
    x"2EF3FF73",
    x"2EF3E0F5",
    x"2EF3C27B",
    x"2EF3A404",
    x"2EF38592",
    x"2EF36723",
    x"2EF348B8",
    x"2EF32A51",
    x"2EF30BED",
    x"2EF2ED8E",
    x"2EF2CF32",
    x"2EF2B0DA",
    x"2EF29286",
    x"2EF27435",
    x"2EF255E9",
    x"2EF237A0",
    x"2EF2195B",
    x"2EF1FB19",
    x"2EF1DCDC",
    x"2EF1BEA2",
    x"2EF1A06C",
    x"2EF1823A",
    x"2EF1640C",
    x"2EF145E1",
    x"2EF127BA",
    x"2EF10997",
    x"2EF0EB78",
    x"2EF0CD5C",
    x"2EF0AF45",
    x"2EF09131",
    x"2EF07320",
    x"2EF05514",
    x"2EF0370B",
    x"2EF01906",
    x"2EEFFB05",
    x"2EEFDD07",
    x"2EEFBF0D",
    x"2EEFA117",
    x"2EEF8325",
    x"2EEF6537",
    x"2EEF474C",
    x"2EEF2965",
    x"2EEF0B82",
    x"2EEEEDA2",
    x"2EEECFC6",
    x"2EEEB1EE",
    x"2EEE941A",
    x"2EEE7649",
    x"2EEE587C",
    x"2EEE3AB3",
    x"2EEE1CED",
    x"2EEDFF2C",
    x"2EEDE16E",
    x"2EEDC3B3",
    x"2EEDA5FD",
    x"2EED884A",
    x"2EED6A9B",
    x"2EED4CEF",
    x"2EED2F47",
    x"2EED11A3",
    x"2EECF403",
    x"2EECD666",
    x"2EECB8CD",
    x"2EEC9B38",
    x"2EEC7DA7",
    x"2EEC6019",
    x"2EEC428F",
    x"2EEC2508",
    x"2EEC0785",
    x"2EEBEA06",
    x"2EEBCC8B",
    x"2EEBAF13",
    x"2EEB919F",
    x"2EEB742F",
    x"2EEB56C2",
    x"2EEB3959",
    x"2EEB1BF4",
    x"2EEAFE92",
    x"2EEAE134",
    x"2EEAC3DA",
    x"2EEAA683",
    x"2EEA8930",
    x"2EEA6BE1",
    x"2EEA4E95",
    x"2EEA314D",
    x"2EEA1409",
    x"2EE9F6C8",
    x"2EE9D98B",
    x"2EE9BC52",
    x"2EE99F1C",
    x"2EE981EA",
    x"2EE964BB",
    x"2EE94791",
    x"2EE92A6A",
    x"2EE90D46",
    x"2EE8F026",
    x"2EE8D30A",
    x"2EE8B5F2",
    x"2EE898DD",
    x"2EE87BCB",
    x"2EE85EBE",
    x"2EE841B4",
    x"2EE824AD",
    x"2EE807AA",
    x"2EE7EAAB",
    x"2EE7CDB0",
    x"2EE7B0B8",
    x"2EE793C4",
    x"2EE776D3",
    x"2EE759E6",
    x"2EE73CFC",
    x"2EE72017",
    x"2EE70334",
    x"2EE6E656",
    x"2EE6C97B",
    x"2EE6ACA3",
    x"2EE68FD0",
    x"2EE67300",
    x"2EE65633",
    x"2EE6396A",
    x"2EE61CA5",
    x"2EE5FFE3",
    x"2EE5E325",
    x"2EE5C66A",
    x"2EE5A9B3",
    x"2EE58D00",
    x"2EE57050",
    x"2EE553A4",
    x"2EE536FB",
    x"2EE51A56",
    x"2EE4FDB4",
    x"2EE4E116",
    x"2EE4C47C",
    x"2EE4A7E5",
    x"2EE48B52",
    x"2EE46EC2",
    x"2EE45236",
    x"2EE435AE",
    x"2EE41929",
    x"2EE3FCA8",
    x"2EE3E02A",
    x"2EE3C3AF",
    x"2EE3A739",
    x"2EE38AC6",
    x"2EE36E56",
    x"2EE351EA",
    x"2EE33582",
    x"2EE3191D",
    x"2EE2FCBB",
    x"2EE2E05E",
    x"2EE2C403",
    x"2EE2A7AD",
    x"2EE28B59",
    x"2EE26F0A",
    x"2EE252BE",
    x"2EE23675",
    x"2EE21A30",
    x"2EE1FDEE",
    x"2EE1E1B0",
    x"2EE1C576",
    x"2EE1A93F",
    x"2EE18D0C",
    x"2EE170DC",
    x"2EE154B0",
    x"2EE13887",
    x"2EE11C61",
    x"2EE10040",
    x"2EE0E421",
    x"2EE0C807",
    x"2EE0ABEF",
    x"2EE08FDC",
    x"2EE073CB",
    x"2EE057BF",
    x"2EE03BB5",
    x"2EE01FB0",
    x"2EE003AD",
    x"2EDFE7AF",
    x"2EDFCBB4",
    x"2EDFAFBC",
    x"2EDF93C8",
    x"2EDF77D7",
    x"2EDF5BEA",
    x"2EDF4000",
    x"2EDF241A",
    x"2EDF0837",
    x"2EDEEC58",
    x"2EDED07C",
    x"2EDEB4A4",
    x"2EDE98CF",
    x"2EDE7CFD",
    x"2EDE612F",
    x"2EDE4565",
    x"2EDE299E",
    x"2EDE0DDB",
    x"2EDDF21B",
    x"2EDDD65E",
    x"2EDDBAA5",
    x"2EDD9EEF",
    x"2EDD833D",
    x"2EDD678F",
    x"2EDD4BE3",
    x"2EDD303C",
    x"2EDD1497",
    x"2EDCF8F6",
    x"2EDCDD59",
    x"2EDCC1BF",
    x"2EDCA629",
    x"2EDC8A96",
    x"2EDC6F06",
    x"2EDC537A",
    x"2EDC37F1",
    x"2EDC1C6C",
    x"2EDC00EA",
    x"2EDBE56C",
    x"2EDBC9F1",
    x"2EDBAE79",
    x"2EDB9305",
    x"2EDB7794",
    x"2EDB5C27",
    x"2EDB40BD",
    x"2EDB2557",
    x"2EDB09F4",
    x"2EDAEE94",
    x"2EDAD338",
    x"2EDAB7E0",
    x"2EDA9C8A",
    x"2EDA8139",
    x"2EDA65EA",
    x"2EDA4A9F",
    x"2EDA2F57",
    x"2EDA1413",
    x"2ED9F8D2",
    x"2ED9DD95",
    x"2ED9C25B",
    x"2ED9A724",
    x"2ED98BF1",
    x"2ED970C1",
    x"2ED95595",
    x"2ED93A6C",
    x"2ED91F46",
    x"2ED90424",
    x"2ED8E905",
    x"2ED8CDEA",
    x"2ED8B2D2",
    x"2ED897BD",
    x"2ED87CAC",
    x"2ED8619E",
    x"2ED84694",
    x"2ED82B8C",
    x"2ED81089",
    x"2ED7F588",
    x"2ED7DA8B",
    x"2ED7BF92",
    x"2ED7A49B",
    x"2ED789A9",
    x"2ED76EB9",
    x"2ED753CD",
    x"2ED738E4",
    x"2ED71DFF",
    x"2ED7031D",
    x"2ED6E83E",
    x"2ED6CD62",
    x"2ED6B28B",
    x"2ED697B6",
    x"2ED67CE5",
    x"2ED66217",
    x"2ED6474C",
    x"2ED62C85",
    x"2ED611C1",
    x"2ED5F700",
    x"2ED5DC43",
    x"2ED5C189",
    x"2ED5A6D3",
    x"2ED58C20",
    x"2ED57170",
    x"2ED556C3",
    x"2ED53C1A",
    x"2ED52174",
    x"2ED506D2",
    x"2ED4EC33",
    x"2ED4D197",
    x"2ED4B6FE",
    x"2ED49C69",
    x"2ED481D7",
    x"2ED46748",
    x"2ED44CBD",
    x"2ED43235",
    x"2ED417B1",
    x"2ED3FD2F",
    x"2ED3E2B1",
    x"2ED3C837",
    x"2ED3ADBF",
    x"2ED3934B",
    x"2ED378DA",
    x"2ED35E6D",
    x"2ED34403",
    x"2ED3299C",
    x"2ED30F38",
    x"2ED2F4D8",
    x"2ED2DA7B",
    x"2ED2C022",
    x"2ED2A5CB",
    x"2ED28B78",
    x"2ED27128",
    x"2ED256DC",
    x"2ED23C93",
    x"2ED2224D",
    x"2ED2080A",
    x"2ED1EDCB",
    x"2ED1D38F",
    x"2ED1B956",
    x"2ED19F20",
    x"2ED184EE",
    x"2ED16ABF",
    x"2ED15093",
    x"2ED1366B",
    x"2ED11C46",
    x"2ED10224",
    x"2ED0E805",
    x"2ED0CDEA",
    x"2ED0B3D2",
    x"2ED099BD",
    x"2ED07FAB",
    x"2ED0659D",
    x"2ED04B92",
    x"2ED0318A",
    x"2ED01785",
    x"2ECFFD84",
    x"2ECFE386",
    x"2ECFC98B",
    x"2ECFAF94",
    x"2ECF959F",
    x"2ECF7BAE",
    x"2ECF61C0",
    x"2ECF47D6",
    x"2ECF2DEF",
    x"2ECF140A",
    x"2ECEFA2A",
    x"2ECEE04C",
    x"2ECEC671",
    x"2ECEAC9A",
    x"2ECE92C6",
    x"2ECE78F6",
    x"2ECE5F28",
    x"2ECE455E",
    x"2ECE2B97",
    x"2ECE11D3",
    x"2ECDF812",
    x"2ECDDE55",
    x"2ECDC49B",
    x"2ECDAAE4",
    x"2ECD9130",
    x"2ECD777F",
    x"2ECD5DD2",
    x"2ECD4428",
    x"2ECD2A81",
    x"2ECD10DD",
    x"2ECCF73D",
    x"2ECCDD9F",
    x"2ECCC405",
    x"2ECCAA6E",
    x"2ECC90DB",
    x"2ECC774A",
    x"2ECC5DBD",
    x"2ECC4433",
    x"2ECC2AAC",
    x"2ECC1128",
    x"2ECBF7A8",
    x"2ECBDE2A",
    x"2ECBC4B0",
    x"2ECBAB39",
    x"2ECB91C5",
    x"2ECB7855",
    x"2ECB5EE7",
    x"2ECB457D",
    x"2ECB2C16",
    x"2ECB12B2",
    x"2ECAF951",
    x"2ECADFF4",
    x"2ECAC699",
    x"2ECAAD42",
    x"2ECA93EE",
    x"2ECA7A9D",
    x"2ECA614F",
    x"2ECA4805",
    x"2ECA2EBD",
    x"2ECA1579",
    x"2EC9FC38",
    x"2EC9E2FA",
    x"2EC9C9BF",
    x"2EC9B087",
    x"2EC99753",
    x"2EC97E22",
    x"2EC964F3",
    x"2EC94BC8",
    x"2EC932A0",
    x"2EC9197C",
    x"2EC9005A",
    x"2EC8E73C",
    x"2EC8CE20",
    x"2EC8B508",
    x"2EC89BF3",
    x"2EC882E1",
    x"2EC869D2",
    x"2EC850C7",
    x"2EC837BE",
    x"2EC81EB9",
    x"2EC805B6",
    x"2EC7ECB7",
    x"2EC7D3BB",
    x"2EC7BAC2",
    x"2EC7A1CD",
    x"2EC788DA",
    x"2EC76FEA",
    x"2EC756FE",
    x"2EC73E15",
    x"2EC7252E",
    x"2EC70C4B",
    x"2EC6F36B",
    x"2EC6DA8E",
    x"2EC6C1B5",
    x"2EC6A8DE",
    x"2EC6900A",
    x"2EC6773A",
    x"2EC65E6D",
    x"2EC645A2",
    x"2EC62CDB",
    x"2EC61417",
    x"2EC5FB56",
    x"2EC5E298",
    x"2EC5C9DE",
    x"2EC5B126",
    x"2EC59871",
    x"2EC57FC0",
    x"2EC56711",
    x"2EC54E66",
    x"2EC535BE",
    x"2EC51D19",
    x"2EC50476",
    x"2EC4EBD7",
    x"2EC4D33C",
    x"2EC4BAA3",
    x"2EC4A20D",
    x"2EC4897A",
    x"2EC470EA",
    x"2EC4585E",
    x"2EC43FD4",
    x"2EC4274E",
    x"2EC40ECB",
    x"2EC3F64A",
    x"2EC3DDCD",
    x"2EC3C553",
    x"2EC3ACDC",
    x"2EC39468",
    x"2EC37BF7",
    x"2EC36389",
    x"2EC34B1E",
    x"2EC332B6",
    x"2EC31A51",
    x"2EC301EF",
    x"2EC2E991",
    x"2EC2D135",
    x"2EC2B8DC",
    x"2EC2A087",
    x"2EC28834",
    x"2EC26FE5",
    x"2EC25798",
    x"2EC23F4F",
    x"2EC22708",
    x"2EC20EC5",
    x"2EC1F685",
    x"2EC1DE47",
    x"2EC1C60D",
    x"2EC1ADD6",
    x"2EC195A2",
    x"2EC17D70",
    x"2EC16542",
    x"2EC14D17",
    x"2EC134EF",
    x"2EC11CCA",
    x"2EC104A8",
    x"2EC0EC89",
    x"2EC0D46D",
    x"2EC0BC54",
    x"2EC0A43E",
    x"2EC08C2A",
    x"2EC0741A",
    x"2EC05C0D",
    x"2EC04403",
    x"2EC02BFC",
    x"2EC013F8",
    x"2EBFFBF7",
    x"2EBFE3F9",
    x"2EBFCBFE",
    x"2EBFB406",
    x"2EBF9C11",
    x"2EBF841F",
    x"2EBF6C30",
    x"2EBF5444",
    x"2EBF3C5B",
    x"2EBF2475",
    x"2EBF0C92",
    x"2EBEF4B2",
    x"2EBEDCD5",
    x"2EBEC4FB",
    x"2EBEAD24",
    x"2EBE9550",
    x"2EBE7D7E",
    x"2EBE65B0",
    x"2EBE4DE5",
    x"2EBE361D",
    x"2EBE1E58",
    x"2EBE0695",
    x"2EBDEED6",
    x"2EBDD71A",
    x"2EBDBF60",
    x"2EBDA7AA",
    x"2EBD8FF6",
    x"2EBD7846",
    x"2EBD6098",
    x"2EBD48EE",
    x"2EBD3146",
    x"2EBD19A1",
    x"2EBD01FF",
    x"2EBCEA61",
    x"2EBCD2C5",
    x"2EBCBB2C",
    x"2EBCA396",
    x"2EBC8C03",
    x"2EBC7473",
    x"2EBC5CE6",
    x"2EBC455C",
    x"2EBC2DD5",
    x"2EBC1650",
    x"2EBBFECF",
    x"2EBBE751",
    x"2EBBCFD5",
    x"2EBBB85D",
    x"2EBBA0E7",
    x"2EBB8975",
    x"2EBB7205",
    x"2EBB5A98",
    x"2EBB432E",
    x"2EBB2BC7",
    x"2EBB1463",
    x"2EBAFD02",
    x"2EBAE5A4",
    x"2EBACE49",
    x"2EBAB6F0",
    x"2EBA9F9B",
    x"2EBA8848",
    x"2EBA70F9",
    x"2EBA59AC",
    x"2EBA4262",
    x"2EBA2B1C",
    x"2EBA13D8",
    x"2EB9FC97",
    x"2EB9E559",
    x"2EB9CE1D",
    x"2EB9B6E5",
    x"2EB99FB0",
    x"2EB9887D",
    x"2EB9714E",
    x"2EB95A21",
    x"2EB942F7",
    x"2EB92BD0",
    x"2EB914AC",
    x"2EB8FD8B",
    x"2EB8E66D",
    x"2EB8CF51",
    x"2EB8B839",
    x"2EB8A123",
    x"2EB88A11",
    x"2EB87301",
    x"2EB85BF4",
    x"2EB844EA",
    x"2EB82DE3",
    x"2EB816DE",
    x"2EB7FFDD",
    x"2EB7E8DE",
    x"2EB7D1E3",
    x"2EB7BAEA",
    x"2EB7A3F4",
    x"2EB78D01",
    x"2EB77611",
    x"2EB75F23",
    x"2EB74839",
    x"2EB73151",
    x"2EB71A6D",
    x"2EB7038B",
    x"2EB6ECAC",
    x"2EB6D5CF",
    x"2EB6BEF6",
    x"2EB6A820",
    x"2EB6914C",
    x"2EB67A7B",
    x"2EB663AE",
    x"2EB64CE2",
    x"2EB6361A",
    x"2EB61F55",
    x"2EB60892",
    x"2EB5F1D3",
    x"2EB5DB16",
    x"2EB5C45C",
    x"2EB5ADA5",
    x"2EB596F1",
    x"2EB5803F",
    x"2EB56991",
    x"2EB552E5",
    x"2EB53C3C",
    x"2EB52596",
    x"2EB50EF2",
    x"2EB4F852",
    x"2EB4E1B4",
    x"2EB4CB1A",
    x"2EB4B482",
    x"2EB49DEC",
    x"2EB4875A",
    x"2EB470CB",
    x"2EB45A3E",
    x"2EB443B4",
    x"2EB42D2D",
    x"2EB416A9",
    x"2EB40027",
    x"2EB3E9A9",
    x"2EB3D32D",
    x"2EB3BCB4",
    x"2EB3A63E",
    x"2EB38FCA",
    x"2EB3795A",
    x"2EB362EC",
    x"2EB34C81",
    x"2EB33619",
    x"2EB31FB4",
    x"2EB30951",
    x"2EB2F2F1",
    x"2EB2DC94",
    x"2EB2C63A",
    x"2EB2AFE3",
    x"2EB2998E",
    x"2EB2833C",
    x"2EB26CED",
    x"2EB256A1",
    x"2EB24058",
    x"2EB22A11",
    x"2EB213CD",
    x"2EB1FD8C",
    x"2EB1E74E",
    x"2EB1D112",
    x"2EB1BAD9",
    x"2EB1A4A3",
    x"2EB18E70",
    x"2EB17840",
    x"2EB16212",
    x"2EB14BE7",
    x"2EB135BF",
    x"2EB11F9A",
    x"2EB10977",
    x"2EB0F358",
    x"2EB0DD3B",
    x"2EB0C720",
    x"2EB0B109",
    x"2EB09AF4",
    x"2EB084E2",
    x"2EB06ED3",
    x"2EB058C6",
    x"2EB042BD",
    x"2EB02CB6",
    x"2EB016B1",
    x"2EB000B0",
    x"2EAFEAB1",
    x"2EAFD4B5",
    x"2EAFBEBC",
    x"2EAFA8C6",
    x"2EAF92D2",
    x"2EAF7CE1",
    x"2EAF66F3",
    x"2EAF5107",
    x"2EAF3B1E",
    x"2EAF2538",
    x"2EAF0F55",
    x"2EAEF975",
    x"2EAEE397",
    x"2EAECDBC",
    x"2EAEB7E3",
    x"2EAEA20E",
    x"2EAE8C3B",
    x"2EAE766B",
    x"2EAE609D",
    x"2EAE4AD2",
    x"2EAE350A",
    x"2EAE1F45",
    x"2EAE0983",
    x"2EADF3C3",
    x"2EADDE06",
    x"2EADC84B",
    x"2EADB294",
    x"2EAD9CDF",
    x"2EAD872C",
    x"2EAD717D",
    x"2EAD5BD0",
    x"2EAD4626",
    x"2EAD307E",
    x"2EAD1ADA",
    x"2EAD0538",
    x"2EACEF98",
    x"2EACD9FC",
    x"2EACC462",
    x"2EACAECB",
    x"2EAC9936",
    x"2EAC83A4",
    x"2EAC6E15",
    x"2EAC5889",
    x"2EAC42FF",
    x"2EAC2D78",
    x"2EAC17F4",
    x"2EAC0272",
    x"2EABECF3",
    x"2EABD777",
    x"2EABC1FD",
    x"2EABAC86",
    x"2EAB9712",
    x"2EAB81A1",
    x"2EAB6C32",
    x"2EAB56C6",
    x"2EAB415C",
    x"2EAB2BF5",
    x"2EAB1691",
    x"2EAB0130",
    x"2EAAEBD1",
    x"2EAAD675",
    x"2EAAC11B",
    x"2EAAABC4",
    x"2EAA9670",
    x"2EAA811F",
    x"2EAA6BD0",
    x"2EAA5684",
    x"2EAA413A",
    x"2EAA2BF4",
    x"2EAA16AF",
    x"2EAA016E",
    x"2EA9EC2F",
    x"2EA9D6F3",
    x"2EA9C1B9",
    x"2EA9AC82",
    x"2EA9974E",
    x"2EA9821D",
    x"2EA96CEE",
    x"2EA957C1",
    x"2EA94298",
    x"2EA92D71",
    x"2EA9184C",
    x"2EA9032B",
    x"2EA8EE0C",
    x"2EA8D8EF",
    x"2EA8C3D5",
    x"2EA8AEBE",
    x"2EA899AA",
    x"2EA88498",
    x"2EA86F88",
    x"2EA85A7C",
    x"2EA84572",
    x"2EA8306A",
    x"2EA81B66",
    x"2EA80664",
    x"2EA7F164",
    x"2EA7DC67",
    x"2EA7C76D",
    x"2EA7B275",
    x"2EA79D80",
    x"2EA7888E",
    x"2EA7739E",
    x"2EA75EB1",
    x"2EA749C7",
    x"2EA734DF",
    x"2EA71FF9",
    x"2EA70B17",
    x"2EA6F637",
    x"2EA6E159",
    x"2EA6CC7E",
    x"2EA6B7A6",
    x"2EA6A2D0",
    x"2EA68DFD",
    x"2EA6792D",
    x"2EA6645F",
    x"2EA64F94",
    x"2EA63ACB",
    x"2EA62605",
    x"2EA61142",
    x"2EA5FC81",
    x"2EA5E7C3",
    x"2EA5D307",
    x"2EA5BE4E",
    x"2EA5A997",
    x"2EA594E3",
    x"2EA58032",
    x"2EA56B83",
    x"2EA556D7",
    x"2EA5422E",
    x"2EA52D87",
    x"2EA518E2",
    x"2EA50440",
    x"2EA4EFA1",
    x"2EA4DB04",
    x"2EA4C66A",
    x"2EA4B1D3",
    x"2EA49D3E",
    x"2EA488AC",
    x"2EA4741C",
    x"2EA45F8F",
    x"2EA44B04",
    x"2EA4367C",
    x"2EA421F6",
    x"2EA40D73",
    x"2EA3F8F3",
    x"2EA3E475",
    x"2EA3CFFA",
    x"2EA3BB81",
    x"2EA3A70B",
    x"2EA39297",
    x"2EA37E26",
    x"2EA369B8",
    x"2EA3554C",
    x"2EA340E2",
    x"2EA32C7C",
    x"2EA31817",
    x"2EA303B6",
    x"2EA2EF56",
    x"2EA2DAFA",
    x"2EA2C6A0",
    x"2EA2B248",
    x"2EA29DF3",
    x"2EA289A1",
    x"2EA27551",
    x"2EA26103",
    x"2EA24CB8",
    x"2EA23870",
    x"2EA2242A",
    x"2EA20FE7",
    x"2EA1FBA6",
    x"2EA1E768",
    x"2EA1D32C",
    x"2EA1BEF3",
    x"2EA1AABD",
    x"2EA19689",
    x"2EA18257",
    x"2EA16E28",
    x"2EA159FC",
    x"2EA145D2",
    x"2EA131AA",
    x"2EA11D85",
    x"2EA10963",
    x"2EA0F543",
    x"2EA0E125",
    x"2EA0CD0B",
    x"2EA0B8F2",
    x"2EA0A4DC",
    x"2EA090C9",
    x"2EA07CB8",
    x"2EA068AA",
    x"2EA0549E",
    x"2EA04095",
    x"2EA02C8E",
    x"2EA01889",
    x"2EA00488",
    x"2E9FF088",
    x"2E9FDC8C",
    x"2E9FC891",
    x"2E9FB499",
    x"2E9FA0A4",
    x"2E9F8CB1",
    x"2E9F78C1",
    x"2E9F64D3",
    x"2E9F50E8",
    x"2E9F3CFF",
    x"2E9F2918",
    x"2E9F1535",
    x"2E9F0153",
    x"2E9EED74",
    x"2E9ED998",
    x"2E9EC5BE",
    x"2E9EB1E6",
    x"2E9E9E11",
    x"2E9E8A3F",
    x"2E9E766F",
    x"2E9E62A1",
    x"2E9E4ED6",
    x"2E9E3B0D",
    x"2E9E2747",
    x"2E9E1384",
    x"2E9DFFC2",
    x"2E9DEC04",
    x"2E9DD847",
    x"2E9DC48E",
    x"2E9DB0D6",
    x"2E9D9D21",
    x"2E9D896F",
    x"2E9D75BF",
    x"2E9D6212",
    x"2E9D4E67",
    x"2E9D3ABE",
    x"2E9D2718",
    x"2E9D1374",
    x"2E9CFFD3",
    x"2E9CEC34",
    x"2E9CD898",
    x"2E9CC4FE",
    x"2E9CB167",
    x"2E9C9DD2",
    x"2E9C8A3F",
    x"2E9C76AF",
    x"2E9C6322",
    x"2E9C4F96",
    x"2E9C3C0E",
    x"2E9C2887",
    x"2E9C1504",
    x"2E9C0182",
    x"2E9BEE03",
    x"2E9BDA87",
    x"2E9BC70D",
    x"2E9BB395",
    x"2E9BA020",
    x"2E9B8CAD",
    x"2E9B793C",
    x"2E9B65CF",
    x"2E9B5263",
    x"2E9B3EFA",
    x"2E9B2B93",
    x"2E9B182F",
    x"2E9B04CD",
    x"2E9AF16E",
    x"2E9ADE11",
    x"2E9ACAB6",
    x"2E9AB75E",
    x"2E9AA409",
    x"2E9A90B5",
    x"2E9A7D64",
    x"2E9A6A16",
    x"2E9A56CA",
    x"2E9A4380",
    x"2E9A3039",
    x"2E9A1CF4",
    x"2E9A09B2",
    x"2E99F672",
    x"2E99E334",
    x"2E99CFF9",
    x"2E99BCC0",
    x"2E99A98A",
    x"2E999656",
    x"2E998324",
    x"2E996FF5",
    x"2E995CC8",
    x"2E99499E",
    x"2E993676",
    x"2E992350",
    x"2E99102D",
    x"2E98FD0C",
    x"2E98E9EE",
    x"2E98D6D2",
    x"2E98C3B8",
    x"2E98B0A1",
    x"2E989D8C",
    x"2E988A79",
    x"2E987769",
    x"2E98645B",
    x"2E985150",
    x"2E983E47",
    x"2E982B40",
    x"2E98183C",
    x"2E98053A",
    x"2E97F23B",
    x"2E97DF3E",
    x"2E97CC43",
    x"2E97B94B",
    x"2E97A655",
    x"2E979361",
    x"2E978070",
    x"2E976D81",
    x"2E975A95",
    x"2E9747AA",
    x"2E9734C3",
    x"2E9721DD",
    x"2E970EFA",
    x"2E96FC1A",
    x"2E96E93B",
    x"2E96D65F",
    x"2E96C386",
    x"2E96B0AE",
    x"2E969DD9",
    x"2E968B07",
    x"2E967837",
    x"2E966569",
    x"2E96529D",
    x"2E963FD4",
    x"2E962D0D",
    x"2E961A49",
    x"2E960787",
    x"2E95F4C7",
    x"2E95E20A",
    x"2E95CF4F",
    x"2E95BC96",
    x"2E95A9DF",
    x"2E95972B",
    x"2E95847A",
    x"2E9571CA",
    x"2E955F1D",
    x"2E954C72",
    x"2E9539CA",
    x"2E952724",
    x"2E951480",
    x"2E9501DF",
    x"2E94EF40",
    x"2E94DCA3",
    x"2E94CA09",
    x"2E94B771",
    x"2E94A4DB",
    x"2E949247",
    x"2E947FB6",
    x"2E946D27",
    x"2E945A9B",
    x"2E944811",
    x"2E943589",
    x"2E942303",
    x"2E941080",
    x"2E93FDFF",
    x"2E93EB81",
    x"2E93D904",
    x"2E93C68A",
    x"2E93B413",
    x"2E93A19D",
    x"2E938F2A",
    x"2E937CBA",
    x"2E936A4B",
    x"2E9357DF",
    x"2E934575",
    x"2E93330E",
    x"2E9320A8",
    x"2E930E45",
    x"2E92FBE5",
    x"2E92E986",
    x"2E92D72A",
    x"2E92C4D1",
    x"2E92B279",
    x"2E92A024",
    x"2E928DD1",
    x"2E927B81",
    x"2E926932",
    x"2E9256E6",
    x"2E92449D",
    x"2E923255",
    x"2E922010",
    x"2E920DCD",
    x"2E91FB8D",
    x"2E91E94E",
    x"2E91D712",
    x"2E91C4D8",
    x"2E91B2A1",
    x"2E91A06C",
    x"2E918E39",
    x"2E917C08",
    x"2E9169DA",
    x"2E9157AE",
    x"2E914584",
    x"2E91335C",
    x"2E912137",
    x"2E910F14",
    x"2E90FCF3",
    x"2E90EAD5",
    x"2E90D8B9",
    x"2E90C69F",
    x"2E90B487",
    x"2E90A272",
    x"2E90905E",
    x"2E907E4D",
    x"2E906C3F",
    x"2E905A32",
    x"2E904828",
    x"2E903620",
    x"2E90241B",
    x"2E901217",
    x"2E900016",
    x"2E8FEE17",
    x"2E8FDC1B",
    x"2E8FCA20",
    x"2E8FB828",
    x"2E8FA632",
    x"2E8F943F",
    x"2E8F824D",
    x"2E8F705E",
    x"2E8F5E71",
    x"2E8F4C86",
    x"2E8F3A9E",
    x"2E8F28B8",
    x"2E8F16D4",
    x"2E8F04F2",
    x"2E8EF313",
    x"2E8EE135",
    x"2E8ECF5A",
    x"2E8EBD81",
    x"2E8EABAB",
    x"2E8E99D7",
    x"2E8E8804",
    x"2E8E7635",
    x"2E8E6467",
    x"2E8E529B",
    x"2E8E40D2",
    x"2E8E2F0B",
    x"2E8E1D46",
    x"2E8E0B84",
    x"2E8DF9C4",
    x"2E8DE805",
    x"2E8DD64A",
    x"2E8DC490",
    x"2E8DB2D8",
    x"2E8DA123",
    x"2E8D8F70",
    x"2E8D7DBF",
    x"2E8D6C11",
    x"2E8D5A64",
    x"2E8D48BA",
    x"2E8D3712",
    x"2E8D256C",
    x"2E8D13C9",
    x"2E8D0227",
    x"2E8CF088",
    x"2E8CDEEB",
    x"2E8CCD50",
    x"2E8CBBB8",
    x"2E8CAA22",
    x"2E8C988D",
    x"2E8C86FB",
    x"2E8C756C",
    x"2E8C63DE",
    x"2E8C5253",
    x"2E8C40C9",
    x"2E8C2F42",
    x"2E8C1DBE",
    x"2E8C0C3B",
    x"2E8BFABB",
    x"2E8BE93C",
    x"2E8BD7C0",
    x"2E8BC646",
    x"2E8BB4CF",
    x"2E8BA359",
    x"2E8B91E6",
    x"2E8B8075",
    x"2E8B6F06",
    x"2E8B5D99",
    x"2E8B4C2E",
    x"2E8B3AC6",
    x"2E8B2960",
    x"2E8B17FC",
    x"2E8B069A",
    x"2E8AF53A",
    x"2E8AE3DC",
    x"2E8AD281",
    x"2E8AC128",
    x"2E8AAFD1",
    x"2E8A9E7C",
    x"2E8A8D29",
    x"2E8A7BD9",
    x"2E8A6A8A",
    x"2E8A593E",
    x"2E8A47F4",
    x"2E8A36AC",
    x"2E8A2566",
    x"2E8A1423",
    x"2E8A02E1",
    x"2E89F1A2",
    x"2E89E065",
    x"2E89CF2A",
    x"2E89BDF1",
    x"2E89ACBA",
    x"2E899B86",
    x"2E898A53",
    x"2E897923",
    x"2E8967F5",
    x"2E8956C9",
    x"2E89459F",
    x"2E893478",
    x"2E892352",
    x"2E89122F",
    x"2E89010E",
    x"2E88EFEF",
    x"2E88DED2",
    x"2E88CDB7",
    x"2E88BC9E",
    x"2E88AB88",
    x"2E889A73",
    x"2E888961",
    x"2E887851",
    x"2E886743",
    x"2E885637",
    x"2E88452E",
    x"2E883426",
    x"2E882321",
    x"2E88121D",
    x"2E88011C",
    x"2E87F01D",
    x"2E87DF20",
    x"2E87CE25",
    x"2E87BD2C",
    x"2E87AC36",
    x"2E879B41",
    x"2E878A4F",
    x"2E87795F",
    x"2E876871",
    x"2E875785",
    x"2E87469B",
    x"2E8735B3",
    x"2E8724CD",
    x"2E8713EA",
    x"2E870308",
    x"2E86F229",
    x"2E86E14C",
    x"2E86D071",
    x"2E86BF98",
    x"2E86AEC1",
    x"2E869DEC",
    x"2E868D19",
    x"2E867C49",
    x"2E866B7A",
    x"2E865AAE",
    x"2E8649E4",
    x"2E86391B",
    x"2E862855",
    x"2E861791",
    x"2E8606CF",
    x"2E85F610",
    x"2E85E552",
    x"2E85D496",
    x"2E85C3DD",
    x"2E85B325",
    x"2E85A270",
    x"2E8591BD",
    x"2E85810C",
    x"2E85705C",
    x"2E855FAF",
    x"2E854F05",
    x"2E853E5C",
    x"2E852DB5",
    x"2E851D10",
    x"2E850C6E",
    x"2E84FBCD",
    x"2E84EB2F",
    x"2E84DA92",
    x"2E84C9F8",
    x"2E84B960",
    x"2E84A8CA",
    x"2E849836",
    x"2E8487A4",
    x"2E847714",
    x"2E846686",
    x"2E8455FA",
    x"2E844570",
    x"2E8434E9",
    x"2E842463",
    x"2E8413E0",
    x"2E84035E",
    x"2E83F2DF",
    x"2E83E262",
    x"2E83D1E6",
    x"2E83C16D",
    x"2E83B0F6",
    x"2E83A081",
    x"2E83900E",
    x"2E837F9D",
    x"2E836F2E",
    x"2E835EC1",
    x"2E834E56",
    x"2E833DED",
    x"2E832D87",
    x"2E831D22",
    x"2E830CBF",
    x"2E82FC5F",
    x"2E82EC00",
    x"2E82DBA4",
    x"2E82CB49",
    x"2E82BAF1",
    x"2E82AA9B",
    x"2E829A46",
    x"2E8289F4",
    x"2E8279A4",
    x"2E826956",
    x"2E82590A",
    x"2E8248BF",
    x"2E823877",
    x"2E822831",
    x"2E8217ED",
    x"2E8207AB",
    x"2E81F76B",
    x"2E81E72D",
    x"2E81D6F2",
    x"2E81C6B8",
    x"2E81B680",
    x"2E81A64A",
    x"2E819616",
    x"2E8185E5",
    x"2E8175B5",
    x"2E816587",
    x"2E81555B",
    x"2E814532",
    x"2E81350A",
    x"2E8124E5",
    x"2E8114C1",
    x"2E81049F",
    x"2E80F480",
    x"2E80E462",
    x"2E80D447",
    x"2E80C42D",
    x"2E80B416",
    x"2E80A400",
    x"2E8093ED",
    x"2E8083DB",
    x"2E8073CC",
    x"2E8063BE",
    x"2E8053B3",
    x"2E8043A9",
    x"2E8033A2",
    x"2E80239C",
    x"2E801399",
    x"2E800398",
    x"2E7FE730",
    x"2E7FC735",
    x"2E7FA73E",
    x"2E7F874B",
    x"2E7F675C",
    x"2E7F4772",
    x"2E7F278B",
    x"2E7F07A8",
    x"2E7EE7C9",
    x"2E7EC7EE",
    x"2E7EA817",
    x"2E7E8844",
    x"2E7E6875",
    x"2E7E48AA",
    x"2E7E28E2",
    x"2E7E091F",
    x"2E7DE960",
    x"2E7DC9A5",
    x"2E7DA9EE",
    x"2E7D8A3B",
    x"2E7D6A8B",
    x"2E7D4AE0",
    x"2E7D2B39",
    x"2E7D0B95",
    x"2E7CEBF6",
    x"2E7CCC5A",
    x"2E7CACC3",
    x"2E7C8D2F",
    x"2E7C6D9F",
    x"2E7C4E14",
    x"2E7C2E8C",
    x"2E7C0F08",
    x"2E7BEF88",
    x"2E7BD00C",
    x"2E7BB094",
    x"2E7B9120",
    x"2E7B71B0",
    x"2E7B5243",
    x"2E7B32DB",
    x"2E7B1377",
    x"2E7AF416",
    x"2E7AD4BA",
    x"2E7AB561",
    x"2E7A960C",
    x"2E7A76BC",
    x"2E7A576F",
    x"2E7A3826",
    x"2E7A18E1",
    x"2E79F99F",
    x"2E79DA62",
    x"2E79BB29",
    x"2E799BF3",
    x"2E797CC2",
    x"2E795D94",
    x"2E793E6A",
    x"2E791F45",
    x"2E790023",
    x"2E78E105",
    x"2E78C1EA",
    x"2E78A2D4",
    x"2E7883C2",
    x"2E7864B3",
    x"2E7845A9",
    x"2E7826A2",
    x"2E78079F",
    x"2E77E8A0",
    x"2E77C9A5",
    x"2E77AAAD",
    x"2E778BBA",
    x"2E776CCB",
    x"2E774DDF",
    x"2E772EF7",
    x"2E771013",
    x"2E76F133",
    x"2E76D257",
    x"2E76B37E",
    x"2E7694AA",
    x"2E7675D9",
    x"2E76570C",
    x"2E763844",
    x"2E76197E",
    x"2E75FABD",
    x"2E75DC00",
    x"2E75BD46",
    x"2E759E90",
    x"2E757FDE",
    x"2E756130",
    x"2E754286",
    x"2E7523E0",
    x"2E75053D",
    x"2E74E69E",
    x"2E74C804",
    x"2E74A96C",
    x"2E748AD9",
    x"2E746C4A",
    x"2E744DBE",
    x"2E742F36",
    x"2E7410B2",
    x"2E73F232",
    x"2E73D3B6",
    x"2E73B53D",
    x"2E7396C8",
    x"2E737858",
    x"2E7359EA",
    x"2E733B81",
    x"2E731D1C",
    x"2E72FEBA",
    x"2E72E05C",
    x"2E72C202",
    x"2E72A3AB",
    x"2E728559",
    x"2E72670A",
    x"2E7248BF",
    x"2E722A78",
    x"2E720C34",
    x"2E71EDF5",
    x"2E71CFB9",
    x"2E71B181",
    x"2E71934D",
    x"2E71751C",
    x"2E7156EF",
    x"2E7138C6",
    x"2E711AA1",
    x"2E70FC80",
    x"2E70DE62",
    x"2E70C048",
    x"2E70A232",
    x"2E70841F",
    x"2E706611",
    x"2E704806",
    x"2E7029FF",
    x"2E700BFB",
    x"2E6FEDFC",
    x"2E6FD000",
    x"2E6FB208",
    x"2E6F9413",
    x"2E6F7623",
    x"2E6F5836",
    x"2E6F3A4D",
    x"2E6F1C67",
    x"2E6EFE86",
    x"2E6EE0A8",
    x"2E6EC2CD",
    x"2E6EA4F7",
    x"2E6E8724",
    x"2E6E6955",
    x"2E6E4B8A",
    x"2E6E2DC2",
    x"2E6E0FFE",
    x"2E6DF23E",
    x"2E6DD482",
    x"2E6DB6C9",
    x"2E6D9914",
    x"2E6D7B63",
    x"2E6D5DB5",
    x"2E6D400C",
    x"2E6D2265",
    x"2E6D04C3",
    x"2E6CE724",
    x"2E6CC989",
    x"2E6CABF2",
    x"2E6C8E5E",
    x"2E6C70CE",
    x"2E6C5342",
    x"2E6C35B9",
    x"2E6C1834",
    x"2E6BFAB3",
    x"2E6BDD36",
    x"2E6BBFBC",
    x"2E6BA246",
    x"2E6B84D3",
    x"2E6B6765",
    x"2E6B49FA",
    x"2E6B2C92",
    x"2E6B0F2E",
    x"2E6AF1CE",
    x"2E6AD472",
    x"2E6AB719",
    x"2E6A99C4",
    x"2E6A7C73",
    x"2E6A5F25",
    x"2E6A41DB",
    x"2E6A2495",
    x"2E6A0752",
    x"2E69EA13",
    x"2E69CCD7",
    x"2E69AFA0",
    x"2E69926B",
    x"2E69753B",
    x"2E69580E",
    x"2E693AE5",
    x"2E691DBF",
    x"2E69009E",
    x"2E68E37F",
    x"2E68C665",
    x"2E68A94E",
    x"2E688C3A",
    x"2E686F2B",
    x"2E68521F",
    x"2E683516",
    x"2E681811",
    x"2E67FB10",
    x"2E67DE13",
    x"2E67C119",
    x"2E67A422",
    x"2E678730",
    x"2E676A40",
    x"2E674D55",
    x"2E67306D",
    x"2E671389",
    x"2E66F6A8",
    x"2E66D9CB",
    x"2E66BCF2",
    x"2E66A01C",
    x"2E66834A",
    x"2E66667B",
    x"2E6649B0",
    x"2E662CE9",
    x"2E661025",
    x"2E65F365",
    x"2E65D6A8",
    x"2E65B9EF",
    x"2E659D3A",
    x"2E658088",
    x"2E6563D9",
    x"2E65472F",
    x"2E652A88",
    x"2E650DE4",
    x"2E64F144",
    x"2E64D4A8",
    x"2E64B80F",
    x"2E649B7A",
    x"2E647EE8",
    x"2E64625A",
    x"2E6445D0",
    x"2E642949",
    x"2E640CC5",
    x"2E63F045",
    x"2E63D3C9",
    x"2E63B750",
    x"2E639ADB",
    x"2E637E6A",
    x"2E6361FC",
    x"2E634591",
    x"2E63292A",
    x"2E630CC7",
    x"2E62F067",
    x"2E62D40B",
    x"2E62B7B2",
    x"2E629B5D",
    x"2E627F0B",
    x"2E6262BD",
    x"2E624673",
    x"2E622A2C",
    x"2E620DE8",
    x"2E61F1A8",
    x"2E61D56C",
    x"2E61B933",
    x"2E619CFD",
    x"2E6180CB",
    x"2E61649D",
    x"2E614872",
    x"2E612C4B",
    x"2E611027",
    x"2E60F407",
    x"2E60D7EA",
    x"2E60BBD1",
    x"2E609FBB",
    x"2E6083A9",
    x"2E60679A",
    x"2E604B8F",
    x"2E602F87",
    x"2E601383",
    x"2E5FF783",
    x"2E5FDB85",
    x"2E5FBF8C",
    x"2E5FA396",
    x"2E5F87A3",
    x"2E5F6BB4",
    x"2E5F4FC8",
    x"2E5F33E0",
    x"2E5F17FB",
    x"2E5EFC1A",
    x"2E5EE03C",
    x"2E5EC462",
    x"2E5EA88B",
    x"2E5E8CB7",
    x"2E5E70E8",
    x"2E5E551B",
    x"2E5E3952",
    x"2E5E1D8D",
    x"2E5E01CB",
    x"2E5DE60C",
    x"2E5DCA51",
    x"2E5DAE9A",
    x"2E5D92E6",
    x"2E5D7735",
    x"2E5D5B88",
    x"2E5D3FDE",
    x"2E5D2438",
    x"2E5D0895",
    x"2E5CECF6",
    x"2E5CD15A",
    x"2E5CB5C2",
    x"2E5C9A2D",
    x"2E5C7E9B",
    x"2E5C630D",
    x"2E5C4782",
    x"2E5C2BFB",
    x"2E5C1077",
    x"2E5BF4F7",
    x"2E5BD97A",
    x"2E5BBE01",
    x"2E5BA28A",
    x"2E5B8718",
    x"2E5B6BA9",
    x"2E5B503D",
    x"2E5B34D5",
    x"2E5B1970",
    x"2E5AFE0E",
    x"2E5AE2B0",
    x"2E5AC756",
    x"2E5AABFE",
    x"2E5A90AB",
    x"2E5A755A",
    x"2E5A5A0D",
    x"2E5A3EC4",
    x"2E5A237E",
    x"2E5A083B",
    x"2E59ECFC",
    x"2E59D1C0",
    x"2E59B687",
    x"2E599B52",
    x"2E598020",
    x"2E5964F2",
    x"2E5949C7",
    x"2E592EA0",
    x"2E59137B",
    x"2E58F85B",
    x"2E58DD3D",
    x"2E58C223",
    x"2E58A70D",
    x"2E588BFA",
    x"2E5870EA",
    x"2E5855DD",
    x"2E583AD4",
    x"2E581FCF",
    x"2E5804CC",
    x"2E57E9CD",
    x"2E57CED2",
    x"2E57B3DA",
    x"2E5798E5",
    x"2E577DF4",
    x"2E576305",
    x"2E57481B",
    x"2E572D33",
    x"2E57124F",
    x"2E56F76F",
    x"2E56DC92",
    x"2E56C1B8",
    x"2E56A6E1",
    x"2E568C0E",
    x"2E56713E",
    x"2E565672",
    x"2E563BA9",
    x"2E5620E3",
    x"2E560620",
    x"2E55EB61",
    x"2E55D0A5",
    x"2E55B5ED",
    x"2E559B38",
    x"2E558086",
    x"2E5565D8",
    x"2E554B2D",
    x"2E553085",
    x"2E5515E1",
    x"2E54FB40",
    x"2E54E0A2",
    x"2E54C607",
    x"2E54AB70",
    x"2E5490DD",
    x"2E54764C",
    x"2E545BBF",
    x"2E544135",
    x"2E5426AF",
    x"2E540C2C",
    x"2E53F1AC",
    x"2E53D72F",
    x"2E53BCB6",
    x"2E53A240",
    x"2E5387CD",
    x"2E536D5E",
    x"2E5352F2",
    x"2E533889",
    x"2E531E24",
    x"2E5303C2",
    x"2E52E963",
    x"2E52CF07",
    x"2E52B4AF",
    x"2E529A5A",
    x"2E528009",
    x"2E5265BA",
    x"2E524B6F",
    x"2E523127",
    x"2E5216E3",
    x"2E51FCA2",
    x"2E51E264",
    x"2E51C829",
    x"2E51ADF2",
    x"2E5193BD",
    x"2E51798D",
    x"2E515F5F",
    x"2E514535",
    x"2E512B0E",
    x"2E5110EA",
    x"2E50F6CA",
    x"2E50DCAC",
    x"2E50C292",
    x"2E50A87C",
    x"2E508E68",
    x"2E507458",
    x"2E505A4B",
    x"2E504042",
    x"2E50263B",
    x"2E500C38",
    x"2E4FF238",
    x"2E4FD83B",
    x"2E4FBE42",
    x"2E4FA44C",
    x"2E4F8A59",
    x"2E4F7069",
    x"2E4F567D",
    x"2E4F3C94",
    x"2E4F22AE",
    x"2E4F08CB",
    x"2E4EEEEC",
    x"2E4ED50F",
    x"2E4EBB36",
    x"2E4EA160",
    x"2E4E878E",
    x"2E4E6DBF",
    x"2E4E53F2",
    x"2E4E3A2A",
    x"2E4E2064",
    x"2E4E06A1",
    x"2E4DECE2",
    x"2E4DD326",
    x"2E4DB96D",
    x"2E4D9FB8",
    x"2E4D8606",
    x"2E4D6C56",
    x"2E4D52AA",
    x"2E4D3902",
    x"2E4D1F5C",
    x"2E4D05BA",
    x"2E4CEC1B",
    x"2E4CD27F",
    x"2E4CB8E6",
    x"2E4C9F51",
    x"2E4C85BE",
    x"2E4C6C2F",
    x"2E4C52A3",
    x"2E4C391B",
    x"2E4C1F95",
    x"2E4C0613",
    x"2E4BEC93",
    x"2E4BD317",
    x"2E4BB99F",
    x"2E4BA029",
    x"2E4B86B7",
    x"2E4B6D47",
    x"2E4B53DB",
    x"2E4B3A72",
    x"2E4B210D",
    x"2E4B07AA",
    x"2E4AEE4B",
    x"2E4AD4EF",
    x"2E4ABB96",
    x"2E4AA240",
    x"2E4A88ED",
    x"2E4A6F9D",
    x"2E4A5651",
    x"2E4A3D08",
    x"2E4A23C2",
    x"2E4A0A7F",
    x"2E49F13F",
    x"2E49D803",
    x"2E49BEC9",
    x"2E49A593",
    x"2E498C60",
    x"2E497330",
    x"2E495A03",
    x"2E4940D9",
    x"2E4927B3",
    x"2E490E8F",
    x"2E48F56F",
    x"2E48DC52",
    x"2E48C338",
    x"2E48AA21",
    x"2E48910E",
    x"2E4877FD",
    x"2E485EF0",
    x"2E4845E5",
    x"2E482CDE",
    x"2E4813DA",
    x"2E47FAD9",
    x"2E47E1DB",
    x"2E47C8E1",
    x"2E47AFE9",
    x"2E4796F5",
    x"2E477E03",
    x"2E476515",
    x"2E474C2A",
    x"2E473342",
    x"2E471A5D",
    x"2E47017C",
    x"2E46E89D",
    x"2E46CFC1",
    x"2E46B6E9",
    x"2E469E14",
    x"2E468541",
    x"2E466C72",
    x"2E4653A6",
    x"2E463ADD",
    x"2E462218",
    x"2E460955",
    x"2E45F095",
    x"2E45D7D9",
    x"2E45BF1F",
    x"2E45A669",
    x"2E458DB6",
    x"2E457506",
    x"2E455C58",
    x"2E4543AE",
    x"2E452B08",
    x"2E451264",
    x"2E44F9C3",
    x"2E44E125",
    x"2E44C88B",
    x"2E44AFF3",
    x"2E44975F",
    x"2E447ECD",
    x"2E44663F",
    x"2E444DB4",
    x"2E44352C",
    x"2E441CA6",
    x"2E440424",
    x"2E43EBA5",
    x"2E43D329",
    x"2E43BAB1",
    x"2E43A23B",
    x"2E4389C8",
    x"2E437158",
    x"2E4358EC",
    x"2E434082",
    x"2E43281C",
    x"2E430FB8",
    x"2E42F758",
    x"2E42DEFA",
    x"2E42C6A0",
    x"2E42AE49",
    x"2E4295F4",
    x"2E427DA3",
    x"2E426555",
    x"2E424D0A",
    x"2E4234C2",
    x"2E421C7D",
    x"2E42043B",
    x"2E41EBFC",
    x"2E41D3C0",
    x"2E41BB87",
    x"2E41A351",
    x"2E418B1E",
    x"2E4172EE",
    x"2E415AC1",
    x"2E414297",
    x"2E412A70",
    x"2E41124D",
    x"2E40FA2C",
    x"2E40E20E",
    x"2E40C9F3",
    x"2E40B1DC",
    x"2E4099C7",
    x"2E4081B5",
    x"2E4069A6",
    x"2E40519B",
    x"2E403992",
    x"2E40218C",
    x"2E40098A",
    x"2E3FF18A",
    x"2E3FD98D",
    x"2E3FC194",
    x"2E3FA99D",
    x"2E3F91A9",
    x"2E3F79B8",
    x"2E3F61CB",
    x"2E3F49E0",
    x"2E3F31F8",
    x"2E3F1A13",
    x"2E3F0232",
    x"2E3EEA53",
    x"2E3ED277",
    x"2E3EBA9E",
    x"2E3EA2C8",
    x"2E3E8AF6",
    x"2E3E7326",
    x"2E3E5B59",
    x"2E3E438F",
    x"2E3E2BC8",
    x"2E3E1404",
    x"2E3DFC43",
    x"2E3DE485",
    x"2E3DCCCA",
    x"2E3DB512",
    x"2E3D9D5D",
    x"2E3D85AA",
    x"2E3D6DFB",
    x"2E3D564F",
    x"2E3D3EA6",
    x"2E3D26FF",
    x"2E3D0F5C",
    x"2E3CF7BB",
    x"2E3CE01E",
    x"2E3CC883",
    x"2E3CB0EC",
    x"2E3C9957",
    x"2E3C81C5",
    x"2E3C6A37",
    x"2E3C52AB",
    x"2E3C3B22",
    x"2E3C239C",
    x"2E3C0C19",
    x"2E3BF499",
    x"2E3BDD1C",
    x"2E3BC5A2",
    x"2E3BAE2B",
    x"2E3B96B6",
    x"2E3B7F45",
    x"2E3B67D6",
    x"2E3B506B",
    x"2E3B3902",
    x"2E3B219D",
    x"2E3B0A3A",
    x"2E3AF2DA",
    x"2E3ADB7D",
    x"2E3AC423",
    x"2E3AACCC",
    x"2E3A9578",
    x"2E3A7E27",
    x"2E3A66D8",
    x"2E3A4F8D",
    x"2E3A3845",
    x"2E3A20FF",
    x"2E3A09BC",
    x"2E39F27D",
    x"2E39DB40",
    x"2E39C406",
    x"2E39ACCF",
    x"2E39959B",
    x"2E397E69",
    x"2E39673B",
    x"2E39500F",
    x"2E3938E7",
    x"2E3921C1",
    x"2E390A9E",
    x"2E38F37F",
    x"2E38DC62",
    x"2E38C548",
    x"2E38AE30",
    x"2E38971C",
    x"2E38800B",
    x"2E3868FC",
    x"2E3851F0",
    x"2E383AE7",
    x"2E3823E2",
    x"2E380CDF",
    x"2E37F5DE",
    x"2E37DEE1",
    x"2E37C7E7",
    x"2E37B0EF",
    x"2E3799FA",
    x"2E378309",
    x"2E376C1A",
    x"2E37552E",
    x"2E373E44",
    x"2E37275E",
    x"2E37107A",
    x"2E36F99A",
    x"2E36E2BC",
    x"2E36CBE1",
    x"2E36B509",
    x"2E369E34",
    x"2E368762",
    x"2E367092",
    x"2E3659C5",
    x"2E3642FC",
    x"2E362C35",
    x"2E361571",
    x"2E35FEAF",
    x"2E35E7F1",
    x"2E35D135",
    x"2E35BA7D",
    x"2E35A3C7",
    x"2E358D14",
    x"2E357663",
    x"2E355FB6",
    x"2E35490C",
    x"2E353264",
    x"2E351BBF",
    x"2E35051D",
    x"2E34EE7E",
    x"2E34D7E1",
    x"2E34C148",
    x"2E34AAB1",
    x"2E34941D",
    x"2E347D8C",
    x"2E3466FE",
    x"2E345072",
    x"2E3439E9",
    x"2E342364",
    x"2E340CE1",
    x"2E33F660",
    x"2E33DFE3",
    x"2E33C968",
    x"2E33B2F1",
    x"2E339C7C",
    x"2E33860A",
    x"2E336F9A",
    x"2E33592E",
    x"2E3342C4",
    x"2E332C5D",
    x"2E3315F9",
    x"2E32FF97",
    x"2E32E939",
    x"2E32D2DD",
    x"2E32BC84",
    x"2E32A62E",
    x"2E328FDB",
    x"2E32798A",
    x"2E32633C",
    x"2E324CF1",
    x"2E3236A9",
    x"2E322064",
    x"2E320A21",
    x"2E31F3E1",
    x"2E31DDA4",
    x"2E31C76A",
    x"2E31B132",
    x"2E319AFD",
    x"2E3184CB",
    x"2E316E9C",
    x"2E315870",
    x"2E314246",
    x"2E312C1F",
    x"2E3115FB",
    x"2E30FFDA",
    x"2E30E9BB",
    x"2E30D39F",
    x"2E30BD86",
    x"2E30A770",
    x"2E30915C",
    x"2E307B4C",
    x"2E30653D",
    x"2E304F32",
    x"2E30392A",
    x"2E302324",
    x"2E300D21",
    x"2E2FF721",
    x"2E2FE123",
    x"2E2FCB28",
    x"2E2FB530",
    x"2E2F9F3B",
    x"2E2F8949",
    x"2E2F7359",
    x"2E2F5D6C",
    x"2E2F4781",
    x"2E2F319A",
    x"2E2F1BB5",
    x"2E2F05D3",
    x"2E2EEFF4",
    x"2E2EDA17",
    x"2E2EC43D",
    x"2E2EAE66",
    x"2E2E9891",
    x"2E2E82C0",
    x"2E2E6CF1",
    x"2E2E5724",
    x"2E2E415B",
    x"2E2E2B94",
    x"2E2E15D0",
    x"2E2E000F",
    x"2E2DEA50",
    x"2E2DD494",
    x"2E2DBEDB",
    x"2E2DA924",
    x"2E2D9371",
    x"2E2D7DBF",
    x"2E2D6811",
    x"2E2D5265",
    x"2E2D3CBD",
    x"2E2D2716",
    x"2E2D1173",
    x"2E2CFBD2",
    x"2E2CE634",
    x"2E2CD098",
    x"2E2CBB00",
    x"2E2CA56A",
    x"2E2C8FD6",
    x"2E2C7A46",
    x"2E2C64B8",
    x"2E2C4F2C",
    x"2E2C39A4",
    x"2E2C241E",
    x"2E2C0E9B",
    x"2E2BF91A",
    x"2E2BE39D",
    x"2E2BCE22",
    x"2E2BB8A9",
    x"2E2BA333",
    x"2E2B8DC0",
    x"2E2B7850",
    x"2E2B62E2",
    x"2E2B4D77",
    x"2E2B380F",
    x"2E2B22A9",
    x"2E2B0D46",
    x"2E2AF7E6",
    x"2E2AE288",
    x"2E2ACD2D",
    x"2E2AB7D5",
    x"2E2AA27F",
    x"2E2A8D2C",
    x"2E2A77DC",
    x"2E2A628E",
    x"2E2A4D43",
    x"2E2A37FB",
    x"2E2A22B5",
    x"2E2A0D72",
    x"2E29F832",
    x"2E29E2F4",
    x"2E29CDB9",
    x"2E29B881",
    x"2E29A34B",
    x"2E298E18",
    x"2E2978E8",
    x"2E2963BA",
    x"2E294E8F",
    x"2E293966",
    x"2E292440",
    x"2E290F1D",
    x"2E28F9FD",
    x"2E28E4DF",
    x"2E28CFC3",
    x"2E28BAAB",
    x"2E28A595",
    x"2E289081",
    x"2E287B71",
    x"2E286662",
    x"2E285157",
    x"2E283C4E",
    x"2E282748",
    x"2E281244",
    x"2E27FD43",
    x"2E27E845",
    x"2E27D349",
    x"2E27BE50",
    x"2E27A95A",
    x"2E279466",
    x"2E277F75",
    x"2E276A86",
    x"2E27559A",
    x"2E2740B1",
    x"2E272BCA",
    x"2E2716E6",
    x"2E270204",
    x"2E26ED25",
    x"2E26D849",
    x"2E26C36F",
    x"2E26AE98",
    x"2E2699C3",
    x"2E2684F1",
    x"2E267022",
    x"2E265B55",
    x"2E26468B",
    x"2E2631C4",
    x"2E261CFF",
    x"2E26083C",
    x"2E25F37D",
    x"2E25DEC0",
    x"2E25CA05",
    x"2E25B54D",
    x"2E25A098",
    x"2E258BE5",
    x"2E257735",
    x"2E256287",
    x"2E254DDC",
    x"2E253934",
    x"2E25248E",
    x"2E250FEB",
    x"2E24FB4A",
    x"2E24E6AC",
    x"2E24D210",
    x"2E24BD77",
    x"2E24A8E1",
    x"2E24944D",
    x"2E247FBC",
    x"2E246B2D",
    x"2E2456A1",
    x"2E244217",
    x"2E242D90",
    x"2E24190C",
    x"2E24048A",
    x"2E23F00B",
    x"2E23DB8E",
    x"2E23C714",
    x"2E23B29C",
    x"2E239E27",
    x"2E2389B5",
    x"2E237545",
    x"2E2360D8",
    x"2E234C6D",
    x"2E233804",
    x"2E23239F",
    x"2E230F3C",
    x"2E22FADB",
    x"2E22E67D",
    x"2E22D221",
    x"2E22BDC8",
    x"2E22A972",
    x"2E22951E",
    x"2E2280CD",
    x"2E226C7E",
    x"2E225831",
    x"2E2243E8",
    x"2E222FA0",
    x"2E221B5C",
    x"2E22071A",
    x"2E21F2DA",
    x"2E21DE9D",
    x"2E21CA62",
    x"2E21B62A",
    x"2E21A1F5",
    x"2E218DC2",
    x"2E217991",
    x"2E216563",
    x"2E215138",
    x"2E213D0F",
    x"2E2128E9",
    x"2E2114C5",
    x"2E2100A4",
    x"2E20EC85",
    x"2E20D868",
    x"2E20C44F",
    x"2E20B037",
    x"2E209C23",
    x"2E208810",
    x"2E207401",
    x"2E205FF3",
    x"2E204BE9",
    x"2E2037E0",
    x"2E2023DB",
    x"2E200FD7",
    x"2E1FFBD7",
    x"2E1FE7D8",
    x"2E1FD3DD",
    x"2E1FBFE3",
    x"2E1FABED",
    x"2E1F97F8",
    x"2E1F8407",
    x"2E1F7017",
    x"2E1F5C2B",
    x"2E1F4840",
    x"2E1F3459",
    x"2E1F2073",
    x"2E1F0C91",
    x"2E1EF8B0",
    x"2E1EE4D2",
    x"2E1ED0F7",
    x"2E1EBD1E",
    x"2E1EA948",
    x"2E1E9574",
    x"2E1E81A2",
    x"2E1E6DD3",
    x"2E1E5A07",
    x"2E1E463D",
    x"2E1E3275",
    x"2E1E1EB0",
    x"2E1E0AEE",
    x"2E1DF72E",
    x"2E1DE370",
    x"2E1DCFB5",
    x"2E1DBBFC",
    x"2E1DA846",
    x"2E1D9492",
    x"2E1D80E1",
    x"2E1D6D32",
    x"2E1D5985",
    x"2E1D45DB",
    x"2E1D3234",
    x"2E1D1E8F",
    x"2E1D0AEC",
    x"2E1CF74C",
    x"2E1CE3AE",
    x"2E1CD013",
    x"2E1CBC7A",
    x"2E1CA8E4",
    x"2E1C9550",
    x"2E1C81BF",
    x"2E1C6E30",
    x"2E1C5AA3",
    x"2E1C4719",
    x"2E1C3391",
    x"2E1C200C",
    x"2E1C0C89",
    x"2E1BF909",
    x"2E1BE58B",
    x"2E1BD210",
    x"2E1BBE96",
    x"2E1BAB20",
    x"2E1B97AC",
    x"2E1B843A",
    x"2E1B70CB",
    x"2E1B5D5E",
    x"2E1B49F3",
    x"2E1B368B",
    x"2E1B2326",
    x"2E1B0FC2",
    x"2E1AFC62",
    x"2E1AE903",
    x"2E1AD5A7",
    x"2E1AC24E",
    x"2E1AAEF7",
    x"2E1A9BA2",
    x"2E1A8850",
    x"2E1A7500",
    x"2E1A61B3",
    x"2E1A4E68",
    x"2E1A3B1F",
    x"2E1A27D9",
    x"2E1A1495",
    x"2E1A0154",
    x"2E19EE15",
    x"2E19DAD8",
    x"2E19C79E",
    x"2E19B466",
    x"2E19A131",
    x"2E198DFE",
    x"2E197ACE",
    x"2E19679F",
    x"2E195474",
    x"2E19414A",
    x"2E192E23",
    x"2E191AFF",
    x"2E1907DD",
    x"2E18F4BD",
    x"2E18E19F",
    x"2E18CE84",
    x"2E18BB6C",
    x"2E18A856",
    x"2E189542",
    x"2E188230",
    x"2E186F21",
    x"2E185C14",
    x"2E18490A",
    x"2E183602",
    x"2E1822FD",
    x"2E180FF9",
    x"2E17FCF9",
    x"2E17E9FA",
    x"2E17D6FE",
    x"2E17C404",
    x"2E17B10D",
    x"2E179E18",
    x"2E178B26",
    x"2E177835",
    x"2E176548",
    x"2E17525C",
    x"2E173F73",
    x"2E172C8C",
    x"2E1719A8",
    x"2E1706C6",
    x"2E16F3E6",
    x"2E16E109",
    x"2E16CE2E",
    x"2E16BB55",
    x"2E16A87F",
    x"2E1695AB",
    x"2E1682DA",
    x"2E16700A",
    x"2E165D3E",
    x"2E164A73",
    x"2E1637AB",
    x"2E1624E5",
    x"2E161222",
    x"2E15FF61",
    x"2E15ECA2",
    x"2E15D9E5",
    x"2E15C72B",
    x"2E15B474",
    x"2E15A1BE",
    x"2E158F0B",
    x"2E157C5B",
    x"2E1569AC",
    x"2E155700",
    x"2E154456",
    x"2E1531AF",
    x"2E151F0A",
    x"2E150C67",
    x"2E14F9C7",
    x"2E14E729",
    x"2E14D48D",
    x"2E14C1F4",
    x"2E14AF5D",
    x"2E149CC8",
    x"2E148A35",
    x"2E1477A5",
    x"2E146518",
    x"2E14528C",
    x"2E144003",
    x"2E142D7C",
    x"2E141AF8",
    x"2E140875",
    x"2E13F5F5",
    x"2E13E378",
    x"2E13D0FD",
    x"2E13BE84",
    x"2E13AC0D",
    x"2E139999",
    x"2E138726",
    x"2E1374B7",
    x"2E136249",
    x"2E134FDE",
    x"2E133D75",
    x"2E132B0F",
    x"2E1318AB",
    x"2E130649",
    x"2E12F3E9",
    x"2E12E18C",
    x"2E12CF31",
    x"2E12BCD8",
    x"2E12AA81",
    x"2E12982D",
    x"2E1285DB",
    x"2E12738C",
    x"2E12613E",
    x"2E124EF3",
    x"2E123CAB",
    x"2E122A64",
    x"2E121820",
    x"2E1205DE",
    x"2E11F39F",
    x"2E11E161",
    x"2E11CF26",
    x"2E11BCEE",
    x"2E11AAB7",
    x"2E119883",
    x"2E118651",
    x"2E117421",
    x"2E1161F4",
    x"2E114FC9",
    x"2E113DA0",
    x"2E112B79",
    x"2E111955",
    x"2E110733",
    x"2E10F513",
    x"2E10E2F6",
    x"2E10D0DB",
    x"2E10BEC2",
    x"2E10ACAB",
    x"2E109A96",
    x"2E108884",
    x"2E107674",
    x"2E106467",
    x"2E10525B",
    x"2E104052",
    x"2E102E4B",
    x"2E101C46",
    x"2E100A44",
    x"2E0FF844",
    x"2E0FE646",
    x"2E0FD44A",
    x"2E0FC251",
    x"2E0FB05A",
    x"2E0F9E65",
    x"2E0F8C72",
    x"2E0F7A82",
    x"2E0F6894",
    x"2E0F56A8",
    x"2E0F44BE",
    x"2E0F32D6",
    x"2E0F20F1",
    x"2E0F0F0E",
    x"2E0EFD2D",
    x"2E0EEB4F",
    x"2E0ED973",
    x"2E0EC798",
    x"2E0EB5C1",
    x"2E0EA3EB",
    x"2E0E9218",
    x"2E0E8047",
    x"2E0E6E78",
    x"2E0E5CAB",
    x"2E0E4AE0",
    x"2E0E3918",
    x"2E0E2752",
    x"2E0E158E",
    x"2E0E03CD",
    x"2E0DF20D",
    x"2E0DE050",
    x"2E0DCE95",
    x"2E0DBCDD",
    x"2E0DAB26",
    x"2E0D9972",
    x"2E0D87C0",
    x"2E0D7610",
    x"2E0D6462",
    x"2E0D52B7",
    x"2E0D410E",
    x"2E0D2F67",
    x"2E0D1DC2",
    x"2E0D0C1F",
    x"2E0CFA7F",
    x"2E0CE8E0",
    x"2E0CD744",
    x"2E0CC5AB",
    x"2E0CB413",
    x"2E0CA27E",
    x"2E0C90EA",
    x"2E0C7F59",
    x"2E0C6DCB",
    x"2E0C5C3E",
    x"2E0C4AB4",
    x"2E0C392B",
    x"2E0C27A5",
    x"2E0C1621",
    x"2E0C04A0",
    x"2E0BF320",
    x"2E0BE1A3",
    x"2E0BD028",
    x"2E0BBEAF",
    x"2E0BAD38",
    x"2E0B9BC4",
    x"2E0B8A51",
    x"2E0B78E1",
    x"2E0B6773",
    x"2E0B5607",
    x"2E0B449D",
    x"2E0B3336",
    x"2E0B21D1",
    x"2E0B106E",
    x"2E0AFF0D",
    x"2E0AEDAE",
    x"2E0ADC51",
    x"2E0ACAF7",
    x"2E0AB99E",
    x"2E0AA848",
    x"2E0A96F4",
    x"2E0A85A3",
    x"2E0A7453",
    x"2E0A6305",
    x"2E0A51BA",
    x"2E0A4071",
    x"2E0A2F2A",
    x"2E0A1DE5",
    x"2E0A0CA3",
    x"2E09FB62",
    x"2E09EA24",
    x"2E09D8E8",
    x"2E09C7AE",
    x"2E09B676",
    x"2E09A540",
    x"2E09940C",
    x"2E0982DB",
    x"2E0971AC",
    x"2E09607E",
    x"2E094F53",
    x"2E093E2B",
    x"2E092D04",
    x"2E091BDF",
    x"2E090ABD",
    x"2E08F99D",
    x"2E08E87F",
    x"2E08D763",
    x"2E08C649",
    x"2E08B531",
    x"2E08A41B",
    x"2E089308",
    x"2E0881F7",
    x"2E0870E7",
    x"2E085FDA",
    x"2E084ED0",
    x"2E083DC7",
    x"2E082CC0",
    x"2E081BBC",
    x"2E080AB9",
    x"2E07F9B9",
    x"2E07E8BB",
    x"2E07D7BF",
    x"2E07C6C5",
    x"2E07B5CD",
    x"2E07A4D7",
    x"2E0793E4",
    x"2E0782F2",
    x"2E077203",
    x"2E076116",
    x"2E07502B",
    x"2E073F42",
    x"2E072E5B",
    x"2E071D76",
    x"2E070C94",
    x"2E06FBB3",
    x"2E06EAD5",
    x"2E06D9F8",
    x"2E06C91E",
    x"2E06B846",
    x"2E06A770",
    x"2E06969C",
    x"2E0685CA",
    x"2E0674FB",
    x"2E06642D",
    x"2E065362",
    x"2E064298",
    x"2E0631D1",
    x"2E06210C",
    x"2E061049",
    x"2E05FF88",
    x"2E05EEC9",
    x"2E05DE0C",
    x"2E05CD51",
    x"2E05BC99",
    x"2E05ABE2",
    x"2E059B2E",
    x"2E058A7B",
    x"2E0579CB",
    x"2E05691D",
    x"2E055871",
    x"2E0547C7",
    x"2E05371F",
    x"2E052679",
    x"2E0515D5",
    x"2E050534",
    x"2E04F494",
    x"2E04E3F7",
    x"2E04D35B",
    x"2E04C2C2",
    x"2E04B22A",
    x"2E04A195",
    x"2E049102",
    x"2E048071",
    x"2E046FE2",
    x"2E045F55",
    x"2E044ECA",
    x"2E043E41",
    x"2E042DBA",
    x"2E041D36",
    x"2E040CB3",
    x"2E03FC33",
    x"2E03EBB4",
    x"2E03DB38",
    x"2E03CABD",
    x"2E03BA45",
    x"2E03A9CF",
    x"2E03995B",
    x"2E0388E8",
    x"2E037878",
    x"2E03680A",
    x"2E03579E",
    x"2E034734",
    x"2E0336CD",
    x"2E032667",
    x"2E031603",
    x"2E0305A1",
    x"2E02F542",
    x"2E02E4E4",
    x"2E02D488",
    x"2E02C42F",
    x"2E02B3D7",
    x"2E02A382",
    x"2E02932E",
    x"2E0282DD",
    x"2E02728E",
    x"2E026240",
    x"2E0251F5",
    x"2E0241AC",
    x"2E023165",
    x"2E022120",
    x"2E0210DC",
    x"2E02009B",
    x"2E01F05C",
    x"2E01E01F",
    x"2E01CFE4",
    x"2E01BFAB",
    x"2E01AF74",
    x"2E019F3F",
    x"2E018F0C",
    x"2E017EDC",
    x"2E016EAD",
    x"2E015E80",
    x"2E014E55",
    x"2E013E2C",
    x"2E012E06",
    x"2E011DE1",
    x"2E010DBE",
    x"2E00FD9D",
    x"2E00ED7F",
    x"2E00DD62",
    x"2E00CD47",
    x"2E00BD2F",
    x"2E00AD18",
    x"2E009D03",
    x"2E008CF1",
    x"2E007CE0",
    x"2E006CD2",
    x"2E005CC5",
    x"2E004CBA",
    x"2E003CB2",
    x"2E002CAB",
    x"2E001CA7",
    x"2E000CA4",
    x"2DFFF947",
    x"2DFFD94A",
    x"2DFFB951",
    x"2DFF995B",
    x"2DFF796A",
    x"2DFF597D",
    x"2DFF3994",
    x"2DFF19AF",
    x"2DFEF9CE",
    x"2DFED9F0",
    x"2DFEBA17",
    x"2DFE9A42",
    x"2DFE7A70",
    x"2DFE5AA3",
    x"2DFE3ADA",
    x"2DFE1B14",
    x"2DFDFB53",
    x"2DFDDB96",
    x"2DFDBBDC",
    x"2DFD9C27",
    x"2DFD7C75",
    x"2DFD5CC8",
    x"2DFD3D1E",
    x"2DFD1D78",
    x"2DFCFDD7",
    x"2DFCDE39",
    x"2DFCBE9F",
    x"2DFC9F09",
    x"2DFC7F77",
    x"2DFC5FE9",
    x"2DFC405F",
    x"2DFC20D9",
    x"2DFC0157",
    x"2DFBE1D9",
    x"2DFBC25F",
    x"2DFBA2E8",
    x"2DFB8376",
    x"2DFB6407",
    x"2DFB449D",
    x"2DFB2536",
    x"2DFB05D4",
    x"2DFAE675",
    x"2DFAC71A",
    x"2DFAA7C3",
    x"2DFA8870",
    x"2DFA6921",
    x"2DFA49D6",
    x"2DFA2A8E",
    x"2DFA0B4B",
    x"2DF9EC0C",
    x"2DF9CCD0",
    x"2DF9AD98",
    x"2DF98E65",
    x"2DF96F35",
    x"2DF95009",
    x"2DF930E1",
    x"2DF911BD",
    x"2DF8F29C",
    x"2DF8D380",
    x"2DF8B467",
    x"2DF89553",
    x"2DF87642",
    x"2DF85735",
    x"2DF8382C",
    x"2DF81927",
    x"2DF7FA26",
    x"2DF7DB29",
    x"2DF7BC2F",
    x"2DF79D3A",
    x"2DF77E48",
    x"2DF75F5A",
    x"2DF74070",
    x"2DF7218A",
    x"2DF702A8",
    x"2DF6E3C9",
    x"2DF6C4EF",
    x"2DF6A618",
    x"2DF68745",
    x"2DF66876",
    x"2DF649AB",
    x"2DF62AE4",
    x"2DF60C20",
    x"2DF5ED61",
    x"2DF5CEA5",
    x"2DF5AFED",
    x"2DF59139",
    x"2DF57289",
    x"2DF553DC",
    x"2DF53534",
    x"2DF5168F",
    x"2DF4F7EE",
    x"2DF4D951",
    x"2DF4BAB8",
    x"2DF49C22",
    x"2DF47D91",
    x"2DF45F03",
    x"2DF44079",
    x"2DF421F3",
    x"2DF40371",
    x"2DF3E4F2",
    x"2DF3C677",
    x"2DF3A800",
    x"2DF3898D",
    x"2DF36B1E",
    x"2DF34CB3",
    x"2DF32E4B",
    x"2DF30FE7",
    x"2DF2F187",
    x"2DF2D32B",
    x"2DF2B4D2",
    x"2DF2967D",
    x"2DF2782D",
    x"2DF259DF",
    x"2DF23B96",
    x"2DF21D51",
    x"2DF1FF0F",
    x"2DF1E0D1",
    x"2DF1C297",
    x"2DF1A460",
    x"2DF1862D",
    x"2DF167FF",
    x"2DF149D3",
    x"2DF12BAC",
    x"2DF10D89",
    x"2DF0EF69",
    x"2DF0D14D",
    x"2DF0B334",
    x"2DF09520",
    x"2DF0770F",
    x"2DF05902",
    x"2DF03AF9",
    x"2DF01CF3",
    x"2DEFFEF2",
    x"2DEFE0F4",
    x"2DEFC2F9",
    x"2DEFA503",
    x"2DEF8710",
    x"2DEF6921",
    x"2DEF4B36",
    x"2DEF2D4E",
    x"2DEF0F6B",
    x"2DEEF18A",
    x"2DEED3AE",
    x"2DEEB5D6",
    x"2DEE9801",
    x"2DEE7A30",
    x"2DEE5C62",
    x"2DEE3E98",
    x"2DEE20D2",
    x"2DEE0310",
    x"2DEDE552",
    x"2DEDC797",
    x"2DEDA9E0",
    x"2DED8C2C",
    x"2DED6E7D",
    x"2DED50D1",
    x"2DED3329",
    x"2DED1584",
    x"2DECF7E3",
    x"2DECDA46",
    x"2DECBCAD",
    x"2DEC9F17",
    x"2DEC8185",
    x"2DEC63F6",
    x"2DEC466C",
    x"2DEC28E5",
    x"2DEC0B62",
    x"2DEBEDE2",
    x"2DEBD066",
    x"2DEBB2EE",
    x"2DEB9579",
    x"2DEB7809",
    x"2DEB5A9B",
    x"2DEB3D32",
    x"2DEB1FCC",
    x"2DEB026A",
    x"2DEAE50C",
    x"2DEAC7B1",
    x"2DEAAA5A",
    x"2DEA8D06",
    x"2DEA6FB6",
    x"2DEA526A",
    x"2DEA3522",
    x"2DEA17DD",
    x"2DE9FA9C",
    x"2DE9DD5E",
    x"2DE9C024",
    x"2DE9A2EE",
    x"2DE985BC",
    x"2DE9688D",
    x"2DE94B62",
    x"2DE92E3A",
    x"2DE91116",
    x"2DE8F3F6",
    x"2DE8D6D9",
    x"2DE8B9C0",
    x"2DE89CAB",
    x"2DE87F99",
    x"2DE8628B",
    x"2DE84580",
    x"2DE82879",
    x"2DE80B76",
    x"2DE7EE76",
    x"2DE7D17A",
    x"2DE7B482",
    x"2DE7978D",
    x"2DE77A9C",
    x"2DE75DAF",
    x"2DE740C5",
    x"2DE723DE",
    x"2DE706FC",
    x"2DE6EA1D",
    x"2DE6CD41",
    x"2DE6B069",
    x"2DE69395",
    x"2DE676C4",
    x"2DE659F7",
    x"2DE63D2E",
    x"2DE62068",
    x"2DE603A6",
    x"2DE5E6E7",
    x"2DE5CA2C",
    x"2DE5AD75",
    x"2DE590C1",
    x"2DE57411",
    x"2DE55764",
    x"2DE53ABB",
    x"2DE51E15",
    x"2DE50173",
    x"2DE4E4D5",
    x"2DE4C83A",
    x"2DE4ABA3",
    x"2DE48F0F",
    x"2DE4727F",
    x"2DE455F2",
    x"2DE43969",
    x"2DE41CE4",
    x"2DE40062",
    x"2DE3E3E4",
    x"2DE3C769",
    x"2DE3AAF2",
    x"2DE38E7E",
    x"2DE3720E",
    x"2DE355A2",
    x"2DE33939",
    x"2DE31CD4",
    x"2DE30072",
    x"2DE2E414",
    x"2DE2C7B9",
    x"2DE2AB62",
    x"2DE28F0E",
    x"2DE272BE",
    x"2DE25671",
    x"2DE23A28",
    x"2DE21DE3",
    x"2DE201A1",
    x"2DE1E562",
    x"2DE1C927",
    x"2DE1ACF0",
    x"2DE190BC",
    x"2DE1748C",
    x"2DE1585F",
    x"2DE13C36",
    x"2DE12010",
    x"2DE103EE",
    x"2DE0E7CF",
    x"2DE0CBB4",
    x"2DE0AF9C",
    x"2DE09388",
    x"2DE07777",
    x"2DE05B6A",
    x"2DE03F60",
    x"2DE0235A",
    x"2DE00758",
    x"2DDFEB58",
    x"2DDFCF5D",
    x"2DDFB365",
    x"2DDF9770",
    x"2DDF7B7F",
    x"2DDF5F91",
    x"2DDF43A7",
    x"2DDF27C0",
    x"2DDF0BDD",
    x"2DDEEFFD",
    x"2DDED421",
    x"2DDEB848",
    x"2DDE9C73",
    x"2DDE80A1",
    x"2DDE64D3",
    x"2DDE4908",
    x"2DDE2D40",
    x"2DDE117C",
    x"2DDDF5BC",
    x"2DDDD9FF",
    x"2DDDBE45",
    x"2DDDA28F",
    x"2DDD86DD",
    x"2DDD6B2E",
    x"2DDD4F82",
    x"2DDD33DA",
    x"2DDD1835",
    x"2DDCFC94",
    x"2DDCE0F6",
    x"2DDCC55C",
    x"2DDCA9C5",
    x"2DDC8E31",
    x"2DDC72A1",
    x"2DDC5714",
    x"2DDC3B8B",
    x"2DDC2006",
    x"2DDC0483",
    x"2DDBE904",
    x"2DDBCD89",
    x"2DDBB211",
    x"2DDB969C",
    x"2DDB7B2B",
    x"2DDB5FBE",
    x"2DDB4453",
    x"2DDB28ED",
    x"2DDB0D89",
    x"2DDAF229",
    x"2DDAD6CD",
    x"2DDABB74",
    x"2DDAA01E",
    x"2DDA84CC",
    x"2DDA697D",
    x"2DDA4E31",
    x"2DDA32E9",
    x"2DDA17A4",
    x"2DD9FC63",
    x"2DD9E125",
    x"2DD9C5EB",
    x"2DD9AAB4",
    x"2DD98F80",
    x"2DD97450",
    x"2DD95923",
    x"2DD93DFA",
    x"2DD922D4",
    x"2DD907B1",
    x"2DD8EC92",
    x"2DD8D176",
    x"2DD8B65D",
    x"2DD89B48",
    x"2DD88037",
    x"2DD86528",
    x"2DD84A1D",
    x"2DD82F16",
    x"2DD81411",
    x"2DD7F911",
    x"2DD7DE13",
    x"2DD7C319",
    x"2DD7A822",
    x"2DD78D2F",
    x"2DD7723F",
    x"2DD75753",
    x"2DD73C69",
    x"2DD72183",
    x"2DD706A1",
    x"2DD6EBC2",
    x"2DD6D0E6",
    x"2DD6B60E",
    x"2DD69B38",
    x"2DD68067",
    x"2DD66598",
    x"2DD64ACD",
    x"2DD63006",
    x"2DD61541",
    x"2DD5FA80",
    x"2DD5DFC3",
    x"2DD5C508",
    x"2DD5AA51",
    x"2DD58F9E",
    x"2DD574EE",
    x"2DD55A41",
    x"2DD53F97",
    x"2DD524F1",
    x"2DD50A4E",
    x"2DD4EFAE",
    x"2DD4D512",
    x"2DD4BA79",
    x"2DD49FE3",
    x"2DD48551",
    x"2DD46AC2",
    x"2DD45036",
    x"2DD435AE",
    x"2DD41B29",
    x"2DD400A7",
    x"2DD3E629",
    x"2DD3CBAD",
    x"2DD3B136",
    x"2DD396C1",
    x"2DD37C50",
    x"2DD361E2",
    x"2DD34778",
    x"2DD32D10",
    x"2DD312AC",
    x"2DD2F84C",
    x"2DD2DDEE",
    x"2DD2C394",
    x"2DD2A93D",
    x"2DD28EEA",
    x"2DD2749A",
    x"2DD25A4D",
    x"2DD24003",
    x"2DD225BD",
    x"2DD20B7A",
    x"2DD1F13A",
    x"2DD1D6FD",
    x"2DD1BCC4",
    x"2DD1A28E",
    x"2DD1885B",
    x"2DD16E2C",
    x"2DD15400",
    x"2DD139D7",
    x"2DD11FB1",
    x"2DD1058F",
    x"2DD0EB70",
    x"2DD0D154",
    x"2DD0B73C",
    x"2DD09D26",
    x"2DD08314",
    x"2DD06906",
    x"2DD04EFA",
    x"2DD034F2",
    x"2DD01AED",
    x"2DD000EB",
    x"2DCFE6ED",
    x"2DCFCCF1",
    x"2DCFB2F9",
    x"2DCF9905",
    x"2DCF7F13",
    x"2DCF6525",
    x"2DCF4B3A",
    x"2DCF3152",
    x"2DCF176E",
    x"2DCEFD8C",
    x"2DCEE3AE",
    x"2DCEC9D3",
    x"2DCEAFFC",
    x"2DCE9627",
    x"2DCE7C56",
    x"2DCE6288",
    x"2DCE48BD",
    x"2DCE2EF6",
    x"2DCE1532",
    x"2DCDFB71",
    x"2DCDE1B3",
    x"2DCDC7F8",
    x"2DCDAE41",
    x"2DCD948D",
    x"2DCD7ADC",
    x"2DCD612E",
    x"2DCD4783",
    x"2DCD2DDC",
    x"2DCD1438",
    x"2DCCFA97",
    x"2DCCE0F9",
    x"2DCCC75F",
    x"2DCCADC8",
    x"2DCC9433",
    x"2DCC7AA2",
    x"2DCC6115",
    x"2DCC478A",
    x"2DCC2E03",
    x"2DCC147F",
    x"2DCBFAFE",
    x"2DCBE180",
    x"2DCBC805",
    x"2DCBAE8E",
    x"2DCB951A",
    x"2DCB7BA9",
    x"2DCB623B",
    x"2DCB48D0",
    x"2DCB2F69",
    x"2DCB1604",
    x"2DCAFCA3",
    x"2DCAE345",
    x"2DCAC9EA",
    x"2DCAB093",
    x"2DCA973E",
    x"2DCA7DED",
    x"2DCA649F",
    x"2DCA4B54",
    x"2DCA320C",
    x"2DCA18C7",
    x"2DC9FF86",
    x"2DC9E647",
    x"2DC9CD0C",
    x"2DC9B3D4",
    x"2DC99A9F",
    x"2DC9816D",
    x"2DC9683F",
    x"2DC94F13",
    x"2DC935EB",
    x"2DC91CC6",
    x"2DC903A4",
    x"2DC8EA85",
    x"2DC8D169",
    x"2DC8B851",
    x"2DC89F3B",
    x"2DC88629",
    x"2DC86D1A",
    x"2DC8540D",
    x"2DC83B04",
    x"2DC821FF",
    x"2DC808FC",
    x"2DC7EFFC",
    x"2DC7D700",
    x"2DC7BE07",
    x"2DC7A510",
    x"2DC78C1D",
    x"2DC7732D",
    x"2DC75A41",
    x"2DC74157",
    x"2DC72870",
    x"2DC70F8D",
    x"2DC6F6AC",
    x"2DC6DDCF",
    x"2DC6C4F5",
    x"2DC6AC1E",
    x"2DC6934A",
    x"2DC67A79",
    x"2DC661AB",
    x"2DC648E1",
    x"2DC63019",
    x"2DC61755",
    x"2DC5FE93",
    x"2DC5E5D5",
    x"2DC5CD1A",
    x"2DC5B462",
    x"2DC59BAD",
    x"2DC582FB",
    x"2DC56A4C",
    x"2DC551A0",
    x"2DC538F8",
    x"2DC52052",
    x"2DC507AF",
    x"2DC4EF10",
    x"2DC4D674",
    x"2DC4BDDA",
    x"2DC4A544",
    x"2DC48CB1",
    x"2DC47421",
    x"2DC45B94",
    x"2DC4430A",
    x"2DC42A83",
    x"2DC41200",
    x"2DC3F97F",
    x"2DC3E101",
    x"2DC3C887",
    x"2DC3B00F",
    x"2DC3979B",
    x"2DC37F29",
    x"2DC366BB",
    x"2DC34E4F",
    x"2DC335E7",
    x"2DC31D82",
    x"2DC30520",
    x"2DC2ECC1",
    x"2DC2D465",
    x"2DC2BC0C",
    x"2DC2A3B6",
    x"2DC28B63",
    x"2DC27313",
    x"2DC25AC6",
    x"2DC2427C",
    x"2DC22A35",
    x"2DC211F2",
    x"2DC1F9B1",
    x"2DC1E173",
    x"2DC1C938",
    x"2DC1B101",
    x"2DC198CC",
    x"2DC1809B",
    x"2DC1686C",
    x"2DC15040",
    x"2DC13818",
    x"2DC11FF2",
    x"2DC107D0",
    x"2DC0EFB0",
    x"2DC0D794",
    x"2DC0BF7B",
    x"2DC0A764",
    x"2DC08F51",
    x"2DC07740",
    x"2DC05F33",
    x"2DC04729",
    x"2DC02F21",
    x"2DC0171D",
    x"2DBFFF1B",
    x"2DBFE71D",
    x"2DBFCF22",
    x"2DBFB729",
    x"2DBF9F34",
    x"2DBF8741",
    x"2DBF6F52",
    x"2DBF5766",
    x"2DBF3F7C",
    x"2DBF2796",
    x"2DBF0FB2",
    x"2DBEF7D2",
    x"2DBEDFF4",
    x"2DBEC81A",
    x"2DBEB042",
    x"2DBE986E",
    x"2DBE809C",
    x"2DBE68CE",
    x"2DBE5102",
    x"2DBE3939",
    x"2DBE2174",
    x"2DBE09B1",
    x"2DBDF1F1",
    x"2DBDDA34",
    x"2DBDC27B",
    x"2DBDAAC4",
    x"2DBD9310",
    x"2DBD7B5F",
    x"2DBD63B1",
    x"2DBD4C06",
    x"2DBD345E",
    x"2DBD1CB9",
    x"2DBD0517",
    x"2DBCED78",
    x"2DBCD5DC",
    x"2DBCBE42",
    x"2DBCA6AC",
    x"2DBC8F19",
    x"2DBC7788",
    x"2DBC5FFB",
    x"2DBC4870",
    x"2DBC30E9",
    x"2DBC1964",
    x"2DBC01E2",
    x"2DBBEA64",
    x"2DBBD2E8",
    x"2DBBBB6F",
    x"2DBBA3F9",
    x"2DBB8C86",
    x"2DBB7516",
    x"2DBB5DA9",
    x"2DBB463E",
    x"2DBB2ED7",
    x"2DBB1773",
    x"2DBB0011",
    x"2DBAE8B3",
    x"2DBAD157",
    x"2DBAB9FE",
    x"2DBAA2A8",
    x"2DBA8B56",
    x"2DBA7406",
    x"2DBA5CB9",
    x"2DBA456E",
    x"2DBA2E27",
    x"2DBA16E3",
    x"2DB9FFA1",
    x"2DB9E863",
    x"2DB9D127",
    x"2DB9B9EF",
    x"2DB9A2B9",
    x"2DB98B86",
    x"2DB97456",
    x"2DB95D29",
    x"2DB945FF",
    x"2DB92ED7",
    x"2DB917B3",
    x"2DB90092",
    x"2DB8E973",
    x"2DB8D257",
    x"2DB8BB3E",
    x"2DB8A428",
    x"2DB88D15",
    x"2DB87605",
    x"2DB85EF8",
    x"2DB847ED",
    x"2DB830E6",
    x"2DB819E1",
    x"2DB802DF",
    x"2DB7EBE0",
    x"2DB7D4E4",
    x"2DB7BDEB",
    x"2DB7A6F5",
    x"2DB79001",
    x"2DB77911",
    x"2DB76223",
    x"2DB74B38",
    x"2DB73450",
    x"2DB71D6B",
    x"2DB70689",
    x"2DB6EFAA",
    x"2DB6D8CD",
    x"2DB6C1F3",
    x"2DB6AB1D",
    x"2DB69449",
    x"2DB67D78",
    x"2DB666A9",
    x"2DB64FDE",
    x"2DB63915",
    x"2DB62250",
    x"2DB60B8D",
    x"2DB5F4CD",
    x"2DB5DE10",
    x"2DB5C755",
    x"2DB5B09E",
    x"2DB599E9",
    x"2DB58337",
    x"2DB56C88",
    x"2DB555DC",
    x"2DB53F33",
    x"2DB5288C",
    x"2DB511E9",
    x"2DB4FB48",
    x"2DB4E4AA",
    x"2DB4CE0F",
    x"2DB4B776",
    x"2DB4A0E1",
    x"2DB48A4E",
    x"2DB473BE",
    x"2DB45D31",
    x"2DB446A7",
    x"2DB4301F",
    x"2DB4199B",
    x"2DB40319",
    x"2DB3EC9A",
    x"2DB3D61E",
    x"2DB3BFA5",
    x"2DB3A92E",
    x"2DB392BA",
    x"2DB37C49",
    x"2DB365DB",
    x"2DB34F70",
    x"2DB33907",
    x"2DB322A2",
    x"2DB30C3F",
    x"2DB2F5DF",
    x"2DB2DF81",
    x"2DB2C927",
    x"2DB2B2CF",
    x"2DB29C7A",
    x"2DB28628",
    x"2DB26FD8",
    x"2DB2598C",
    x"2DB24342",
    x"2DB22CFB",
    x"2DB216B7",
    x"2DB20075",
    x"2DB1EA37",
    x"2DB1D3FB",
    x"2DB1BDC2",
    x"2DB1A78B",
    x"2DB19158",
    x"2DB17B27",
    x"2DB164F9",
    x"2DB14ECE",
    x"2DB138A5",
    x"2DB12280",
    x"2DB10C5D",
    x"2DB0F63C",
    x"2DB0E01F",
    x"2DB0CA04",
    x"2DB0B3ED",
    x"2DB09DD7",
    x"2DB087C5",
    x"2DB071B6",
    x"2DB05BA9",
    x"2DB0459F",
    x"2DB02F97",
    x"2DB01993",
    x"2DB00391",
    x"2DAFED92",
    x"2DAFD796",
    x"2DAFC19C",
    x"2DAFABA5",
    x"2DAF95B1",
    x"2DAF7FC0",
    x"2DAF69D1",
    x"2DAF53E5",
    x"2DAF3DFC",
    x"2DAF2816",
    x"2DAF1232",
    x"2DAEFC51",
    x"2DAEE673",
    x"2DAED098",
    x"2DAEBABF",
    x"2DAEA4E9",
    x"2DAE8F16",
    x"2DAE7945",
    x"2DAE6377",
    x"2DAE4DAC",
    x"2DAE37E4",
    x"2DAE221E",
    x"2DAE0C5B",
    x"2DADF69B",
    x"2DADE0DE",
    x"2DADCB23",
    x"2DADB56B",
    x"2DAD9FB6",
    x"2DAD8A03",
    x"2DAD7453",
    x"2DAD5EA6",
    x"2DAD48FB",
    x"2DAD3354",
    x"2DAD1DAF",
    x"2DAD080C",
    x"2DACF26D",
    x"2DACDCD0",
    x"2DACC735",
    x"2DACB19E",
    x"2DAC9C09",
    x"2DAC8677",
    x"2DAC70E7",
    x"2DAC5B5B",
    x"2DAC45D1",
    x"2DAC3049",
    x"2DAC1AC4",
    x"2DAC0542",
    x"2DABEFC3",
    x"2DABDA47",
    x"2DABC4CD",
    x"2DABAF55",
    x"2DAB99E1",
    x"2DAB846F",
    x"2DAB6F00",
    x"2DAB5993",
    x"2DAB4429",
    x"2DAB2EC2",
    x"2DAB195E",
    x"2DAB03FC",
    x"2DAAEE9D",
    x"2DAAD940",
    x"2DAAC3E6",
    x"2DAAAE8F",
    x"2DAA993B",
    x"2DAA83E9",
    x"2DAA6E9A",
    x"2DAA594D",
    x"2DAA4403",
    x"2DAA2EBC",
    x"2DAA1978",
    x"2DAA0436",
    x"2DA9EEF7",
    x"2DA9D9BA",
    x"2DA9C480",
    x"2DA9AF49",
    x"2DA99A14",
    x"2DA984E2",
    x"2DA96FB3",
    x"2DA95A86",
    x"2DA9455C",
    x"2DA93035",
    x"2DA91B10",
    x"2DA905EE",
    x"2DA8F0CF",
    x"2DA8DBB2",
    x"2DA8C698",
    x"2DA8B180",
    x"2DA89C6C",
    x"2DA88759",
    x"2DA8724A",
    x"2DA85D3D",
    x"2DA84832",
    x"2DA8332B",
    x"2DA81E26",
    x"2DA80923",
    x"2DA7F423",
    x"2DA7DF26",
    x"2DA7CA2C",
    x"2DA7B534",
    x"2DA7A03E",
    x"2DA78B4C",
    x"2DA7765B",
    x"2DA7616E",
    x"2DA74C83",
    x"2DA7379B",
    x"2DA722B5",
    x"2DA70DD2",
    x"2DA6F8F2",
    x"2DA6E414",
    x"2DA6CF39",
    x"2DA6BA60",
    x"2DA6A58A",
    x"2DA690B7",
    x"2DA67BE6",
    x"2DA66718",
    x"2DA6524C",
    x"2DA63D83",
    x"2DA628BD",
    x"2DA613F9",
    x"2DA5FF38",
    x"2DA5EA79",
    x"2DA5D5BD",
    x"2DA5C104",
    x"2DA5AC4D",
    x"2DA59799",
    x"2DA582E7",
    x"2DA56E38",
    x"2DA5598C",
    x"2DA544E2",
    x"2DA5303A",
    x"2DA51B96",
    x"2DA506F3",
    x"2DA4F254",
    x"2DA4DDB7",
    x"2DA4C91C",
    x"2DA4B485",
    x"2DA49FEF",
    x"2DA48B5D",
    x"2DA476CC",
    x"2DA4623F",
    x"2DA44DB4",
    x"2DA4392B",
    x"2DA424A6",
    x"2DA41022",
    x"2DA3FBA2",
    x"2DA3E723",
    x"2DA3D2A8",
    x"2DA3BE2F",
    x"2DA3A9B8",
    x"2DA39544",
    x"2DA380D3",
    x"2DA36C64",
    x"2DA357F8",
    x"2DA3438E",
    x"2DA32F27",
    x"2DA31AC2",
    x"2DA30660",
    x"2DA2F201",
    x"2DA2DDA4",
    x"2DA2C949",
    x"2DA2B4F1",
    x"2DA2A09C",
    x"2DA28C49",
    x"2DA277F9",
    x"2DA263AB",
    x"2DA24F60",
    x"2DA23B17",
    x"2DA226D1",
    x"2DA2128E",
    x"2DA1FE4D",
    x"2DA1EA0E",
    x"2DA1D5D2",
    x"2DA1C199",
    x"2DA1AD62",
    x"2DA1992D",
    x"2DA184FB",
    x"2DA170CC",
    x"2DA15C9F",
    x"2DA14875",
    x"2DA1344D",
    x"2DA12028",
    x"2DA10C05",
    x"2DA0F7E5",
    x"2DA0E3C7",
    x"2DA0CFAC",
    x"2DA0BB93",
    x"2DA0A77D",
    x"2DA09369",
    x"2DA07F58",
    x"2DA06B49",
    x"2DA0573D",
    x"2DA04334",
    x"2DA02F2D",
    x"2DA01B28",
    x"2DA00726",
    x"2D9FF326",
    x"2D9FDF29",
    x"2D9FCB2E",
    x"2D9FB736",
    x"2D9FA340",
    x"2D9F8F4D",
    x"2D9F7B5D",
    x"2D9F676E",
    x"2D9F5383",
    x"2D9F3F9A",
    x"2D9F2BB3",
    x"2D9F17CF",
    x"2D9F03ED",
    x"2D9EF00E",
    x"2D9EDC31",
    x"2D9EC857",
    x"2D9EB47F",
    x"2D9EA0AA",
    x"2D9E8CD7",
    x"2D9E7906",
    x"2D9E6538",
    x"2D9E516D",
    x"2D9E3DA4",
    x"2D9E29DE",
    x"2D9E161A",
    x"2D9E0258",
    x"2D9DEE99",
    x"2D9DDADC",
    x"2D9DC722",
    x"2D9DB36B",
    x"2D9D9FB5",
    x"2D9D8C03",
    x"2D9D7852",
    x"2D9D64A5",
    x"2D9D50F9",
    x"2D9D3D50",
    x"2D9D29AA",
    x"2D9D1606",
    x"2D9D0264",
    x"2D9CEEC5",
    x"2D9CDB29",
    x"2D9CC78F",
    x"2D9CB3F7",
    x"2D9CA062",
    x"2D9C8CCF",
    x"2D9C793E",
    x"2D9C65B0",
    x"2D9C5225",
    x"2D9C3E9C",
    x"2D9C2B15",
    x"2D9C1791",
    x"2D9C040F",
    x"2D9BF090",
    x"2D9BDD13",
    x"2D9BC999",
    x"2D9BB621",
    x"2D9BA2AB",
    x"2D9B8F38",
    x"2D9B7BC8",
    x"2D9B6859",
    x"2D9B54ED",
    x"2D9B4184",
    x"2D9B2E1D",
    x"2D9B1AB9",
    x"2D9B0756",
    x"2D9AF3F7",
    x"2D9AE099",
    x"2D9ACD3F",
    x"2D9AB9E6",
    x"2D9AA690",
    x"2D9A933C",
    x"2D9A7FEB",
    x"2D9A6C9C",
    x"2D9A5950",
    x"2D9A4606",
    x"2D9A32BF",
    x"2D9A1F79",
    x"2D9A0C37",
    x"2D99F8F6",
    x"2D99E5B8",
    x"2D99D27D",
    x"2D99BF44",
    x"2D99AC0D",
    x"2D9998D9",
    x"2D9985A7",
    x"2D997277",
    x"2D995F4A",
    x"2D994C20",
    x"2D9938F7",
    x"2D9925D1",
    x"2D9912AE",
    x"2D98FF8D",
    x"2D98EC6E",
    x"2D98D952",
    x"2D98C638",
    x"2D98B320",
    x"2D98A00B",
    x"2D988CF8",
    x"2D9879E8",
    x"2D9866DA",
    x"2D9853CE",
    x"2D9840C5",
    x"2D982DBE",
    x"2D981AB9",
    x"2D9807B7",
    x"2D97F4B7",
    x"2D97E1BA",
    x"2D97CEBF",
    x"2D97BBC6",
    x"2D97A8D0",
    x"2D9795DC",
    x"2D9782EA",
    x"2D976FFB",
    x"2D975D0E",
    x"2D974A24",
    x"2D97373C",
    x"2D972456",
    x"2D971173",
    x"2D96FE92",
    x"2D96EBB3",
    x"2D96D8D7",
    x"2D96C5FD",
    x"2D96B325",
    x"2D96A050",
    x"2D968D7D",
    x"2D967AAD",
    x"2D9667DF",
    x"2D965513",
    x"2D964249",
    x"2D962F82",
    x"2D961CBD",
    x"2D9609FB",
    x"2D95F73B",
    x"2D95E47D",
    x"2D95D1C2",
    x"2D95BF09",
    x"2D95AC52",
    x"2D95999E",
    x"2D9586EC",
    x"2D95743C",
    x"2D95618F",
    x"2D954EE4",
    x"2D953C3B",
    x"2D952995",
    x"2D9516F0",
    x"2D95044F",
    x"2D94F1AF",
    x"2D94DF12",
    x"2D94CC78",
    x"2D94B9DF",
    x"2D94A749",
    x"2D9494B5",
    x"2D948224",
    x"2D946F95",
    x"2D945D08",
    x"2D944A7E",
    x"2D9437F5",
    x"2D942570",
    x"2D9412EC",
    x"2D94006B",
    x"2D93EDEC",
    x"2D93DB6F",
    x"2D93C8F5",
    x"2D93B67D",
    x"2D93A408",
    x"2D939194",
    x"2D937F23",
    x"2D936CB4",
    x"2D935A48",
    x"2D9347DE",
    x"2D933576",
    x"2D932310",
    x"2D9310AD",
    x"2D92FE4C",
    x"2D92EBEE",
    x"2D92D991",
    x"2D92C737",
    x"2D92B4DF",
    x"2D92A28A",
    x"2D929037",
    x"2D927DE6",
    x"2D926B97",
    x"2D92594B",
    x"2D924701",
    x"2D9234B9",
    x"2D922274",
    x"2D921031",
    x"2D91FDF0",
    x"2D91EBB1",
    x"2D91D975",
    x"2D91C73B",
    x"2D91B503",
    x"2D91A2CE",
    x"2D91909A",
    x"2D917E69",
    x"2D916C3B",
    x"2D915A0E",
    x"2D9147E4",
    x"2D9135BC",
    x"2D912397",
    x"2D911174",
    x"2D90FF52",
    x"2D90ED34",
    x"2D90DB17",
    x"2D90C8FD",
    x"2D90B6E5",
    x"2D90A4CF",
    x"2D9092BC",
    x"2D9080AB",
    x"2D906E9C",
    x"2D905C8F",
    x"2D904A84",
    x"2D90387C",
    x"2D902676",
    x"2D901473",
    x"2D900271",
    x"2D8FF072",
    x"2D8FDE75",
    x"2D8FCC7A",
    x"2D8FBA82",
    x"2D8FA88C",
    x"2D8F9698",
    x"2D8F84A6",
    x"2D8F72B7",
    x"2D8F60C9",
    x"2D8F4EDE",
    x"2D8F3CF6",
    x"2D8F2B0F",
    x"2D8F192B",
    x"2D8F0749",
    x"2D8EF569",
    x"2D8EE38C",
    x"2D8ED1B0",
    x"2D8EBFD7",
    x"2D8EAE00",
    x"2D8E9C2C",
    x"2D8E8A59",
    x"2D8E7889",
    x"2D8E66BB",
    x"2D8E54EF",
    x"2D8E4326",
    x"2D8E315F",
    x"2D8E1F9A",
    x"2D8E0DD7",
    x"2D8DFC16",
    x"2D8DEA58",
    x"2D8DD89B",
    x"2D8DC6E2",
    x"2D8DB52A",
    x"2D8DA374",
    x"2D8D91C1",
    x"2D8D8010",
    x"2D8D6E61",
    x"2D8D5CB4",
    x"2D8D4B0A",
    x"2D8D3961",
    x"2D8D27BB",
    x"2D8D1618",
    x"2D8D0476",
    x"2D8CF2D6",
    x"2D8CE139",
    x"2D8CCF9E",
    x"2D8CBE05",
    x"2D8CAC6F",
    x"2D8C9ADA",
    x"2D8C8948",
    x"2D8C77B8",
    x"2D8C662A",
    x"2D8C549E",
    x"2D8C4315",
    x"2D8C318D",
    x"2D8C2008",
    x"2D8C0E85",
    x"2D8BFD05",
    x"2D8BEB86",
    x"2D8BDA0A",
    x"2D8BC890",
    x"2D8BB718",
    x"2D8BA5A2",
    x"2D8B942E",
    x"2D8B82BD",
    x"2D8B714E",
    x"2D8B5FE1",
    x"2D8B4E76",
    x"2D8B3D0D",
    x"2D8B2BA6",
    x"2D8B1A42",
    x"2D8B08E0",
    x"2D8AF780",
    x"2D8AE622",
    x"2D8AD4C6",
    x"2D8AC36D",
    x"2D8AB215",
    x"2D8AA0C0",
    x"2D8A8F6D",
    x"2D8A7E1C",
    x"2D8A6CCE",
    x"2D8A5B81",
    x"2D8A4A37",
    x"2D8A38EF",
    x"2D8A27A9",
    x"2D8A1665",
    x"2D8A0523",
    x"2D89F3E3",
    x"2D89E2A6",
    x"2D89D16B",
    x"2D89C032",
    x"2D89AEFB",
    x"2D899DC6",
    x"2D898C93",
    x"2D897B63",
    x"2D896A34",
    x"2D895908",
    x"2D8947DE",
    x"2D8936B6",
    x"2D892591",
    x"2D89146D",
    x"2D89034B",
    x"2D88F22C",
    x"2D88E10F",
    x"2D88CFF4",
    x"2D88BEDB",
    x"2D88ADC4",
    x"2D889CAF",
    x"2D888B9D",
    x"2D887A8D",
    x"2D88697E",
    x"2D885872",
    x"2D884768",
    x"2D883660",
    x"2D88255B",
    x"2D881457",
    x"2D880355",
    x"2D87F256",
    x"2D87E159",
    x"2D87D05E",
    x"2D87BF65",
    x"2D87AE6E",
    x"2D879D79",
    x"2D878C87",
    x"2D877B96",
    x"2D876AA8",
    x"2D8759BB",
    x"2D8748D1",
    x"2D8737E9",
    x"2D872703",
    x"2D87161F",
    x"2D87053E",
    x"2D86F45E",
    x"2D86E381",
    x"2D86D2A5",
    x"2D86C1CC",
    x"2D86B0F5",
    x"2D86A020",
    x"2D868F4D",
    x"2D867E7C",
    x"2D866DAD",
    x"2D865CE0",
    x"2D864C16",
    x"2D863B4D",
    x"2D862A87",
    x"2D8619C3",
    x"2D860901",
    x"2D85F841",
    x"2D85E783",
    x"2D85D6C7",
    x"2D85C60D",
    x"2D85B555",
    x"2D85A4A0",
    x"2D8593EC",
    x"2D85833B",
    x"2D85728B",
    x"2D8561DE",
    x"2D855133",
    x"2D85408A",
    x"2D852FE3",
    x"2D851F3E",
    x"2D850E9B",
    x"2D84FDFA",
    x"2D84ED5B",
    x"2D84DCBF",
    x"2D84CC24",
    x"2D84BB8C",
    x"2D84AAF5",
    x"2D849A61",
    x"2D8489CF",
    x"2D84793E",
    x"2D8468B0",
    x"2D845824",
    x"2D84479A",
    x"2D843712",
    x"2D84268D",
    x"2D841609",
    x"2D840587",
    x"2D83F507",
    x"2D83E48A",
    x"2D83D40E",
    x"2D83C395",
    x"2D83B31D",
    x"2D83A2A8",
    x"2D839235",
    x"2D8381C3",
    x"2D837154",
    x"2D8360E7",
    x"2D83507C",
    x"2D834013",
    x"2D832FAC",
    x"2D831F47",
    x"2D830EE4",
    x"2D82FE83",
    x"2D82EE25",
    x"2D82DDC8",
    x"2D82CD6D",
    x"2D82BD14",
    x"2D82ACBE",
    x"2D829C69",
    x"2D828C17",
    x"2D827BC6",
    x"2D826B78",
    x"2D825B2B",
    x"2D824AE1",
    x"2D823A99",
    x"2D822A52",
    x"2D821A0E",
    x"2D8209CC",
    x"2D81F98C",
    x"2D81E94D",
    x"2D81D911",
    x"2D81C8D7",
    x"2D81B89F",
    x"2D81A869",
    x"2D819835",
    x"2D818803",
    x"2D8177D3",
    x"2D8167A5",
    x"2D815779",
    x"2D81474F",
    x"2D813727",
    x"2D812701",
    x"2D8116DD",
    x"2D8106BC",
    x"2D80F69C",
    x"2D80E67E",
    x"2D80D662",
    x"2D80C648",
    x"2D80B631",
    x"2D80A61B",
    x"2D809607",
    x"2D8085F5",
    x"2D8075E6",
    x"2D8065D8",
    x"2D8055CC",
    x"2D8045C2",
    x"2D8035BB",
    x"2D8025B5",
    x"2D8015B1",
    x"2D8005B0",
    x"2D7FEB60",
    x"2D7FCB64",
    x"2D7FAB6D",
    x"2D7F8B79",
    x"2D7F6B8A",
    x"2D7F4B9F",
    x"2D7F2BB7",
    x"2D7F0BD4",
    x"2D7EEBF4",
    x"2D7ECC19",
    x"2D7EAC41",
    x"2D7E8C6E",
    x"2D7E6C9E",
    x"2D7E4CD2",
    x"2D7E2D0B",
    x"2D7E0D47",
    x"2D7DED87",
    x"2D7DCDCC",
    x"2D7DAE14",
    x"2D7D8E60",
    x"2D7D6EB0",
    x"2D7D4F05",
    x"2D7D2F5D",
    x"2D7D0FB9",
    x"2D7CF019",
    x"2D7CD07D",
    x"2D7CB0E5",
    x"2D7C9150",
    x"2D7C71C0",
    x"2D7C5234",
    x"2D7C32AC",
    x"2D7C1327",
    x"2D7BF3A7",
    x"2D7BD42A",
    x"2D7BB4B2",
    x"2D7B953D",
    x"2D7B75CD",
    x"2D7B5660",
    x"2D7B36F7",
    x"2D7B1792",
    x"2D7AF831",
    x"2D7AD8D4",
    x"2D7AB97B",
    x"2D7A9A26",
    x"2D7A7AD4",
    x"2D7A5B87",
    x"2D7A3C3D",
    x"2D7A1CF8",
    x"2D79FDB6",
    x"2D79DE78",
    x"2D79BF3F",
    x"2D79A009",
    x"2D7980D7",
    x"2D7961A8",
    x"2D79427E",
    x"2D792358",
    x"2D790435",
    x"2D78E517",
    x"2D78C5FC",
    x"2D78A6E5",
    x"2D7887D2",
    x"2D7868C3",
    x"2D7849B8",
    x"2D782AB1",
    x"2D780BAD",
    x"2D77ECAE",
    x"2D77CDB2",
    x"2D77AEBB",
    x"2D778FC7",
    x"2D7770D7",
    x"2D7751EA",
    x"2D773302",
    x"2D77141E",
    x"2D76F53D",
    x"2D76D660",
    x"2D76B787",
    x"2D7698B2",
    x"2D7679E1",
    x"2D765B14",
    x"2D763C4B",
    x"2D761D85",
    x"2D75FEC3",
    x"2D75E005",
    x"2D75C14B",
    x"2D75A295",
    x"2D7583E2",
    x"2D756534",
    x"2D754689",
    x"2D7527E2",
    x"2D75093F",
    x"2D74EAA0",
    x"2D74CC05",
    x"2D74AD6D",
    x"2D748ED9",
    x"2D747049",
    x"2D7451BD",
    x"2D743335",
    x"2D7414B0",
    x"2D73F630",
    x"2D73D7B3",
    x"2D73B93A",
    x"2D739AC4",
    x"2D737C53",
    x"2D735DE5",
    x"2D733F7C",
    x"2D732116",
    x"2D7302B3",
    x"2D72E455",
    x"2D72C5FA",
    x"2D72A7A3",
    x"2D728950",
    x"2D726B01",
    x"2D724CB6",
    x"2D722E6E",
    x"2D72102A",
    x"2D71F1EA",
    x"2D71D3AD",
    x"2D71B575",
    x"2D719740",
    x"2D71790F",
    x"2D715AE2",
    x"2D713CB8",
    x"2D711E93",
    x"2D710071",
    x"2D70E253",
    x"2D70C438",
    x"2D70A621",
    x"2D70880F",
    x"2D7069FF",
    x"2D704BF4",
    x"2D702DEC",
    x"2D700FE9",
    x"2D6FF1E9",
    x"2D6FD3EC",
    x"2D6FB5F4",
    x"2D6F97FF",
    x"2D6F7A0E",
    x"2D6F5C20",
    x"2D6F3E36",
    x"2D6F2051",
    x"2D6F026E",
    x"2D6EE490",
    x"2D6EC6B5",
    x"2D6EA8DE",
    x"2D6E8B0B",
    x"2D6E6D3C",
    x"2D6E4F70",
    x"2D6E31A8",
    x"2D6E13E3",
    x"2D6DF623",
    x"2D6DD866",
    x"2D6DBAAD",
    x"2D6D9CF7",
    x"2D6D7F45",
    x"2D6D6197",
    x"2D6D43ED",
    x"2D6D2646",
    x"2D6D08A3",
    x"2D6CEB04",
    x"2D6CCD69",
    x"2D6CAFD1",
    x"2D6C923D",
    x"2D6C74AC",
    x"2D6C5720",
    x"2D6C3996",
    x"2D6C1C11",
    x"2D6BFE8F",
    x"2D6BE111",
    x"2D6BC397",
    x"2D6BA621",
    x"2D6B88AE",
    x"2D6B6B3E",
    x"2D6B4DD3",
    x"2D6B306B",
    x"2D6B1307",
    x"2D6AF5A6",
    x"2D6AD849",
    x"2D6ABAF0",
    x"2D6A9D9B",
    x"2D6A8049",
    x"2D6A62FB",
    x"2D6A45B0",
    x"2D6A2869",
    x"2D6A0B26",
    x"2D69EDE6",
    x"2D69D0AA",
    x"2D69B372",
    x"2D69963E",
    x"2D69790D",
    x"2D695BDF",
    x"2D693EB6",
    x"2D692190",
    x"2D69046D",
    x"2D68E74E",
    x"2D68CA33",
    x"2D68AD1C",
    x"2D689008",
    x"2D6872F8",
    x"2D6855EB",
    x"2D6838E2",
    x"2D681BDD",
    x"2D67FEDB",
    x"2D67E1DD",
    x"2D67C4E3",
    x"2D67A7EC",
    x"2D678AF9",
    x"2D676E09",
    x"2D67511E",
    x"2D673435",
    x"2D671750",
    x"2D66FA6F",
    x"2D66DD92",
    x"2D66C0B8",
    x"2D66A3E2",
    x"2D66870F",
    x"2D666A40",
    x"2D664D74",
    x"2D6630AD",
    x"2D6613E8",
    x"2D65F728",
    x"2D65DA6A",
    x"2D65BDB1",
    x"2D65A0FB",
    x"2D658449",
    x"2D65679A",
    x"2D654AEF",
    x"2D652E47",
    x"2D6511A3",
    x"2D64F503",
    x"2D64D866",
    x"2D64BBCD",
    x"2D649F37",
    x"2D6482A5",
    x"2D646616",
    x"2D64498B",
    x"2D642D04",
    x"2D641080",
    x"2D63F400",
    x"2D63D783",
    x"2D63BB0A",
    x"2D639E94",
    x"2D638222",
    x"2D6365B4",
    x"2D634949",
    x"2D632CE2",
    x"2D63107E",
    x"2D62F41D",
    x"2D62D7C1",
    x"2D62BB67",
    x"2D629F12",
    x"2D6282C0",
    x"2D626671",
    x"2D624A26",
    x"2D622DDF",
    x"2D62119B",
    x"2D61F55A",
    x"2D61D91D",
    x"2D61BCE4",
    x"2D61A0AE",
    x"2D61847C",
    x"2D61684D",
    x"2D614C22",
    x"2D612FFA",
    x"2D6113D6",
    x"2D60F7B5",
    x"2D60DB98",
    x"2D60BF7E",
    x"2D60A368",
    x"2D608755",
    x"2D606B46",
    x"2D604F3A",
    x"2D603332",
    x"2D60172E",
    x"2D5FFB2C",
    x"2D5FDF2F",
    x"2D5FC335",
    x"2D5FA73E",
    x"2D5F8B4B",
    x"2D5F6F5B",
    x"2D5F536F",
    x"2D5F3786",
    x"2D5F1BA1",
    x"2D5EFFBF",
    x"2D5EE3E1",
    x"2D5EC806",
    x"2D5EAC2F",
    x"2D5E905B",
    x"2D5E748B",
    x"2D5E58BE",
    x"2D5E3CF5",
    x"2D5E212F",
    x"2D5E056D",
    x"2D5DE9AE",
    x"2D5DCDF2",
    x"2D5DB23A",
    x"2D5D9686",
    x"2D5D7AD5",
    x"2D5D5F27",
    x"2D5D437D",
    x"2D5D27D6",
    x"2D5D0C33",
    x"2D5CF093",
    x"2D5CD4F7",
    x"2D5CB95E",
    x"2D5C9DC8",
    x"2D5C8236",
    x"2D5C66A8",
    x"2D5C4B1D",
    x"2D5C2F95",
    x"2D5C1411",
    x"2D5BF890",
    x"2D5BDD13",
    x"2D5BC199",
    x"2D5BA622",
    x"2D5B8AAF",
    x"2D5B6F40",
    x"2D5B53D3",
    x"2D5B386B",
    x"2D5B1D05",
    x"2D5B01A3",
    x"2D5AE645",
    x"2D5ACAEA",
    x"2D5AAF92",
    x"2D5A943E",
    x"2D5A78ED",
    x"2D5A5DA0",
    x"2D5A4256",
    x"2D5A270F",
    x"2D5A0BCC",
    x"2D59F08C",
    x"2D59D550",
    x"2D59BA17",
    x"2D599EE1",
    x"2D5983AF",
    x"2D596880",
    x"2D594D55",
    x"2D59322D",
    x"2D591708",
    x"2D58FBE7",
    x"2D58E0C9",
    x"2D58C5AF",
    x"2D58AA98",
    x"2D588F84",
    x"2D587474",
    x"2D585967",
    x"2D583E5E",
    x"2D582358",
    x"2D580855",
    x"2D57ED56",
    x"2D57D25A",
    x"2D57B761",
    x"2D579C6C",
    x"2D57817A",
    x"2D57668B",
    x"2D574BA0",
    x"2D5730B8",
    x"2D5715D4",
    x"2D56FAF3",
    x"2D56E015",
    x"2D56C53B",
    x"2D56AA64",
    x"2D568F90",
    x"2D5674C0",
    x"2D5659F3",
    x"2D563F2A",
    x"2D562463",
    x"2D5609A1",
    x"2D55EEE1",
    x"2D55D425",
    x"2D55B96C",
    x"2D559EB6",
    x"2D558404",
    x"2D556955",
    x"2D554EAA",
    x"2D553402",
    x"2D55195D",
    x"2D54FEBB",
    x"2D54E41D",
    x"2D54C982",
    x"2D54AEEB",
    x"2D549457",
    x"2D5479C6",
    x"2D545F38",
    x"2D5444AE",
    x"2D542A27",
    x"2D540FA3",
    x"2D53F523",
    x"2D53DAA6",
    x"2D53C02C",
    x"2D53A5B6",
    x"2D538B43",
    x"2D5370D3",
    x"2D535667",
    x"2D533BFE",
    x"2D532198",
    x"2D530735",
    x"2D52ECD6",
    x"2D52D27A",
    x"2D52B821",
    x"2D529DCC",
    x"2D52837A",
    x"2D52692B",
    x"2D524EE0",
    x"2D523497",
    x"2D521A53",
    x"2D520011",
    x"2D51E5D3",
    x"2D51CB97",
    x"2D51B160",
    x"2D51972B",
    x"2D517CFA",
    x"2D5162CC",
    x"2D5148A1",
    x"2D512E7A",
    x"2D511456",
    x"2D50FA35",
    x"2D50E017",
    x"2D50C5FD",
    x"2D50ABE5",
    x"2D5091D2",
    x"2D5077C1",
    x"2D505DB4",
    x"2D5043AA",
    x"2D5029A3",
    x"2D500F9F",
    x"2D4FF59F",
    x"2D4FDBA2",
    x"2D4FC1A8",
    x"2D4FA7B1",
    x"2D4F8DBE",
    x"2D4F73CE",
    x"2D4F59E1",
    x"2D4F3FF7",
    x"2D4F2611",
    x"2D4F0C2E",
    x"2D4EF24E",
    x"2D4ED871",
    x"2D4EBE98",
    x"2D4EA4C2",
    x"2D4E8AEF",
    x"2D4E711F",
    x"2D4E5752",
    x"2D4E3D89",
    x"2D4E23C3",
    x"2D4E0A00",
    x"2D4DF041",
    x"2D4DD684",
    x"2D4DBCCB",
    x"2D4DA315",
    x"2D4D8962",
    x"2D4D6FB3",
    x"2D4D5606",
    x"2D4D3C5D",
    x"2D4D22B7",
    x"2D4D0914",
    x"2D4CEF75",
    x"2D4CD5D9",
    x"2D4CBC3F",
    x"2D4CA2A9",
    x"2D4C8917",
    x"2D4C6F87",
    x"2D4C55FB",
    x"2D4C3C72",
    x"2D4C22EC",
    x"2D4C0969",
    x"2D4BEFE9",
    x"2D4BD66D",
    x"2D4BBCF4",
    x"2D4BA37E",
    x"2D4B8A0B",
    x"2D4B709B",
    x"2D4B572F",
    x"2D4B3DC5",
    x"2D4B245F",
    x"2D4B0AFC",
    x"2D4AF19D",
    x"2D4AD840",
    x"2D4ABEE6",
    x"2D4AA590",
    x"2D4A8C3D",
    x"2D4A72ED",
    x"2D4A59A0",
    x"2D4A4057",
    x"2D4A2710",
    x"2D4A0DCD",
    x"2D49F48D",
    x"2D49DB50",
    x"2D49C216",
    x"2D49A8DF",
    x"2D498FAC",
    x"2D49767B",
    x"2D495D4E",
    x"2D494424",
    x"2D492AFD",
    x"2D4911D9",
    x"2D48F8B9",
    x"2D48DF9B",
    x"2D48C681",
    x"2D48AD6A",
    x"2D489455",
    x"2D487B44",
    x"2D486237",
    x"2D48492C",
    x"2D483024",
    x"2D481720",
    x"2D47FE1F",
    x"2D47E520",
    x"2D47CC25",
    x"2D47B32D",
    x"2D479A38",
    x"2D478147",
    x"2D476858",
    x"2D474F6D",
    x"2D473684",
    x"2D471D9F",
    x"2D4704BD",
    x"2D46EBDE",
    x"2D46D302",
    x"2D46BA29",
    x"2D46A153",
    x"2D468881",
    x"2D466FB1",
    x"2D4656E5",
    x"2D463E1C",
    x"2D462555",
    x"2D460C92",
    x"2D45F3D2",
    x"2D45DB15",
    x"2D45C25B",
    x"2D45A9A5",
    x"2D4590F1",
    x"2D457840",
    x"2D455F93",
    x"2D4546E8",
    x"2D452E41",
    x"2D45159D",
    x"2D44FCFC",
    x"2D44E45E",
    x"2D44CBC3",
    x"2D44B32B",
    x"2D449A96",
    x"2D448204",
    x"2D446975",
    x"2D4450EA",
    x"2D443861",
    x"2D441FDC",
    x"2D440759",
    x"2D43EEDA",
    x"2D43D65D",
    x"2D43BDE4",
    x"2D43A56E",
    x"2D438CFB",
    x"2D43748B",
    x"2D435C1E",
    x"2D4343B4",
    x"2D432B4D",
    x"2D4312E9",
    x"2D42FA88",
    x"2D42E22A",
    x"2D42C9D0",
    x"2D42B178",
    x"2D429923",
    x"2D4280D2",
    x"2D426883",
    x"2D425037",
    x"2D4237EF",
    x"2D421FA9",
    x"2D420767",
    x"2D41EF28",
    x"2D41D6EB",
    x"2D41BEB2",
    x"2D41A67C",
    x"2D418E48",
    x"2D417618",
    x"2D415DEB",
    x"2D4145C0",
    x"2D412D99",
    x"2D411575",
    x"2D40FD54",
    x"2D40E536",
    x"2D40CD1B",
    x"2D40B502",
    x"2D409CED",
    x"2D4084DB",
    x"2D406CCC",
    x"2D4054C0",
    x"2D403CB7",
    x"2D4024B1",
    x"2D400CAE",
    x"2D3FF4AE",
    x"2D3FDCB1",
    x"2D3FC4B6",
    x"2D3FACBF",
    x"2D3F94CB",
    x"2D3F7CDA",
    x"2D3F64EC",
    x"2D3F4D01",
    x"2D3F3519",
    x"2D3F1D34",
    x"2D3F0552",
    x"2D3EED72",
    x"2D3ED596",
    x"2D3EBDBD",
    x"2D3EA5E7",
    x"2D3E8E14",
    x"2D3E7643",
    x"2D3E5E76",
    x"2D3E46AC",
    x"2D3E2EE4",
    x"2D3E1720",
    x"2D3DFF5E",
    x"2D3DE7A0",
    x"2D3DCFE5",
    x"2D3DB82C",
    x"2D3DA077",
    x"2D3D88C4",
    x"2D3D7114",
    x"2D3D5968",
    x"2D3D41BE",
    x"2D3D2A17",
    x"2D3D1273",
    x"2D3CFAD3",
    x"2D3CE335",
    x"2D3CCB9A",
    x"2D3CB402",
    x"2D3C9C6D",
    x"2D3C84DB",
    x"2D3C6D4C",
    x"2D3C55BF",
    x"2D3C3E36",
    x"2D3C26B0",
    x"2D3C0F2D",
    x"2D3BF7AC",
    x"2D3BE02F",
    x"2D3BC8B4",
    x"2D3BB13C",
    x"2D3B99C8",
    x"2D3B8256",
    x"2D3B6AE7",
    x"2D3B537B",
    x"2D3B3C12",
    x"2D3B24AC",
    x"2D3B0D49",
    x"2D3AF5E9",
    x"2D3ADE8C",
    x"2D3AC731",
    x"2D3AAFDA",
    x"2D3A9885",
    x"2D3A8134",
    x"2D3A69E5",
    x"2D3A5299",
    x"2D3A3B50",
    x"2D3A240A",
    x"2D3A0CC7",
    x"2D39F587",
    x"2D39DE4A",
    x"2D39C710",
    x"2D39AFD8",
    x"2D3998A4",
    x"2D398172",
    x"2D396A43",
    x"2D395317",
    x"2D393BEF",
    x"2D3924C8",
    x"2D390DA5",
    x"2D38F685",
    x"2D38DF68",
    x"2D38C84D",
    x"2D38B136",
    x"2D389A21",
    x"2D38830F",
    x"2D386C00",
    x"2D3854F4",
    x"2D383DEB",
    x"2D3826E5",
    x"2D380FE1",
    x"2D37F8E1",
    x"2D37E1E3",
    x"2D37CAE8",
    x"2D37B3F0",
    x"2D379CFB",
    x"2D378609",
    x"2D376F1A",
    x"2D37582D",
    x"2D374144",
    x"2D372A5D",
    x"2D371379",
    x"2D36FC98",
    x"2D36E5BA",
    x"2D36CEDF",
    x"2D36B806",
    x"2D36A131",
    x"2D368A5E",
    x"2D36738E",
    x"2D365CC1",
    x"2D3645F7",
    x"2D362F2F",
    x"2D36186B",
    x"2D3601A9",
    x"2D35EAEB",
    x"2D35D42F",
    x"2D35BD76",
    x"2D35A6BF",
    x"2D35900C",
    x"2D35795B",
    x"2D3562AE",
    x"2D354C03",
    x"2D35355B",
    x"2D351EB5",
    x"2D350813",
    x"2D34F173",
    x"2D34DAD6",
    x"2D34C43D",
    x"2D34ADA5",
    x"2D349711",
    x"2D348080",
    x"2D3469F1",
    x"2D345365",
    x"2D343CDC",
    x"2D342656",
    x"2D340FD3",
    x"2D33F952",
    x"2D33E2D4",
    x"2D33CC59",
    x"2D33B5E1",
    x"2D339F6C",
    x"2D3388F9",
    x"2D33728A",
    x"2D335C1D",
    x"2D3345B3",
    x"2D332F4B",
    x"2D3318E7",
    x"2D330285",
    x"2D32EC26",
    x"2D32D5CA",
    x"2D32BF71",
    x"2D32A91A",
    x"2D3292C6",
    x"2D327C75",
    x"2D326627",
    x"2D324FDC",
    x"2D323993",
    x"2D32234D",
    x"2D320D0A",
    x"2D31F6CA",
    x"2D31E08D",
    x"2D31CA52",
    x"2D31B41A",
    x"2D319DE5",
    x"2D3187B3",
    x"2D317183",
    x"2D315B56",
    x"2D31452C",
    x"2D312F05",
    x"2D3118E1",
    x"2D3102BF",
    x"2D30ECA0",
    x"2D30D684",
    x"2D30C06A",
    x"2D30AA54",
    x"2D309440",
    x"2D307E2F",
    x"2D306820",
    x"2D305214",
    x"2D303C0C",
    x"2D302605",
    x"2D301002",
    x"2D2FFA01",
    x"2D2FE404",
    x"2D2FCE08",
    x"2D2FB810",
    x"2D2FA21A",
    x"2D2F8C28",
    x"2D2F7637",
    x"2D2F604A",
    x"2D2F4A5F",
    x"2D2F3477",
    x"2D2F1E92",
    x"2D2F08B0",
    x"2D2EF2D0",
    x"2D2EDCF3",
    x"2D2EC719",
    x"2D2EB141",
    x"2D2E9B6C",
    x"2D2E859A",
    x"2D2E6FCB",
    x"2D2E59FE",
    x"2D2E4435",
    x"2D2E2E6D",
    x"2D2E18A9",
    x"2D2E02E7",
    x"2D2DED28",
    x"2D2DD76C",
    x"2D2DC1B2",
    x"2D2DABFC",
    x"2D2D9647",
    x"2D2D8096",
    x"2D2D6AE7",
    x"2D2D553B",
    x"2D2D3F92",
    x"2D2D29EB",
    x"2D2D1447",
    x"2D2CFEA6",
    x"2D2CE908",
    x"2D2CD36C",
    x"2D2CBDD3",
    x"2D2CA83D",
    x"2D2C92A9",
    x"2D2C7D18",
    x"2D2C678A",
    x"2D2C51FE",
    x"2D2C3C75",
    x"2D2C26EF",
    x"2D2C116B",
    x"2D2BFBEB",
    x"2D2BE66C",
    x"2D2BD0F1",
    x"2D2BBB78",
    x"2D2BA602",
    x"2D2B908F",
    x"2D2B7B1E",
    x"2D2B65B0",
    x"2D2B5045",
    x"2D2B3ADC",
    x"2D2B2576",
    x"2D2B1012",
    x"2D2AFAB2",
    x"2D2AE554",
    x"2D2ACFF8",
    x"2D2ABAA0",
    x"2D2AA54A",
    x"2D2A8FF6",
    x"2D2A7AA6",
    x"2D2A6558",
    x"2D2A500C",
    x"2D2A3AC4",
    x"2D2A257E",
    x"2D2A103A",
    x"2D29FAFA",
    x"2D29E5BC",
    x"2D29D080",
    x"2D29BB48",
    x"2D29A611",
    x"2D2990DE",
    x"2D297BAD",
    x"2D29667F",
    x"2D295154",
    x"2D293C2B",
    x"2D292705",
    x"2D2911E1",
    x"2D28FCC0",
    x"2D28E7A2",
    x"2D28D286",
    x"2D28BD6D",
    x"2D28A857",
    x"2D289343",
    x"2D287E32",
    x"2D286924",
    x"2D285418",
    x"2D283F0F",
    x"2D282A08",
    x"2D281504",
    x"2D280003",
    x"2D27EB04",
    x"2D27D608",
    x"2D27C10F",
    x"2D27AC18",
    x"2D279723",
    x"2D278232",
    x"2D276D43",
    x"2D275857",
    x"2D27436D",
    x"2D272E86",
    x"2D2719A1",
    x"2D2704BF",
    x"2D26EFE0",
    x"2D26DB03",
    x"2D26C629",
    x"2D26B152",
    x"2D269C7D",
    x"2D2687AB",
    x"2D2672DB",
    x"2D265E0E",
    x"2D264944",
    x"2D26347C",
    x"2D261FB6",
    x"2D260AF4",
    x"2D25F634",
    x"2D25E176",
    x"2D25CCBB",
    x"2D25B803",
    x"2D25A34D",
    x"2D258E9A",
    x"2D2579EA",
    x"2D25653C",
    x"2D255090",
    x"2D253BE8",
    x"2D252741",
    x"2D25129E",
    x"2D24FDFD",
    x"2D24E95E",
    x"2D24D4C2",
    x"2D24C029",
    x"2D24AB92",
    x"2D2496FE",
    x"2D24826D",
    x"2D246DDE",
    x"2D245951",
    x"2D2444C7",
    x"2D243040",
    x"2D241BBB",
    x"2D240739",
    x"2D23F2B9",
    x"2D23DE3C",
    x"2D23C9C2",
    x"2D23B54A",
    x"2D23A0D4",
    x"2D238C62",
    x"2D2377F1",
    x"2D236384",
    x"2D234F19",
    x"2D233AB0",
    x"2D23264A",
    x"2D2311E6",
    x"2D22FD85",
    x"2D22E927",
    x"2D22D4CB",
    x"2D22C072",
    x"2D22AC1B",
    x"2D2297C7",
    x"2D228375",
    x"2D226F26",
    x"2D225AD9",
    x"2D22468F",
    x"2D223248",
    x"2D221E03",
    x"2D2209C0",
    x"2D21F580",
    x"2D21E143",
    x"2D21CD08",
    x"2D21B8CF",
    x"2D21A49A",
    x"2D219066",
    x"2D217C36",
    x"2D216807",
    x"2D2153DB",
    x"2D213FB2",
    x"2D212B8C",
    x"2D211767",
    x"2D210346",
    x"2D20EF27",
    x"2D20DB0A",
    x"2D20C6F0",
    x"2D20B2D8",
    x"2D209EC3",
    x"2D208AB1",
    x"2D2076A0",
    x"2D206293",
    x"2D204E88",
    x"2D203A7F",
    x"2D202679",
    x"2D201276",
    x"2D1FFE75",
    x"2D1FEA76",
    x"2D1FD67A",
    x"2D1FC280",
    x"2D1FAE89",
    x"2D1F9A95",
    x"2D1F86A3",
    x"2D1F72B3",
    x"2D1F5EC6",
    x"2D1F4ADB",
    x"2D1F36F3",
    x"2D1F230E",
    x"2D1F0F2B",
    x"2D1EFB4A",
    x"2D1EE76C",
    x"2D1ED390",
    x"2D1EBFB7",
    x"2D1EABE0",
    x"2D1E980C",
    x"2D1E843A",
    x"2D1E706B",
    x"2D1E5C9E",
    x"2D1E48D4",
    x"2D1E350C",
    x"2D1E2146",
    x"2D1E0D83",
    x"2D1DF9C3",
    x"2D1DE605",
    x"2D1DD249",
    x"2D1DBE90",
    x"2D1DAADA",
    x"2D1D9726",
    x"2D1D8374",
    x"2D1D6FC5",
    x"2D1D5C18",
    x"2D1D486E",
    x"2D1D34C6",
    x"2D1D2121",
    x"2D1D0D7E",
    x"2D1CF9DD",
    x"2D1CE63F",
    x"2D1CD2A4",
    x"2D1CBF0B",
    x"2D1CAB74",
    x"2D1C97E0",
    x"2D1C844E",
    x"2D1C70BF",
    x"2D1C5D32",
    x"2D1C49A7",
    x"2D1C361F",
    x"2D1C229A",
    x"2D1C0F17",
    x"2D1BFB96",
    x"2D1BE818",
    x"2D1BD49C",
    x"2D1BC123",
    x"2D1BADAC",
    x"2D1B9A37",
    x"2D1B86C5",
    x"2D1B7356",
    x"2D1B5FE8",
    x"2D1B4C7E",
    x"2D1B3915",
    x"2D1B25AF",
    x"2D1B124C",
    x"2D1AFEEB",
    x"2D1AEB8C",
    x"2D1AD830",
    x"2D1AC4D6",
    x"2D1AB17F",
    x"2D1A9E2A",
    x"2D1A8AD7",
    x"2D1A7787",
    x"2D1A6439",
    x"2D1A50EE",
    x"2D1A3DA5",
    x"2D1A2A5E",
    x"2D1A171A",
    x"2D1A03D9",
    x"2D19F099",
    x"2D19DD5D",
    x"2D19CA22",
    x"2D19B6EA",
    x"2D19A3B4",
    x"2D199081",
    x"2D197D50",
    x"2D196A22",
    x"2D1956F6",
    x"2D1943CC",
    x"2D1930A5",
    x"2D191D80",
    x"2D190A5D",
    x"2D18F73D",
    x"2D18E420",
    x"2D18D104",
    x"2D18BDEB",
    x"2D18AAD5",
    x"2D1897C1",
    x"2D1884AF",
    x"2D18719F",
    x"2D185E92",
    x"2D184B88",
    x"2D183880",
    x"2D18257A",
    x"2D181276",
    x"2D17FF75",
    x"2D17EC76",
    x"2D17D97A",
    x"2D17C680",
    x"2D17B388",
    x"2D17A093",
    x"2D178DA0",
    x"2D177AB0",
    x"2D1767C1",
    x"2D1754D6",
    x"2D1741EC",
    x"2D172F05",
    x"2D171C21",
    x"2D17093E",
    x"2D16F65E",
    x"2D16E381",
    x"2D16D0A5",
    x"2D16BDCC",
    x"2D16AAF6",
    x"2D169822",
    x"2D168550",
    x"2D167280",
    x"2D165FB3",
    x"2D164CE8",
    x"2D163A20",
    x"2D16275A",
    x"2D161496",
    x"2D1601D5",
    x"2D15EF16",
    x"2D15DC59",
    x"2D15C99F",
    x"2D15B6E7",
    x"2D15A431",
    x"2D15917E",
    x"2D157ECC",
    x"2D156C1E",
    x"2D155971",
    x"2D1546C7",
    x"2D153420",
    x"2D15217A",
    x"2D150ED7",
    x"2D14FC37",
    x"2D14E998",
    x"2D14D6FC",
    x"2D14C463",
    x"2D14B1CB",
    x"2D149F36",
    x"2D148CA3",
    x"2D147A13",
    x"2D146785",
    x"2D1454F9",
    x"2D144270",
    x"2D142FE9",
    x"2D141D64",
    x"2D140AE1",
    x"2D13F861",
    x"2D13E5E3",
    x"2D13D367",
    x"2D13C0EE",
    x"2D13AE77",
    x"2D139C03",
    x"2D138990",
    x"2D137720",
    x"2D1364B2",
    x"2D135247",
    x"2D133FDE",
    x"2D132D77",
    x"2D131B13",
    x"2D1308B0",
    x"2D12F650",
    x"2D12E3F3",
    x"2D12D197",
    x"2D12BF3E",
    x"2D12ACE8",
    x"2D129A93",
    x"2D128841",
    x"2D1275F1",
    x"2D1263A3",
    x"2D125158",
    x"2D123F0F",
    x"2D122CC8",
    x"2D121A84",
    x"2D120842",
    x"2D11F602",
    x"2D11E3C4",
    x"2D11D189",
    x"2D11BF50",
    x"2D11AD19",
    x"2D119AE5",
    x"2D1188B2",
    x"2D117682",
    x"2D116455",
    x"2D115229",
    x"2D114000",
    x"2D112DD9",
    x"2D111BB5",
    x"2D110992",
    x"2D10F772",
    x"2D10E555",
    x"2D10D339",
    x"2D10C120",
    x"2D10AF09",
    x"2D109CF4",
    x"2D108AE1",
    x"2D1078D1",
    x"2D1066C3",
    x"2D1054B8",
    x"2D1042AE",
    x"2D1030A7",
    x"2D101EA2",
    x"2D100C9F",
    x"2D0FFA9F",
    x"2D0FE8A1",
    x"2D0FD6A5",
    x"2D0FC4AB",
    x"2D0FB2B3",
    x"2D0FA0BE",
    x"2D0F8ECB",
    x"2D0F7CDB",
    x"2D0F6AEC",
    x"2D0F5900",
    x"2D0F4716",
    x"2D0F352E",
    x"2D0F2348",
    x"2D0F1165",
    x"2D0EFF84",
    x"2D0EEDA5",
    x"2D0EDBC9",
    x"2D0EC9EE",
    x"2D0EB816",
    x"2D0EA640",
    x"2D0E946D",
    x"2D0E829B",
    x"2D0E70CC",
    x"2D0E5EFF",
    x"2D0E4D34",
    x"2D0E3B6C",
    x"2D0E29A5",
    x"2D0E17E1",
    x"2D0E061F",
    x"2D0DF460",
    x"2D0DE2A2",
    x"2D0DD0E7",
    x"2D0DBF2E",
    x"2D0DAD77",
    x"2D0D9BC3",
    x"2D0D8A10",
    x"2D0D7860",
    x"2D0D66B2",
    x"2D0D5507",
    x"2D0D435D",
    x"2D0D31B6",
    x"2D0D2011",
    x"2D0D0E6E",
    x"2D0CFCCD",
    x"2D0CEB2F",
    x"2D0CD992",
    x"2D0CC7F8",
    x"2D0CB660",
    x"2D0CA4CB",
    x"2D0C9337",
    x"2D0C81A6",
    x"2D0C7017",
    x"2D0C5E8A",
    x"2D0C4CFF",
    x"2D0C3B76",
    x"2D0C29F0",
    x"2D0C186C",
    x"2D0C06EA",
    x"2D0BF56A",
    x"2D0BE3ED",
    x"2D0BD271",
    x"2D0BC0F8",
    x"2D0BAF81",
    x"2D0B9E0C",
    x"2D0B8C9A",
    x"2D0B7B29",
    x"2D0B69BB",
    x"2D0B584F",
    x"2D0B46E5",
    x"2D0B357D",
    x"2D0B2417",
    x"2D0B12B4",
    x"2D0B0153",
    x"2D0AEFF4",
    x"2D0ADE97",
    x"2D0ACD3C",
    x"2D0ABBE3",
    x"2D0AAA8D",
    x"2D0A9939",
    x"2D0A87E7",
    x"2D0A7697",
    x"2D0A6549",
    x"2D0A53FD",
    x"2D0A42B4",
    x"2D0A316D",
    x"2D0A2028",
    x"2D0A0EE5",
    x"2D09FDA4",
    x"2D09EC65",
    x"2D09DB29",
    x"2D09C9EE",
    x"2D09B8B6",
    x"2D09A780",
    x"2D09964C",
    x"2D09851B",
    x"2D0973EB",
    x"2D0962BE",
    x"2D095192",
    x"2D094069",
    x"2D092F42",
    x"2D091E1D",
    x"2D090CFB",
    x"2D08FBDA",
    x"2D08EABC",
    x"2D08D9A0",
    x"2D08C885",
    x"2D08B76D",
    x"2D08A658",
    x"2D089544",
    x"2D088432",
    x"2D087323",
    x"2D086215",
    x"2D08510A",
    x"2D084001",
    x"2D082EFA",
    x"2D081DF5",
    x"2D080CF3",
    x"2D07FBF2",
    x"2D07EAF4",
    x"2D07D9F7",
    x"2D07C8FD",
    x"2D07B805",
    x"2D07A70F",
    x"2D07961B",
    x"2D07852A",
    x"2D07743A",
    x"2D07634D",
    x"2D075261",
    x"2D074178",
    x"2D073091",
    x"2D071FAC",
    x"2D070EC9",
    x"2D06FDE8",
    x"2D06ED0A",
    x"2D06DC2D",
    x"2D06CB53",
    x"2D06BA7A",
    x"2D06A9A4",
    x"2D0698D0",
    x"2D0687FE",
    x"2D06772E",
    x"2D066660",
    x"2D065594",
    x"2D0644CB",
    x"2D063403",
    x"2D06233E",
    x"2D06127A",
    x"2D0601B9",
    x"2D05F0FA",
    x"2D05E03D",
    x"2D05CF82",
    x"2D05BEC9",
    x"2D05AE12",
    x"2D059D5D",
    x"2D058CAB",
    x"2D057BFA",
    x"2D056B4C",
    x"2D055A9F",
    x"2D0549F5",
    x"2D05394D",
    x"2D0528A7",
    x"2D051803",
    x"2D050761",
    x"2D04F6C1",
    x"2D04E623",
    x"2D04D587",
    x"2D04C4EE",
    x"2D04B456",
    x"2D04A3C1",
    x"2D04932D",
    x"2D04829C",
    x"2D04720C",
    x"2D04617F",
    x"2D0450F4",
    x"2D04406B",
    x"2D042FE4",
    x"2D041F5F",
    x"2D040EDC",
    x"2D03FE5B",
    x"2D03EDDD",
    x"2D03DD60",
    x"2D03CCE5",
    x"2D03BC6D",
    x"2D03ABF6",
    x"2D039B82",
    x"2D038B0F",
    x"2D037A9F",
    x"2D036A31",
    x"2D0359C4",
    x"2D03495A",
    x"2D0338F2",
    x"2D03288C",
    x"2D031828",
    x"2D0307C6",
    x"2D02F766",
    x"2D02E708",
    x"2D02D6AC",
    x"2D02C652",
    x"2D02B5FB",
    x"2D02A5A5",
    x"2D029551",
    x"2D0284FF",
    x"2D0274B0",
    x"2D026462",
    x"2D025417",
    x"2D0243CD",
    x"2D023386",
    x"2D022340",
    x"2D0212FD",
    x"2D0202BC",
    x"2D01F27C",
    x"2D01E23F",
    x"2D01D204",
    x"2D01C1CB",
    x"2D01B193",
    x"2D01A15E",
    x"2D01912B",
    x"2D0180FA",
    x"2D0170CB",
    x"2D01609E",
    x"2D015073",
    x"2D01404A",
    x"2D013023",
    x"2D011FFE",
    x"2D010FDB",
    x"2D00FFBA",
    x"2D00EF9B",
    x"2D00DF7E",
    x"2D00CF63",
    x"2D00BF4A",
    x"2D00AF33",
    x"2D009F1E",
    x"2D008F0B",
    x"2D007EFA",
    x"2D006EEB",
    x"2D005EDE",
    x"2D004ED4",
    x"2D003ECB",
    x"2D002EC4",
    x"2D001EBF",
    x"2D000EBC",
    x"2CFFFD77",
    x"2CFFDD79",
    x"2CFFBD7F",
    x"2CFF9D8A",
    x"2CFF7D98",
    x"2CFF5DAA",
    x"2CFF3DC1",
    x"2CFF1DDB",
    x"2CFEFDF9",
    x"2CFEDE1B",
    x"2CFEBE42",
    x"2CFE9E6C",
    x"2CFE7E9A",
    x"2CFE5ECC",
    x"2CFE3F02",
    x"2CFE1F3C",
    x"2CFDFF7B",
    x"2CFDDFBD",
    x"2CFDC003",
    x"2CFDA04D",
    x"2CFD809B",
    x"2CFD60EC",
    x"2CFD4142",
    x"2CFD219C",
    x"2CFD01FA",
    x"2CFCE25C",
    x"2CFCC2C1",
    x"2CFCA32B",
    x"2CFC8399",
    x"2CFC640A",
    x"2CFC4480",
    x"2CFC24F9",
    x"2CFC0576",
    x"2CFBE5F8",
    x"2CFBC67D",
    x"2CFBA706",
    x"2CFB8793",
    x"2CFB6824",
    x"2CFB48B9",
    x"2CFB2952",
    x"2CFB09EF",
    x"2CFAEA8F",
    x"2CFACB34",
    x"2CFAABDD",
    x"2CFA8C89",
    x"2CFA6D39",
    x"2CFA4DEE",
    x"2CFA2EA6",
    x"2CFA0F62",
    x"2CF9F022",
    x"2CF9D0E6",
    x"2CF9B1AE",
    x"2CF9927A",
    x"2CF97349",
    x"2CF9541D",
    x"2CF934F4",
    x"2CF915D0",
    x"2CF8F6AF",
    x"2CF8D792",
    x"2CF8B879",
    x"2CF89964",
    x"2CF87A53",
    x"2CF85B45",
    x"2CF83C3C",
    x"2CF81D36",
    x"2CF7FE34",
    x"2CF7DF37",
    x"2CF7C03D",
    x"2CF7A147",
    x"2CF78254",
    x"2CF76366",
    x"2CF7447B",
    x"2CF72595",
    x"2CF706B2",
    x"2CF6E7D3",
    x"2CF6C8F8",
    x"2CF6AA21",
    x"2CF68B4E",
    x"2CF66C7E",
    x"2CF64DB2",
    x"2CF62EEB",
    x"2CF61027",
    x"2CF5F167",
    x"2CF5D2AA",
    x"2CF5B3F2",
    x"2CF5953D",
    x"2CF5768D",
    x"2CF557E0",
    x"2CF53937",
    x"2CF51A91",
    x"2CF4FBF0",
    x"2CF4DD52",
    x"2CF4BEB9",
    x"2CF4A023",
    x"2CF48191",
    x"2CF46302",
    x"2CF44478",
    x"2CF425F1",
    x"2CF4076E",
    x"2CF3E8EF",
    x"2CF3CA74",
    x"2CF3ABFD",
    x"2CF38D89",
    x"2CF36F19",
    x"2CF350AD",
    x"2CF33245",
    x"2CF313E1",
    x"2CF2F580",
    x"2CF2D723",
    x"2CF2B8CA",
    x"2CF29A75",
    x"2CF27C24",
    x"2CF25DD6",
    x"2CF23F8C",
    x"2CF22146",
    x"2CF20304",
    x"2CF1E4C6",
    x"2CF1C68B",
    x"2CF1A854",
    x"2CF18A21",
    x"2CF16BF1",
    x"2CF14DC6",
    x"2CF12F9E",
    x"2CF1117A",
    x"2CF0F35A",
    x"2CF0D53D",
    x"2CF0B724",
    x"2CF0990F",
    x"2CF07AFE",
    x"2CF05CF1",
    x"2CF03EE7",
    x"2CF020E1",
    x"2CF002DF",
    x"2CEFE4E0",
    x"2CEFC6E5",
    x"2CEFA8EE",
    x"2CEF8AFB",
    x"2CEF6D0C",
    x"2CEF4F20",
    x"2CEF3138",
    x"2CEF1354",
    x"2CEEF573",
    x"2CEED796",
    x"2CEEB9BD",
    x"2CEE9BE8",
    x"2CEE7E16",
    x"2CEE6048",
    x"2CEE427E",
    x"2CEE24B8",
    x"2CEE06F5",
    x"2CEDE936",
    x"2CEDCB7B",
    x"2CEDADC3",
    x"2CED900F",
    x"2CED725F",
    x"2CED54B3",
    x"2CED370A",
    x"2CED1965",
    x"2CECFBC3",
    x"2CECDE26",
    x"2CECC08C",
    x"2CECA2F6",
    x"2CEC8563",
    x"2CEC67D4",
    x"2CEC4A49",
    x"2CEC2CC2",
    x"2CEC0F3E",
    x"2CEBF1BE",
    x"2CEBD442",
    x"2CEBB6C9",
    x"2CEB9954",
    x"2CEB7BE3",
    x"2CEB5E75",
    x"2CEB410B",
    x"2CEB23A5",
    x"2CEB0642",
    x"2CEAE8E3",
    x"2CEACB88",
    x"2CEAAE30",
    x"2CEA90DC",
    x"2CEA738C",
    x"2CEA563F",
    x"2CEA38F6",
    x"2CEA1BB1",
    x"2CE9FE70",
    x"2CE9E132",
    x"2CE9C3F7",
    x"2CE9A6C1",
    x"2CE9898E",
    x"2CE96C5E",
    x"2CE94F32",
    x"2CE9320A",
    x"2CE914E6",
    x"2CE8F7C5",
    x"2CE8DAA8",
    x"2CE8BD8E",
    x"2CE8A079",
    x"2CE88366",
    x"2CE86658",
    x"2CE8494D",
    x"2CE82C45",
    x"2CE80F42",
    x"2CE7F242",
    x"2CE7D545",
    x"2CE7B84C",
    x"2CE79B57",
    x"2CE77E65",
    x"2CE76177",
    x"2CE7448D",
    x"2CE727A6",
    x"2CE70AC3",
    x"2CE6EDE4",
    x"2CE6D108",
    x"2CE6B42F",
    x"2CE6975B",
    x"2CE67A8A",
    x"2CE65DBC",
    x"2CE640F2",
    x"2CE6242C",
    x"2CE60769",
    x"2CE5EAAA",
    x"2CE5CDEE",
    x"2CE5B136",
    x"2CE59482",
    x"2CE577D1",
    x"2CE55B24",
    x"2CE53E7B",
    x"2CE521D5",
    x"2CE50532",
    x"2CE4E893",
    x"2CE4CBF8",
    x"2CE4AF60",
    x"2CE492CC",
    x"2CE4763C",
    x"2CE459AF",
    x"2CE43D25",
    x"2CE4209F",
    x"2CE4041D",
    x"2CE3E79E",
    x"2CE3CB23",
    x"2CE3AEAB",
    x"2CE39237",
    x"2CE375C7",
    x"2CE3595A",
    x"2CE33CF1",
    x"2CE3208B",
    x"2CE30428",
    x"2CE2E7CA",
    x"2CE2CB6E",
    x"2CE2AF17",
    x"2CE292C3",
    x"2CE27672",
    x"2CE25A25",
    x"2CE23DDC",
    x"2CE22196",
    x"2CE20553",
    x"2CE1E914",
    x"2CE1CCD9",
    x"2CE1B0A1",
    x"2CE1946D",
    x"2CE1783C",
    x"2CE15C0F",
    x"2CE13FE5",
    x"2CE123BF",
    x"2CE1079C",
    x"2CE0EB7D",
    x"2CE0CF61",
    x"2CE0B349",
    x"2CE09734",
    x"2CE07B23",
    x"2CE05F16",
    x"2CE0430B",
    x"2CE02705",
    x"2CE00B02",
    x"2CDFEF02",
    x"2CDFD306",
    x"2CDFB70D",
    x"2CDF9B18",
    x"2CDF7F26",
    x"2CDF6338",
    x"2CDF474E",
    x"2CDF2B66",
    x"2CDF0F83",
    x"2CDEF3A3",
    x"2CDED7C6",
    x"2CDEBBED",
    x"2CDEA017",
    x"2CDE8445",
    x"2CDE6876",
    x"2CDE4CAB",
    x"2CDE30E3",
    x"2CDE151E",
    x"2CDDF95D",
    x"2CDDDDA0",
    x"2CDDC1E6",
    x"2CDDA62F",
    x"2CDD8A7C",
    x"2CDD6ECD",
    x"2CDD5321",
    x"2CDD3778",
    x"2CDD1BD3",
    x"2CDD0031",
    x"2CDCE493",
    x"2CDCC8F8",
    x"2CDCAD61",
    x"2CDC91CD",
    x"2CDC763C",
    x"2CDC5AAF",
    x"2CDC3F25",
    x"2CDC239F",
    x"2CDC081D",
    x"2CDBEC9D",
    x"2CDBD121",
    x"2CDBB5A9",
    x"2CDB9A34",
    x"2CDB7EC2",
    x"2CDB6354",
    x"2CDB47EA",
    x"2CDB2C82",
    x"2CDB111E",
    x"2CDAF5BE",
    x"2CDADA61",
    x"2CDABF07",
    x"2CDAA3B1",
    x"2CDA885F",
    x"2CDA6D0F",
    x"2CDA51C3",
    x"2CDA367B",
    x"2CDA1B36",
    x"2CD9FFF4",
    x"2CD9E4B6",
    x"2CD9C97B",
    x"2CD9AE43",
    x"2CD9930F",
    x"2CD977DF",
    x"2CD95CB1",
    x"2CD94187",
    x"2CD92661",
    x"2CD90B3E",
    x"2CD8F01E",
    x"2CD8D502",
    x"2CD8B9E9",
    x"2CD89ED3",
    x"2CD883C1",
    x"2CD868B2",
    x"2CD84DA7",
    x"2CD8329F",
    x"2CD8179A",
    x"2CD7FC99",
    x"2CD7E19B",
    x"2CD7C6A1",
    x"2CD7ABA9",
    x"2CD790B6",
    x"2CD775C5",
    x"2CD75AD8",
    x"2CD73FEF",
    x"2CD72508",
    x"2CD70A25",
    x"2CD6EF46",
    x"2CD6D469",
    x"2CD6B991",
    x"2CD69EBB",
    x"2CD683E9",
    x"2CD6691A",
    x"2CD64E4F",
    x"2CD63387",
    x"2CD618C2",
    x"2CD5FE00",
    x"2CD5E342",
    x"2CD5C888",
    x"2CD5ADD0",
    x"2CD5931C",
    x"2CD5786B",
    x"2CD55DBE",
    x"2CD54314",
    x"2CD5286D",
    x"2CD50DCA",
    x"2CD4F32A",
    x"2CD4D88D",
    x"2CD4BDF4",
    x"2CD4A35E",
    x"2CD488CB",
    x"2CD46E3B",
    x"2CD453AF",
    x"2CD43926",
    x"2CD41EA1",
    x"2CD4041F",
    x"2CD3E9A0",
    x"2CD3CF24",
    x"2CD3B4AC",
    x"2CD39A37",
    x"2CD37FC6",
    x"2CD36557",
    x"2CD34AEC",
    x"2CD33084",
    x"2CD31620",
    x"2CD2FBBF",
    x"2CD2E161",
    x"2CD2C707",
    x"2CD2ACAF",
    x"2CD2925B",
    x"2CD2780B",
    x"2CD25DBD",
    x"2CD24373",
    x"2CD2292D",
    x"2CD20EE9",
    x"2CD1F4A9",
    x"2CD1DA6C",
    x"2CD1C032",
    x"2CD1A5FC",
    x"2CD18BC9",
    x"2CD17199",
    x"2CD1576C",
    x"2CD13D43",
    x"2CD1231D",
    x"2CD108FA",
    x"2CD0EEDB",
    x"2CD0D4BF",
    x"2CD0BAA6",
    x"2CD0A090",
    x"2CD0867D",
    x"2CD06C6E",
    x"2CD05262",
    x"2CD0385A",
    x"2CD01E54",
    x"2CD00452",
    x"2CCFEA53",
    x"2CCFD058",
    x"2CCFB65F",
    x"2CCF9C6A",
    x"2CCF8278",
    x"2CCF6889",
    x"2CCF4E9E",
    x"2CCF34B6",
    x"2CCF1AD1",
    x"2CCF00EF",
    x"2CCEE710",
    x"2CCECD35",
    x"2CCEB35D",
    x"2CCE9988",
    x"2CCE7FB7",
    x"2CCE65E8",
    x"2CCE4C1D",
    x"2CCE3255",
    x"2CCE1891",
    x"2CCDFECF",
    x"2CCDE511",
    x"2CCDCB56",
    x"2CCDB19E",
    x"2CCD97EA",
    x"2CCD7E38",
    x"2CCD648A",
    x"2CCD4ADF",
    x"2CCD3137",
    x"2CCD1793",
    x"2CCCFDF1",
    x"2CCCE453",
    x"2CCCCAB8",
    x"2CCCB121",
    x"2CCC978C",
    x"2CCC7DFB",
    x"2CCC646D",
    x"2CCC4AE2",
    x"2CCC315A",
    x"2CCC17D5",
    x"2CCBFE54",
    x"2CCBE4D6",
    x"2CCBCB5B",
    x"2CCBB1E3",
    x"2CCB986E",
    x"2CCB7EFD",
    x"2CCB658E",
    x"2CCB4C23",
    x"2CCB32BB",
    x"2CCB1957",
    x"2CCAFFF5",
    x"2CCAE697",
    x"2CCACD3B",
    x"2CCAB3E3",
    x"2CCA9A8E",
    x"2CCA813D",
    x"2CCA67EE",
    x"2CCA4EA3",
    x"2CCA355A",
    x"2CCA1C15",
    x"2CCA02D3",
    x"2CC9E995",
    x"2CC9D059",
    x"2CC9B721",
    x"2CC99DEB",
    x"2CC984B9",
    x"2CC96B8A",
    x"2CC9525E",
    x"2CC93935",
    x"2CC92010",
    x"2CC906ED",
    x"2CC8EDCE",
    x"2CC8D4B2",
    x"2CC8BB99",
    x"2CC8A283",
    x"2CC88970",
    x"2CC87061",
    x"2CC85754",
    x"2CC83E4B",
    x"2CC82545",
    x"2CC80C42",
    x"2CC7F342",
    x"2CC7DA45",
    x"2CC7C14B",
    x"2CC7A854",
    x"2CC78F61",
    x"2CC77671",
    x"2CC75D83",
    x"2CC74499",
    x"2CC72BB2",
    x"2CC712CE",
    x"2CC6F9EE",
    x"2CC6E110",
    x"2CC6C835",
    x"2CC6AF5E",
    x"2CC69689",
    x"2CC67DB8",
    x"2CC664EA",
    x"2CC64C1F",
    x"2CC63357",
    x"2CC61A92",
    x"2CC601D0",
    x"2CC5E912",
    x"2CC5D056",
    x"2CC5B79E",
    x"2CC59EE8",
    x"2CC58636",
    x"2CC56D87",
    x"2CC554DA",
    x"2CC53C31",
    x"2CC5238B",
    x"2CC50AE8",
    x"2CC4F249",
    x"2CC4D9AC",
    x"2CC4C112",
    x"2CC4A87C",
    x"2CC48FE8",
    x"2CC47758",
    x"2CC45ECA",
    x"2CC44640",
    x"2CC42DB9",
    x"2CC41535",
    x"2CC3FCB3",
    x"2CC3E435",
    x"2CC3CBBA",
    x"2CC3B342",
    x"2CC39ACE",
    x"2CC3825C",
    x"2CC369ED",
    x"2CC35181",
    x"2CC33919",
    x"2CC320B3",
    x"2CC30850",
    x"2CC2EFF1",
    x"2CC2D794",
    x"2CC2BF3B",
    x"2CC2A6E5",
    x"2CC28E91",
    x"2CC27641",
    x"2CC25DF4",
    x"2CC245A9",
    x"2CC22D62",
    x"2CC2151E",
    x"2CC1FCDD",
    x"2CC1E49F",
    x"2CC1CC64",
    x"2CC1B42C",
    x"2CC19BF7",
    x"2CC183C5",
    x"2CC16B96",
    x"2CC1536A",
    x"2CC13B41",
    x"2CC1231B",
    x"2CC10AF8",
    x"2CC0F2D8",
    x"2CC0DABC",
    x"2CC0C2A2",
    x"2CC0AA8B",
    x"2CC09277",
    x"2CC07A66",
    x"2CC06258",
    x"2CC04A4E",
    x"2CC03246",
    x"2CC01A41",
    x"2CC0023F",
    x"2CBFEA41",
    x"2CBFD245",
    x"2CBFBA4C",
    x"2CBFA256",
    x"2CBF8A63",
    x"2CBF7274",
    x"2CBF5A87",
    x"2CBF429D",
    x"2CBF2AB6",
    x"2CBF12D2",
    x"2CBEFAF1",
    x"2CBEE314",
    x"2CBECB39",
    x"2CBEB361",
    x"2CBE9B8C",
    x"2CBE83BA",
    x"2CBE6BEB",
    x"2CBE541F",
    x"2CBE3C56",
    x"2CBE2490",
    x"2CBE0CCD",
    x"2CBDF50D",
    x"2CBDDD4F",
    x"2CBDC595",
    x"2CBDADDE",
    x"2CBD962A",
    x"2CBD7E79",
    x"2CBD66CA",
    x"2CBD4F1F",
    x"2CBD3776",
    x"2CBD1FD1",
    x"2CBD082E",
    x"2CBCF08F",
    x"2CBCD8F2",
    x"2CBCC159",
    x"2CBCA9C2",
    x"2CBC922E",
    x"2CBC7A9D",
    x"2CBC6310",
    x"2CBC4B85",
    x"2CBC33FD",
    x"2CBC1C78",
    x"2CBC04F6",
    x"2CBBED76",
    x"2CBBD5FA",
    x"2CBBBE81",
    x"2CBBA70B",
    x"2CBB8F97",
    x"2CBB7827",
    x"2CBB60B9",
    x"2CBB494E",
    x"2CBB31E7",
    x"2CBB1A82",
    x"2CBB0320",
    x"2CBAEBC1",
    x"2CBAD465",
    x"2CBABD0C",
    x"2CBAA5B6",
    x"2CBA8E63",
    x"2CBA7712",
    x"2CBA5FC5",
    x"2CBA487A",
    x"2CBA3133",
    x"2CBA19EE",
    x"2CBA02AC",
    x"2CB9EB6D",
    x"2CB9D431",
    x"2CB9BCF8",
    x"2CB9A5C2",
    x"2CB98E8F",
    x"2CB9775F",
    x"2CB96031",
    x"2CB94907",
    x"2CB931DF",
    x"2CB91ABA",
    x"2CB90398",
    x"2CB8EC79",
    x"2CB8D55D",
    x"2CB8BE44",
    x"2CB8A72D",
    x"2CB8901A",
    x"2CB87909",
    x"2CB861FC",
    x"2CB84AF1",
    x"2CB833E9",
    x"2CB81CE4",
    x"2CB805E2",
    x"2CB7EEE3",
    x"2CB7D7E6",
    x"2CB7C0ED",
    x"2CB7A9F6",
    x"2CB79302",
    x"2CB77C11",
    x"2CB76523",
    x"2CB74E38",
    x"2CB7374F",
    x"2CB7206A",
    x"2CB70987",
    x"2CB6F2A8",
    x"2CB6DBCB",
    x"2CB6C4F1",
    x"2CB6AE19",
    x"2CB69745",
    x"2CB68074",
    x"2CB669A5",
    x"2CB652D9",
    x"2CB63C10",
    x"2CB6254A",
    x"2CB60E87",
    x"2CB5F7C7",
    x"2CB5E109",
    x"2CB5CA4E",
    x"2CB5B396",
    x"2CB59CE1",
    x"2CB5862F",
    x"2CB56F80",
    x"2CB558D3",
    x"2CB5422A",
    x"2CB52B83",
    x"2CB514DF",
    x"2CB4FE3E",
    x"2CB4E79F",
    x"2CB4D104",
    x"2CB4BA6B",
    x"2CB4A3D5",
    x"2CB48D42",
    x"2CB476B2",
    x"2CB46024",
    x"2CB4499A",
    x"2CB43312",
    x"2CB41C8D",
    x"2CB4060B",
    x"2CB3EF8B",
    x"2CB3D90F",
    x"2CB3C295",
    x"2CB3AC1E",
    x"2CB395AA",
    x"2CB37F39",
    x"2CB368CA",
    x"2CB3525F",
    x"2CB33BF6",
    x"2CB32590",
    x"2CB30F2C",
    x"2CB2F8CC",
    x"2CB2E26E",
    x"2CB2CC13",
    x"2CB2B5BB",
    x"2CB29F66",
    x"2CB28913",
    x"2CB272C4",
    x"2CB25C77",
    x"2CB2462C",
    x"2CB22FE5",
    x"2CB219A0",
    x"2CB2035F",
    x"2CB1ED20",
    x"2CB1D6E3",
    x"2CB1C0AA",
    x"2CB1AA73",
    x"2CB1943F",
    x"2CB17E0E",
    x"2CB167E0",
    x"2CB151B4",
    x"2CB13B8B",
    x"2CB12565",
    x"2CB10F42",
    x"2CB0F922",
    x"2CB0E304",
    x"2CB0CCE9",
    x"2CB0B6D1",
    x"2CB0A0BB",
    x"2CB08AA8",
    x"2CB07498",
    x"2CB05E8B",
    x"2CB04881",
    x"2CB03279",
    x"2CB01C74",
    x"2CB00672",
    x"2CAFF073",
    x"2CAFDA76",
    x"2CAFC47C",
    x"2CAFAE85",
    x"2CAF9890",
    x"2CAF829F",
    x"2CAF6CB0",
    x"2CAF56C3",
    x"2CAF40DA",
    x"2CAF2AF3",
    x"2CAF150F",
    x"2CAEFF2E",
    x"2CAEE94F",
    x"2CAED374",
    x"2CAEBD9B",
    x"2CAEA7C4",
    x"2CAE91F1",
    x"2CAE7C20",
    x"2CAE6652",
    x"2CAE5086",
    x"2CAE3ABD",
    x"2CAE24F7",
    x"2CAE0F34",
    x"2CADF974",
    x"2CADE3B6",
    x"2CADCDFB",
    x"2CADB842",
    x"2CADA28D",
    x"2CAD8CDA",
    x"2CAD7729",
    x"2CAD617C",
    x"2CAD4BD1",
    x"2CAD3629",
    x"2CAD2084",
    x"2CAD0AE1",
    x"2CACF541",
    x"2CACDFA3",
    x"2CACCA09",
    x"2CACB471",
    x"2CAC9EDC",
    x"2CAC8949",
    x"2CAC73B9",
    x"2CAC5E2C",
    x"2CAC48A2",
    x"2CAC331A",
    x"2CAC1D95",
    x"2CAC0813",
    x"2CABF293",
    x"2CABDD16",
    x"2CABC79C",
    x"2CABB224",
    x"2CAB9CAF",
    x"2CAB873D",
    x"2CAB71CE",
    x"2CAB5C61",
    x"2CAB46F6",
    x"2CAB318F",
    x"2CAB1C2A",
    x"2CAB06C8",
    x"2CAAF168",
    x"2CAADC0B",
    x"2CAAC6B1",
    x"2CAAB15A",
    x"2CAA9C05",
    x"2CAA86B3",
    x"2CAA7163",
    x"2CAA5C16",
    x"2CAA46CC",
    x"2CAA3185",
    x"2CAA1C40",
    x"2CAA06FE",
    x"2CA9F1BE",
    x"2CA9DC81",
    x"2CA9C747",
    x"2CA9B20F",
    x"2CA99CDB",
    x"2CA987A8",
    x"2CA97279",
    x"2CA95D4C",
    x"2CA94821",
    x"2CA932FA",
    x"2CA91DD5",
    x"2CA908B2",
    x"2CA8F392",
    x"2CA8DE75",
    x"2CA8C95B",
    x"2CA8B443",
    x"2CA89F2E",
    x"2CA88A1B",
    x"2CA8750B",
    x"2CA85FFE",
    x"2CA84AF3",
    x"2CA835EB",
    x"2CA820E6",
    x"2CA80BE3",
    x"2CA7F6E3",
    x"2CA7E1E5",
    x"2CA7CCEA",
    x"2CA7B7F2",
    x"2CA7A2FC",
    x"2CA78E09",
    x"2CA77919",
    x"2CA7642B",
    x"2CA74F40",
    x"2CA73A57",
    x"2CA72571",
    x"2CA7108E",
    x"2CA6FBAD",
    x"2CA6E6CF",
    x"2CA6D1F3",
    x"2CA6BD1A",
    x"2CA6A844",
    x"2CA69370",
    x"2CA67E9F",
    x"2CA669D1",
    x"2CA65505",
    x"2CA6403B",
    x"2CA62B75",
    x"2CA616B0",
    x"2CA601EF",
    x"2CA5ED30",
    x"2CA5D874",
    x"2CA5C3BA",
    x"2CA5AF03",
    x"2CA59A4E",
    x"2CA5859C",
    x"2CA570ED",
    x"2CA55C40",
    x"2CA54796",
    x"2CA532EE",
    x"2CA51E49",
    x"2CA509A6",
    x"2CA4F507",
    x"2CA4E069",
    x"2CA4CBCE",
    x"2CA4B736",
    x"2CA4A2A1",
    x"2CA48E0E",
    x"2CA4797D",
    x"2CA464EF",
    x"2CA45064",
    x"2CA43BDB",
    x"2CA42755",
    x"2CA412D1",
    x"2CA3FE50",
    x"2CA3E9D2",
    x"2CA3D556",
    x"2CA3C0DC",
    x"2CA3AC66",
    x"2CA397F1",
    x"2CA38380",
    x"2CA36F10",
    x"2CA35AA4",
    x"2CA3463A",
    x"2CA331D2",
    x"2CA31D6D",
    x"2CA3090B",
    x"2CA2F4AB",
    x"2CA2E04E",
    x"2CA2CBF3",
    x"2CA2B79B",
    x"2CA2A345",
    x"2CA28EF2",
    x"2CA27AA1",
    x"2CA26653",
    x"2CA25208",
    x"2CA23DBF",
    x"2CA22978",
    x"2CA21534",
    x"2CA200F3",
    x"2CA1ECB4",
    x"2CA1D878",
    x"2CA1C43E",
    x"2CA1B007",
    x"2CA19BD2",
    x"2CA187A0",
    x"2CA17370",
    x"2CA15F43",
    x"2CA14B18",
    x"2CA136F0",
    x"2CA122CB",
    x"2CA10EA7",
    x"2CA0FA87",
    x"2CA0E669",
    x"2CA0D24D",
    x"2CA0BE34",
    x"2CA0AA1E",
    x"2CA0960A",
    x"2CA081F8",
    x"2CA06DE9",
    x"2CA059DD",
    x"2CA045D3",
    x"2CA031CB",
    x"2CA01DC6",
    x"2CA009C4",
    x"2C9FF5C4",
    x"2C9FE1C6",
    x"2C9FCDCB",
    x"2C9FB9D3",
    x"2C9FA5DD",
    x"2C9F91E9",
    x"2C9F7DF8",
    x"2C9F6A0A",
    x"2C9F561E",
    x"2C9F4234",
    x"2C9F2E4D",
    x"2C9F1A69",
    x"2C9F0687",
    x"2C9EF2A7",
    x"2C9EDECA",
    x"2C9ECAF0",
    x"2C9EB717",
    x"2C9EA342",
    x"2C9E8F6F",
    x"2C9E7B9E",
    x"2C9E67D0",
    x"2C9E5404",
    x"2C9E403B",
    x"2C9E2C74",
    x"2C9E18B0",
    x"2C9E04EE",
    x"2C9DF12E",
    x"2C9DDD71",
    x"2C9DC9B7",
    x"2C9DB5FF",
    x"2C9DA249",
    x"2C9D8E96",
    x"2C9D7AE6",
    x"2C9D6738",
    x"2C9D538C",
    x"2C9D3FE3",
    x"2C9D2C3C",
    x"2C9D1898",
    x"2C9D04F6",
    x"2C9CF157",
    x"2C9CDDBA",
    x"2C9CCA1F",
    x"2C9CB687",
    x"2C9CA2F1",
    x"2C9C8F5E",
    x"2C9C7BCE",
    x"2C9C683F",
    x"2C9C54B4",
    x"2C9C412A",
    x"2C9C2DA3",
    x"2C9C1A1F",
    x"2C9C069D",
    x"2C9BF31D",
    x"2C9BDFA0",
    x"2C9BCC25",
    x"2C9BB8AD",
    x"2C9BA537",
    x"2C9B91C4",
    x"2C9B7E53",
    x"2C9B6AE4",
    x"2C9B5778",
    x"2C9B440E",
    x"2C9B30A7",
    x"2C9B1D42",
    x"2C9B09E0",
    x"2C9AF680",
    x"2C9AE322",
    x"2C9ACFC7",
    x"2C9ABC6E",
    x"2C9AA918",
    x"2C9A95C4",
    x"2C9A8272",
    x"2C9A6F23",
    x"2C9A5BD6",
    x"2C9A488C",
    x"2C9A3544",
    x"2C9A21FF",
    x"2C9A0EBC",
    x"2C99FB7B",
    x"2C99E83D",
    x"2C99D501",
    x"2C99C1C8",
    x"2C99AE91",
    x"2C999B5C",
    x"2C99882A",
    x"2C9974FA",
    x"2C9961CD",
    x"2C994EA2",
    x"2C993B79",
    x"2C992853",
    x"2C99152F",
    x"2C99020D",
    x"2C98EEEE",
    x"2C98DBD2",
    x"2C98C8B7",
    x"2C98B59F",
    x"2C98A28A",
    x"2C988F77",
    x"2C987C66",
    x"2C986958",
    x"2C98564C",
    x"2C984342",
    x"2C98303B",
    x"2C981D36",
    x"2C980A34",
    x"2C97F734",
    x"2C97E436",
    x"2C97D13A",
    x"2C97BE41",
    x"2C97AB4B",
    x"2C979857",
    x"2C978565",
    x"2C977275",
    x"2C975F88",
    x"2C974C9D",
    x"2C9739B5",
    x"2C9726CF",
    x"2C9713EB",
    x"2C97010A",
    x"2C96EE2B",
    x"2C96DB4E",
    x"2C96C874",
    x"2C96B59C",
    x"2C96A2C7",
    x"2C968FF4",
    x"2C967D23",
    x"2C966A54",
    x"2C965788",
    x"2C9644BF",
    x"2C9631F7",
    x"2C961F32",
    x"2C960C6F",
    x"2C95F9AF",
    x"2C95E6F1",
    x"2C95D435",
    x"2C95C17C",
    x"2C95AEC5",
    x"2C959C10",
    x"2C95895E",
    x"2C9576AE",
    x"2C956400",
    x"2C955155",
    x"2C953EAC",
    x"2C952C05",
    x"2C951961",
    x"2C9506BF",
    x"2C94F41F",
    x"2C94E182",
    x"2C94CEE7",
    x"2C94BC4E",
    x"2C94A9B8",
    x"2C949724",
    x"2C948492",
    x"2C947202",
    x"2C945F75",
    x"2C944CEB",
    x"2C943A62",
    x"2C9427DC",
    x"2C941558",
    x"2C9402D7",
    x"2C93F057",
    x"2C93DDDB",
    x"2C93CB60",
    x"2C93B8E8",
    x"2C93A672",
    x"2C9393FE",
    x"2C93818D",
    x"2C936F1E",
    x"2C935CB1",
    x"2C934A47",
    x"2C9337DE",
    x"2C932579",
    x"2C931315",
    x"2C9300B4",
    x"2C92EE55",
    x"2C92DBF8",
    x"2C92C99E",
    x"2C92B746",
    x"2C92A4F0",
    x"2C92929D",
    x"2C92804B",
    x"2C926DFD",
    x"2C925BB0",
    x"2C924966",
    x"2C92371E",
    x"2C9224D8",
    x"2C921294",
    x"2C920053",
    x"2C91EE14",
    x"2C91DBD8",
    x"2C91C99D",
    x"2C91B765",
    x"2C91A52F",
    x"2C9192FC",
    x"2C9180CB",
    x"2C916E9C",
    x"2C915C6F",
    x"2C914A45",
    x"2C91381C",
    x"2C9125F7",
    x"2C9113D3",
    x"2C9101B2",
    x"2C90EF93",
    x"2C90DD76",
    x"2C90CB5B",
    x"2C90B943",
    x"2C90A72D",
    x"2C909519",
    x"2C908308",
    x"2C9070F8",
    x"2C905EEB",
    x"2C904CE1",
    x"2C903AD8",
    x"2C9028D2",
    x"2C9016CE",
    x"2C9004CC",
    x"2C8FF2CD",
    x"2C8FE0D0",
    x"2C8FCED5",
    x"2C8FBCDC",
    x"2C8FAAE5",
    x"2C8F98F1",
    x"2C8F86FF",
    x"2C8F750F",
    x"2C8F6322",
    x"2C8F5137",
    x"2C8F3F4E",
    x"2C8F2D67",
    x"2C8F1B82",
    x"2C8F09A0",
    x"2C8EF7C0",
    x"2C8EE5E2",
    x"2C8ED406",
    x"2C8EC22D",
    x"2C8EB056",
    x"2C8E9E81",
    x"2C8E8CAE",
    x"2C8E7ADE",
    x"2C8E690F",
    x"2C8E5743",
    x"2C8E457A",
    x"2C8E33B2",
    x"2C8E21ED",
    x"2C8E102A",
    x"2C8DFE69",
    x"2C8DECAA",
    x"2C8DDAED",
    x"2C8DC933",
    x"2C8DB77B",
    x"2C8DA5C5",
    x"2C8D9412",
    x"2C8D8260",
    x"2C8D70B1",
    x"2C8D5F04",
    x"2C8D4D59",
    x"2C8D3BB1",
    x"2C8D2A0A",
    x"2C8D1866",
    x"2C8D06C4",
    x"2C8CF525",
    x"2C8CE387",
    x"2C8CD1EC",
    x"2C8CC053",
    x"2C8CAEBC",
    x"2C8C9D27",
    x"2C8C8B94",
    x"2C8C7A04",
    x"2C8C6876",
    x"2C8C56EA",
    x"2C8C4560",
    x"2C8C33D9",
    x"2C8C2253",
    x"2C8C10D0",
    x"2C8BFF4F",
    x"2C8BEDD0",
    x"2C8BDC53",
    x"2C8BCAD9",
    x"2C8BB961",
    x"2C8BA7EB",
    x"2C8B9677",
    x"2C8B8505",
    x"2C8B7396",
    x"2C8B6228",
    x"2C8B50BD",
    x"2C8B3F54",
    x"2C8B2DED",
    x"2C8B1C89",
    x"2C8B0B26",
    x"2C8AF9C6",
    x"2C8AE868",
    x"2C8AD70C",
    x"2C8AC5B2",
    x"2C8AB45A",
    x"2C8AA305",
    x"2C8A91B1",
    x"2C8A8060",
    x"2C8A6F11",
    x"2C8A5DC5",
    x"2C8A4C7A",
    x"2C8A3B31",
    x"2C8A29EB",
    x"2C8A18A7",
    x"2C8A0765",
    x"2C89F625",
    x"2C89E4E7",
    x"2C89D3AC",
    x"2C89C272",
    x"2C89B13B",
    x"2C89A006",
    x"2C898ED3",
    x"2C897DA2",
    x"2C896C74",
    x"2C895B47",
    x"2C894A1D",
    x"2C8938F5",
    x"2C8927CF",
    x"2C8916AB",
    x"2C890589",
    x"2C88F46A",
    x"2C88E34C",
    x"2C88D231",
    x"2C88C117",
    x"2C88B000",
    x"2C889EEB",
    x"2C888DD9",
    x"2C887CC8",
    x"2C886BB9",
    x"2C885AAD",
    x"2C8849A3",
    x"2C88389B",
    x"2C882795",
    x"2C881691",
    x"2C88058F",
    x"2C87F48F",
    x"2C87E392",
    x"2C87D296",
    x"2C87C19D",
    x"2C87B0A6",
    x"2C879FB1",
    x"2C878EBE",
    x"2C877DCD",
    x"2C876CDF",
    x"2C875BF2",
    x"2C874B08",
    x"2C873A1F",
    x"2C872939",
    x"2C871855",
    x"2C870773",
    x"2C86F693",
    x"2C86E5B5",
    x"2C86D4DA",
    x"2C86C400",
    x"2C86B329",
    x"2C86A253",
    x"2C869180",
    x"2C8680AF",
    x"2C866FE0",
    x"2C865F13",
    x"2C864E48",
    x"2C863D80",
    x"2C862CB9",
    x"2C861BF4",
    x"2C860B32",
    x"2C85FA72",
    x"2C85E9B3",
    x"2C85D8F7",
    x"2C85C83D",
    x"2C85B785",
    x"2C85A6CF",
    x"2C85961B",
    x"2C85856A",
    x"2C8574BA",
    x"2C85640C",
    x"2C855361",
    x"2C8542B8",
    x"2C853210",
    x"2C85216B",
    x"2C8510C8",
    x"2C850027",
    x"2C84EF88",
    x"2C84DEEB",
    x"2C84CE50",
    x"2C84BDB7",
    x"2C84AD21",
    x"2C849C8C",
    x"2C848BFA",
    x"2C847B69",
    x"2C846ADB",
    x"2C845A4E",
    x"2C8449C4",
    x"2C84393C",
    x"2C8428B6",
    x"2C841832",
    x"2C8407B0",
    x"2C83F730",
    x"2C83E6B2",
    x"2C83D636",
    x"2C83C5BD",
    x"2C83B545",
    x"2C83A4CF",
    x"2C83945C",
    x"2C8383EA",
    x"2C83737B",
    x"2C83630D",
    x"2C8352A2",
    x"2C834239",
    x"2C8331D1",
    x"2C83216C",
    x"2C831109",
    x"2C8300A8",
    x"2C82F049",
    x"2C82DFEC",
    x"2C82CF91",
    x"2C82BF38",
    x"2C82AEE1",
    x"2C829E8C",
    x"2C828E39",
    x"2C827DE9",
    x"2C826D9A",
    x"2C825D4D",
    x"2C824D03",
    x"2C823CBA",
    x"2C822C73",
    x"2C821C2F",
    x"2C820BEC",
    x"2C81FBAC",
    x"2C81EB6D",
    x"2C81DB31",
    x"2C81CAF7",
    x"2C81BABE",
    x"2C81AA88",
    x"2C819A54",
    x"2C818A21",
    x"2C8179F1",
    x"2C8169C3",
    x"2C815997",
    x"2C81496C",
    x"2C813944",
    x"2C81291E",
    x"2C8118FA",
    x"2C8108D8",
    x"2C80F8B8",
    x"2C80E89A",
    x"2C80D87E",
    x"2C80C864",
    x"2C80B84C",
    x"2C80A836",
    x"2C809822",
    x"2C808810",
    x"2C807800",
    x"2C8067F2",
    x"2C8057E6",
    x"2C8047DC",
    x"2C8037D4",
    x"2C8027CE",
    x"2C8017CA",
    x"2C8007C8",
    x"2C7FEF8F",
    x"2C7FCF93",
    x"2C7FAF9B",
    x"2C7F8FA7",
    x"2C7F6FB8",
    x"2C7F4FCC",
    x"2C7F2FE4",
    x"2C7F1000",
    x"2C7EF020",
    x"2C7ED044",
    x"2C7EB06B",
    x"2C7E9097",
    x"2C7E70C7",
    x"2C7E50FB",
    x"2C7E3133",
    x"2C7E116F",
    x"2C7DF1AF",
    x"2C7DD1F3",
    x"2C7DB23A",
    x"2C7D9286",
    x"2C7D72D6",
    x"2C7D5329",
    x"2C7D3381",
    x"2C7D13DC",
    x"2C7CF43C",
    x"2C7CD49F",
    x"2C7CB507",
    x"2C7C9572",
    x"2C7C75E1",
    x"2C7C5655",
    x"2C7C36CC",
    x"2C7C1747",
    x"2C7BF7C6",
    x"2C7BD849",
    x"2C7BB8D0",
    x"2C7B995B",
    x"2C7B79EA",
    x"2C7B5A7C",
    x"2C7B3B13",
    x"2C7B1BAD",
    x"2C7AFC4C",
    x"2C7ADCEE",
    x"2C7ABD95",
    x"2C7A9E3F",
    x"2C7A7EED",
    x"2C7A5F9F",
    x"2C7A4055",
    x"2C7A210F",
    x"2C7A01CD",
    x"2C79E28F",
    x"2C79C354",
    x"2C79A41E",
    x"2C7984EB",
    x"2C7965BD",
    x"2C794692",
    x"2C79276B",
    x"2C790848",
    x"2C78E929",
    x"2C78CA0E",
    x"2C78AAF6",
    x"2C788BE3",
    x"2C786CD3",
    x"2C784DC8",
    x"2C782EC0",
    x"2C780FBC",
    x"2C77F0BC",
    x"2C77D1C0",
    x"2C77B2C8",
    x"2C7793D3",
    x"2C7774E3",
    x"2C7755F6",
    x"2C77370D",
    x"2C771828",
    x"2C76F947",
    x"2C76DA6A",
    x"2C76BB91",
    x"2C769CBB",
    x"2C767DE9",
    x"2C765F1C",
    x"2C764052",
    x"2C76218B",
    x"2C7602C9",
    x"2C75E40B",
    x"2C75C550",
    x"2C75A699",
    x"2C7587E7",
    x"2C756937",
    x"2C754A8C",
    x"2C752BE5",
    x"2C750D41",
    x"2C74EEA2",
    x"2C74D006",
    x"2C74B16E",
    x"2C7492D9",
    x"2C747449",
    x"2C7455BC",
    x"2C743733",
    x"2C7418AE",
    x"2C73FA2D",
    x"2C73DBB0",
    x"2C73BD36",
    x"2C739EC1",
    x"2C73804F",
    x"2C7361E0",
    x"2C734376",
    x"2C732510",
    x"2C7306AD",
    x"2C72E84E",
    x"2C72C9F3",
    x"2C72AB9B",
    x"2C728D48",
    x"2C726EF8",
    x"2C7250AC",
    x"2C723264",
    x"2C721420",
    x"2C71F5DF",
    x"2C71D7A2",
    x"2C71B969",
    x"2C719B34",
    x"2C717D02",
    x"2C715ED4",
    x"2C7140AB",
    x"2C712284",
    x"2C710462",
    x"2C70E643",
    x"2C70C828",
    x"2C70AA11",
    x"2C708BFE",
    x"2C706DEE",
    x"2C704FE2",
    x"2C7031DA",
    x"2C7013D6",
    x"2C6FF5D5",
    x"2C6FD7D8",
    x"2C6FB9DF",
    x"2C6F9BEA",
    x"2C6F7DF8",
    x"2C6F600A",
    x"2C6F4220",
    x"2C6F243A",
    x"2C6F0657",
    x"2C6EE878",
    x"2C6ECA9D",
    x"2C6EACC6",
    x"2C6E8EF2",
    x"2C6E7122",
    x"2C6E5356",
    x"2C6E358D",
    x"2C6E17C8",
    x"2C6DFA07",
    x"2C6DDC4A",
    x"2C6DBE90",
    x"2C6DA0DA",
    x"2C6D8328",
    x"2C6D6579",
    x"2C6D47CE",
    x"2C6D2A27",
    x"2C6D0C84",
    x"2C6CEEE4",
    x"2C6CD148",
    x"2C6CB3B0",
    x"2C6C961B",
    x"2C6C788A",
    x"2C6C5AFD",
    x"2C6C3D74",
    x"2C6C1FEE",
    x"2C6C026C",
    x"2C6BE4ED",
    x"2C6BC772",
    x"2C6BA9FB",
    x"2C6B8C88",
    x"2C6B6F18",
    x"2C6B51AC",
    x"2C6B3444",
    x"2C6B16DF",
    x"2C6AF97E",
    x"2C6ADC21",
    x"2C6ABEC7",
    x"2C6AA171",
    x"2C6A841F",
    x"2C6A66D0",
    x"2C6A4985",
    x"2C6A2C3E",
    x"2C6A0EFA",
    x"2C69F1BA",
    x"2C69D47D",
    x"2C69B745",
    x"2C699A10",
    x"2C697CDE",
    x"2C695FB0",
    x"2C694286",
    x"2C692560",
    x"2C69083D",
    x"2C68EB1E",
    x"2C68CE02",
    x"2C68B0EA",
    x"2C6893D6",
    x"2C6876C5",
    x"2C6859B8",
    x"2C683CAF",
    x"2C681FA9",
    x"2C6802A7",
    x"2C67E5A8",
    x"2C67C8AE",
    x"2C67ABB6",
    x"2C678EC3",
    x"2C6771D3",
    x"2C6754E6",
    x"2C6737FD",
    x"2C671B18",
    x"2C66FE37",
    x"2C66E159",
    x"2C66C47E",
    x"2C66A7A7",
    x"2C668AD4",
    x"2C666E05",
    x"2C665139",
    x"2C663470",
    x"2C6617AC",
    x"2C65FAEB",
    x"2C65DE2D",
    x"2C65C173",
    x"2C65A4BD",
    x"2C65880A",
    x"2C656B5B",
    x"2C654EAF",
    x"2C653207",
    x"2C651562",
    x"2C64F8C2",
    x"2C64DC24",
    x"2C64BF8B",
    x"2C64A2F4",
    x"2C648662",
    x"2C6469D3",
    x"2C644D47",
    x"2C6430BF",
    x"2C64143B",
    x"2C63F7BA",
    x"2C63DB3D",
    x"2C63BEC4",
    x"2C63A24E",
    x"2C6385DB",
    x"2C63696C",
    x"2C634D01",
    x"2C633099",
    x"2C631435",
    x"2C62F7D4",
    x"2C62DB77",
    x"2C62BF1D",
    x"2C62A2C7",
    x"2C628674",
    x"2C626A25",
    x"2C624DDA",
    x"2C623192",
    x"2C62154D",
    x"2C61F90C",
    x"2C61DCCF",
    x"2C61C095",
    x"2C61A45F",
    x"2C61882C",
    x"2C616BFD",
    x"2C614FD1",
    x"2C6133A9",
    x"2C611784",
    x"2C60FB63",
    x"2C60DF45",
    x"2C60C32B",
    x"2C60A715",
    x"2C608B01",
    x"2C606EF2",
    x"2C6052E6",
    x"2C6036DD",
    x"2C601AD8",
    x"2C5FFED6",
    x"2C5FE2D8",
    x"2C5FC6DE",
    x"2C5FAAE7",
    x"2C5F8EF3",
    x"2C5F7303",
    x"2C5F5716",
    x"2C5F3B2D",
    x"2C5F1F47",
    x"2C5F0365",
    x"2C5EE786",
    x"2C5ECBAB",
    x"2C5EAFD4",
    x"2C5E93FF",
    x"2C5E782F",
    x"2C5E5C61",
    x"2C5E4097",
    x"2C5E24D1",
    x"2C5E090E",
    x"2C5DED4F",
    x"2C5DD193",
    x"2C5DB5DA",
    x"2C5D9A25",
    x"2C5D7E74",
    x"2C5D62C6",
    x"2C5D471B",
    x"2C5D2B74",
    x"2C5D0FD0",
    x"2C5CF430",
    x"2C5CD893",
    x"2C5CBCFA",
    x"2C5CA164",
    x"2C5C85D2",
    x"2C5C6A43",
    x"2C5C4EB7",
    x"2C5C332F",
    x"2C5C17AA",
    x"2C5BFC29",
    x"2C5BE0AB",
    x"2C5BC531",
    x"2C5BA9BA",
    x"2C5B8E46",
    x"2C5B72D6",
    x"2C5B576A",
    x"2C5B3C01",
    x"2C5B209B",
    x"2C5B0538",
    x"2C5AE9D9",
    x"2C5ACE7E",
    x"2C5AB326",
    x"2C5A97D1",
    x"2C5A7C80",
    x"2C5A6132",
    x"2C5A45E8",
    x"2C5A2AA1",
    x"2C5A0F5D",
    x"2C59F41D",
    x"2C59D8E0",
    x"2C59BDA6",
    x"2C59A270",
    x"2C59873E",
    x"2C596C0F",
    x"2C5950E3",
    x"2C5935BA",
    x"2C591A95",
    x"2C58FF74",
    x"2C58E456",
    x"2C58C93B",
    x"2C58AE23",
    x"2C58930F",
    x"2C5877FE",
    x"2C585CF1",
    x"2C5841E7",
    x"2C5826E1",
    x"2C580BDE",
    x"2C57F0DE",
    x"2C57D5E1",
    x"2C57BAE8",
    x"2C579FF3",
    x"2C578500",
    x"2C576A11",
    x"2C574F26",
    x"2C57343E",
    x"2C571959",
    x"2C56FE77",
    x"2C56E399",
    x"2C56C8BE",
    x"2C56ADE7",
    x"2C569313",
    x"2C567842",
    x"2C565D75",
    x"2C5642AB",
    x"2C5627E4",
    x"2C560D21",
    x"2C55F261",
    x"2C55D7A4",
    x"2C55BCEB",
    x"2C55A235",
    x"2C558782",
    x"2C556CD3",
    x"2C555227",
    x"2C55377F",
    x"2C551CD9",
    x"2C550237",
    x"2C54E799",
    x"2C54CCFD",
    x"2C54B265",
    x"2C5497D1",
    x"2C547D3F",
    x"2C5462B2",
    x"2C544827",
    x"2C542D9F",
    x"2C54131B",
    x"2C53F89B",
    x"2C53DE1D",
    x"2C53C3A3",
    x"2C53A92C",
    x"2C538EB9",
    x"2C537449",
    x"2C5359DC",
    x"2C533F72",
    x"2C53250C",
    x"2C530AA9",
    x"2C52F049",
    x"2C52D5ED",
    x"2C52BB94",
    x"2C52A13E",
    x"2C5286EB",
    x"2C526C9C",
    x"2C525250",
    x"2C523808",
    x"2C521DC2",
    x"2C520380",
    x"2C51E941",
    x"2C51CF06",
    x"2C51B4CE",
    x"2C519A99",
    x"2C518067",
    x"2C516639",
    x"2C514C0D",
    x"2C5131E6",
    x"2C5117C1",
    x"2C50FDA0",
    x"2C50E382",
    x"2C50C967",
    x"2C50AF4F",
    x"2C50953B",
    x"2C507B2A",
    x"2C50611C",
    x"2C504712",
    x"2C502D0A",
    x"2C501306",
    x"2C4FF906",
    x"2C4FDF08",
    x"2C4FC50E",
    x"2C4FAB17",
    x"2C4F9123",
    x"2C4F7733",
    x"2C4F5D45",
    x"2C4F435B",
    x"2C4F2974",
    x"2C4F0F91",
    x"2C4EF5B1",
    x"2C4EDBD3",
    x"2C4EC1FA",
    x"2C4EA823",
    x"2C4E8E50",
    x"2C4E747F",
    x"2C4E5AB2",
    x"2C4E40E9",
    x"2C4E2722",
    x"2C4E0D5F",
    x"2C4DF39F",
    x"2C4DD9E2",
    x"2C4DC028",
    x"2C4DA672",
    x"2C4D8CBF",
    x"2C4D730F",
    x"2C4D5962",
    x"2C4D3FB8",
    x"2C4D2612",
    x"2C4D0C6F",
    x"2C4CF2CF",
    x"2C4CD932",
    x"2C4CBF99",
    x"2C4CA602",
    x"2C4C8C6F",
    x"2C4C72DF",
    x"2C4C5952",
    x"2C4C3FC9",
    x"2C4C2643",
    x"2C4C0CBF",
    x"2C4BF33F",
    x"2C4BD9C3",
    x"2C4BC049",
    x"2C4BA6D2",
    x"2C4B8D5F",
    x"2C4B73EF",
    x"2C4B5A82",
    x"2C4B4118",
    x"2C4B27B2",
    x"2C4B0E4F",
    x"2C4AF4EE",
    x"2C4ADB91",
    x"2C4AC237",
    x"2C4AA8E1",
    x"2C4A8F8D",
    x"2C4A763D",
    x"2C4A5CF0",
    x"2C4A43A6",
    x"2C4A2A5F",
    x"2C4A111B",
    x"2C49F7DB",
    x"2C49DE9D",
    x"2C49C563",
    x"2C49AC2C",
    x"2C4992F8",
    x"2C4979C7",
    x"2C496099",
    x"2C49476F",
    x"2C492E48",
    x"2C491523",
    x"2C48FC02",
    x"2C48E2E4",
    x"2C48C9C9",
    x"2C48B0B2",
    x"2C48979D",
    x"2C487E8C",
    x"2C48657E",
    x"2C484C73",
    x"2C48336B",
    x"2C481A66",
    x"2C480164",
    x"2C47E865",
    x"2C47CF6A",
    x"2C47B672",
    x"2C479D7C",
    x"2C47848A",
    x"2C476B9B",
    x"2C4752AF",
    x"2C4739C6",
    x"2C4720E1",
    x"2C4707FE",
    x"2C46EF1F",
    x"2C46D642",
    x"2C46BD69",
    x"2C46A493",
    x"2C468BC0",
    x"2C4672F0",
    x"2C465A23",
    x"2C46415A",
    x"2C462893",
    x"2C460FCF",
    x"2C45F70F",
    x"2C45DE52",
    x"2C45C597",
    x"2C45ACE0",
    x"2C45942C",
    x"2C457B7B",
    x"2C4562CD",
    x"2C454A23",
    x"2C45317B",
    x"2C4518D6",
    x"2C450035",
    x"2C44E796",
    x"2C44CEFB",
    x"2C44B662",
    x"2C449DCD",
    x"2C44853B",
    x"2C446CAC",
    x"2C445420",
    x"2C443B97",
    x"2C442311",
    x"2C440A8E",
    x"2C43F20E",
    x"2C43D992",
    x"2C43C118",
    x"2C43A8A1",
    x"2C43902E",
    x"2C4377BD",
    x"2C435F50",
    x"2C4346E5",
    x"2C432E7E",
    x"2C43161A",
    x"2C42FDB9",
    x"2C42E55A",
    x"2C42CCFF",
    x"2C42B4A7",
    x"2C429C52",
    x"2C428400",
    x"2C426BB1",
    x"2C425365",
    x"2C423B1C",
    x"2C4222D6",
    x"2C420A93",
    x"2C41F254",
    x"2C41DA17",
    x"2C41C1DD",
    x"2C41A9A6",
    x"2C419173",
    x"2C417942",
    x"2C416114",
    x"2C4148EA",
    x"2C4130C2",
    x"2C41189E",
    x"2C41007C",
    x"2C40E85D",
    x"2C40D042",
    x"2C40B829",
    x"2C40A014",
    x"2C408801",
    x"2C406FF2",
    x"2C4057E5",
    x"2C403FDC",
    x"2C4027D5",
    x"2C400FD2",
    x"2C3FF7D1",
    x"2C3FDFD4",
    x"2C3FC7DA",
    x"2C3FAFE2",
    x"2C3F97EE",
    x"2C3F7FFC",
    x"2C3F680E",
    x"2C3F5022",
    x"2C3F383A",
    x"2C3F2054",
    x"2C3F0871",
    x"2C3EF092",
    x"2C3ED8B5",
    x"2C3EC0DC",
    x"2C3EA905",
    x"2C3E9131",
    x"2C3E7961",
    x"2C3E6193",
    x"2C3E49C8",
    x"2C3E3201",
    x"2C3E1A3C",
    x"2C3E027A",
    x"2C3DEABB",
    x"2C3DD2FF",
    x"2C3DBB47",
    x"2C3DA391",
    x"2C3D8BDE",
    x"2C3D742E",
    x"2C3D5C81",
    x"2C3D44D6",
    x"2C3D2D2F",
    x"2C3D158B",
    x"2C3CFDEA",
    x"2C3CE64C",
    x"2C3CCEB0",
    x"2C3CB718",
    x"2C3C9F83",
    x"2C3C87F0",
    x"2C3C7061",
    x"2C3C58D4",
    x"2C3C414A",
    x"2C3C29C4",
    x"2C3C1240",
    x"2C3BFABF",
    x"2C3BE341",
    x"2C3BCBC6",
    x"2C3BB44E",
    x"2C3B9CD9",
    x"2C3B8567",
    x"2C3B6DF8",
    x"2C3B568C",
    x"2C3B3F22",
    x"2C3B27BC",
    x"2C3B1058",
    x"2C3AF8F8",
    x"2C3AE19A",
    x"2C3ACA3F",
    x"2C3AB2E8",
    x"2C3A9B93",
    x"2C3A8441",
    x"2C3A6CF2",
    x"2C3A55A5",
    x"2C3A3E5C",
    x"2C3A2716",
    x"2C3A0FD2",
    x"2C39F892",
    x"2C39E154",
    x"2C39CA1A",
    x"2C39B2E2",
    x"2C399BAD",
    x"2C39847B",
    x"2C396D4C",
    x"2C39561F",
    x"2C393EF6",
    x"2C3927D0",
    x"2C3910AC",
    x"2C38F98C",
    x"2C38E26E",
    x"2C38CB53",
    x"2C38B43B",
    x"2C389D26",
    x"2C388614",
    x"2C386F04",
    x"2C3857F8",
    x"2C3840EE",
    x"2C3829E8",
    x"2C3812E4",
    x"2C37FBE3",
    x"2C37E4E5",
    x"2C37CDEA",
    x"2C37B6F1",
    x"2C379FFC",
    x"2C378909",
    x"2C37721A",
    x"2C375B2D",
    x"2C374443",
    x"2C372D5C",
    x"2C371678",
    x"2C36FF96",
    x"2C36E8B8",
    x"2C36D1DC",
    x"2C36BB03",
    x"2C36A42D",
    x"2C368D5A",
    x"2C36768A",
    x"2C365FBD",
    x"2C3648F2",
    x"2C36322A",
    x"2C361B66",
    x"2C3604A4",
    x"2C35EDE4",
    x"2C35D728",
    x"2C35C06F",
    x"2C35A9B8",
    x"2C359304",
    x"2C357C53",
    x"2C3565A5",
    x"2C354EFA",
    x"2C353851",
    x"2C3521AC",
    x"2C350B09",
    x"2C34F469",
    x"2C34DDCC",
    x"2C34C731",
    x"2C34B09A",
    x"2C349A05",
    x"2C348373",
    x"2C346CE4",
    x"2C345658",
    x"2C343FCF",
    x"2C342948",
    x"2C3412C5",
    x"2C33FC44",
    x"2C33E5C5",
    x"2C33CF4A",
    x"2C33B8D2",
    x"2C33A25C",
    x"2C338BE9",
    x"2C337579",
    x"2C335F0C",
    x"2C3348A1",
    x"2C33323A",
    x"2C331BD5",
    x"2C330573",
    x"2C32EF13",
    x"2C32D8B7",
    x"2C32C25D",
    x"2C32AC06",
    x"2C3295B2",
    x"2C327F61",
    x"2C326912",
    x"2C3252C7",
    x"2C323C7E",
    x"2C322637",
    x"2C320FF4",
    x"2C31F9B3",
    x"2C31E376",
    x"2C31CD3B",
    x"2C31B702",
    x"2C31A0CD",
    x"2C318A9A",
    x"2C31746A",
    x"2C315E3D",
    x"2C314813",
    x"2C3131EB",
    x"2C311BC6",
    x"2C3105A4",
    x"2C30EF85",
    x"2C30D968",
    x"2C30C34E",
    x"2C30AD37",
    x"2C309723",
    x"2C308112",
    x"2C306B03",
    x"2C3054F7",
    x"2C303EEE",
    x"2C3028E7",
    x"2C3012E3",
    x"2C2FFCE2",
    x"2C2FE6E4",
    x"2C2FD0E9",
    x"2C2FBAF0",
    x"2C2FA4FA",
    x"2C2F8F07",
    x"2C2F7916",
    x"2C2F6328",
    x"2C2F4D3D",
    x"2C2F3755",
    x"2C2F216F",
    x"2C2F0B8D",
    x"2C2EF5AD",
    x"2C2EDFCF",
    x"2C2EC9F5",
    x"2C2EB41D",
    x"2C2E9E48",
    x"2C2E8875",
    x"2C2E72A6",
    x"2C2E5CD9",
    x"2C2E470E",
    x"2C2E3147",
    x"2C2E1B82",
    x"2C2E05C0",
    x"2C2DF001",
    x"2C2DDA44",
    x"2C2DC48A",
    x"2C2DAED3",
    x"2C2D991E",
    x"2C2D836C",
    x"2C2D6DBD",
    x"2C2D5811",
    x"2C2D4267",
    x"2C2D2CC0",
    x"2C2D171C",
    x"2C2D017B",
    x"2C2CEBDC",
    x"2C2CD640",
    x"2C2CC0A6",
    x"2C2CAB10",
    x"2C2C957C",
    x"2C2C7FEA",
    x"2C2C6A5C",
    x"2C2C54D0",
    x"2C2C3F46",
    x"2C2C29C0",
    x"2C2C143C",
    x"2C2BFEBB",
    x"2C2BE93C",
    x"2C2BD3C0",
    x"2C2BBE47",
    x"2C2BA8D1",
    x"2C2B935D",
    x"2C2B7DEC",
    x"2C2B687E",
    x"2C2B5312",
    x"2C2B3DA9",
    x"2C2B2842",
    x"2C2B12DF",
    x"2C2AFD7E",
    x"2C2AE81F",
    x"2C2AD2C4",
    x"2C2ABD6B",
    x"2C2AA814",
    x"2C2A92C1",
    x"2C2A7D70",
    x"2C2A6821",
    x"2C2A52D6",
    x"2C2A3D8D",
    x"2C2A2846",
    x"2C2A1303",
    x"2C29FDC1",
    x"2C29E883",
    x"2C29D347",
    x"2C29BE0E",
    x"2C29A8D8",
    x"2C2993A4",
    x"2C297E73",
    x"2C296944",
    x"2C295419",
    x"2C293EEF",
    x"2C2929C9",
    x"2C2914A5",
    x"2C28FF84",
    x"2C28EA65",
    x"2C28D549",
    x"2C28C030",
    x"2C28AB19",
    x"2C289605",
    x"2C2880F4",
    x"2C286BE5",
    x"2C2856D9",
    x"2C2841CF",
    x"2C282CC8",
    x"2C2817C4",
    x"2C2802C2",
    x"2C27EDC3",
    x"2C27D8C7",
    x"2C27C3CD",
    x"2C27AED6",
    x"2C2799E1",
    x"2C2784EF",
    x"2C277000",
    x"2C275B13",
    x"2C274629",
    x"2C273142",
    x"2C271C5D",
    x"2C27077B",
    x"2C26F29B",
    x"2C26DDBE",
    x"2C26C8E4",
    x"2C26B40C",
    x"2C269F37",
    x"2C268A64",
    x"2C267594",
    x"2C2660C7",
    x"2C264BFC",
    x"2C263734",
    x"2C26226E",
    x"2C260DAB",
    x"2C25F8EB",
    x"2C25E42D",
    x"2C25CF72",
    x"2C25BAB9",
    x"2C25A603",
    x"2C25914F",
    x"2C257C9F",
    x"2C2567F0",
    x"2C255345",
    x"2C253E9B",
    x"2C2529F5",
    x"2C251551",
    x"2C2500B0",
    x"2C24EC11",
    x"2C24D775",
    x"2C24C2DB",
    x"2C24AE44",
    x"2C2499AF",
    x"2C24851D",
    x"2C24708E",
    x"2C245C01",
    x"2C244777",
    x"2C2432EF",
    x"2C241E6A",
    x"2C2409E8",
    x"2C23F568",
    x"2C23E0EA",
    x"2C23CC70",
    x"2C23B7F7",
    x"2C23A382",
    x"2C238F0E",
    x"2C237A9E",
    x"2C236630",
    x"2C2351C4",
    x"2C233D5B",
    x"2C2328F5",
    x"2C231491",
    x"2C230030",
    x"2C22EBD1",
    x"2C22D775",
    x"2C22C31B",
    x"2C22AEC4",
    x"2C229A70",
    x"2C22861E",
    x"2C2271CE",
    x"2C225D81",
    x"2C224937",
    x"2C2234EF",
    x"2C2220A9",
    x"2C220C67",
    x"2C21F826",
    x"2C21E3E9",
    x"2C21CFAD",
    x"2C21BB75",
    x"2C21A73E",
    x"2C21930B",
    x"2C217EDA",
    x"2C216AAB",
    x"2C21567F",
    x"2C214255",
    x"2C212E2E",
    x"2C211A0A",
    x"2C2105E8",
    x"2C20F1C8",
    x"2C20DDAB",
    x"2C20C991",
    x"2C20B579",
    x"2C20A164",
    x"2C208D51",
    x"2C207940",
    x"2C206532",
    x"2C205127",
    x"2C203D1E",
    x"2C202918",
    x"2C201514",
    x"2C200113",
    x"2C1FED14",
    x"2C1FD917",
    x"2C1FC51D",
    x"2C1FB126",
    x"2C1F9D31",
    x"2C1F893F",
    x"2C1F754F",
    x"2C1F6161",
    x"2C1F4D76",
    x"2C1F398E",
    x"2C1F25A8",
    x"2C1F11C5",
    x"2C1EFDE4",
    x"2C1EEA05",
    x"2C1ED629",
    x"2C1EC250",
    x"2C1EAE78",
    x"2C1E9AA4",
    x"2C1E86D2",
    x"2C1E7302",
    x"2C1E5F35",
    x"2C1E4B6A",
    x"2C1E37A2",
    x"2C1E23DC",
    x"2C1E1019",
    x"2C1DFC58",
    x"2C1DE89A",
    x"2C1DD4DE",
    x"2C1DC125",
    x"2C1DAD6E",
    x"2C1D99BA",
    x"2C1D8608",
    x"2C1D7258",
    x"2C1D5EAB",
    x"2C1D4B00",
    x"2C1D3758",
    x"2C1D23B3",
    x"2C1D100F",
    x"2C1CFC6F",
    x"2C1CE8D0",
    x"2C1CD534",
    x"2C1CC19B",
    x"2C1CAE04",
    x"2C1C9A6F",
    x"2C1C86DD",
    x"2C1C734E",
    x"2C1C5FC1",
    x"2C1C4C36",
    x"2C1C38AD",
    x"2C1C2528",
    x"2C1C11A4",
    x"2C1BFE23",
    x"2C1BEAA5",
    x"2C1BD729",
    x"2C1BC3AF",
    x"2C1BB038",
    x"2C1B9CC3",
    x"2C1B8950",
    x"2C1B75E0",
    x"2C1B6273",
    x"2C1B4F08",
    x"2C1B3B9F",
    x"2C1B2839",
    x"2C1B14D5",
    x"2C1B0174",
    x"2C1AEE15",
    x"2C1ADAB8",
    x"2C1AC75E",
    x"2C1AB406",
    x"2C1AA0B1",
    x"2C1A8D5E",
    x"2C1A7A0E",
    x"2C1A66C0",
    x"2C1A5374",
    x"2C1A402B",
    x"2C1A2CE4",
    x"2C1A19A0",
    x"2C1A065E",
    x"2C19F31E",
    x"2C19DFE1",
    x"2C19CCA6",
    x"2C19B96E",
    x"2C19A638",
    x"2C199304",
    x"2C197FD3",
    x"2C196CA4",
    x"2C195978",
    x"2C19464E",
    x"2C193326",
    x"2C192001",
    x"2C190CDE",
    x"2C18F9BE",
    x"2C18E6A0",
    x"2C18D384",
    x"2C18C06B",
    x"2C18AD54",
    x"2C189A40",
    x"2C18872D",
    x"2C18741E",
    x"2C186110",
    x"2C184E05",
    x"2C183AFD",
    x"2C1827F7",
    x"2C1814F3",
    x"2C1801F1",
    x"2C17EEF2",
    x"2C17DBF6",
    x"2C17C8FB",
    x"2C17B604",
    x"2C17A30E",
    x"2C17901B",
    x"2C177D2A",
    x"2C176A3B",
    x"2C17574F",
    x"2C174466",
    x"2C17317E",
    x"2C171E99",
    x"2C170BB7",
    x"2C16F8D6",
    x"2C16E5F8",
    x"2C16D31D",
    x"2C16C044",
    x"2C16AD6D",
    x"2C169A98",
    x"2C1687C6",
    x"2C1674F6",
    x"2C166229",
    x"2C164F5E",
    x"2C163C95",
    x"2C1629CF",
    x"2C16170B",
    x"2C160449",
    x"2C15F18A",
    x"2C15DECC",
    x"2C15CC12",
    x"2C15B959",
    x"2C15A6A3",
    x"2C1593F0",
    x"2C15813E",
    x"2C156E90",
    x"2C155BE3",
    x"2C154939",
    x"2C153691",
    x"2C1523EB",
    x"2C151148",
    x"2C14FEA7",
    x"2C14EC08",
    x"2C14D96C",
    x"2C14C6D2",
    x"2C14B43A",
    x"2C14A1A4",
    x"2C148F11",
    x"2C147C81",
    x"2C1469F2",
    x"2C145766",
    x"2C1444DC",
    x"2C143255",
    x"2C141FD0",
    x"2C140D4D",
    x"2C13FACD",
    x"2C13E84E",
    x"2C13D5D2",
    x"2C13C359",
    x"2C13B0E2",
    x"2C139E6D",
    x"2C138BFA",
    x"2C13798A",
    x"2C13671C",
    x"2C1354B0",
    x"2C134246",
    x"2C132FDF",
    x"2C131D7B",
    x"2C130B18",
    x"2C12F8B8",
    x"2C12E65A",
    x"2C12D3FE",
    x"2C12C1A5",
    x"2C12AF4E",
    x"2C129CF9",
    x"2C128AA6",
    x"2C127856",
    x"2C126608",
    x"2C1253BD",
    x"2C124173",
    x"2C122F2C",
    x"2C121CE8",
    x"2C120AA5",
    x"2C11F865",
    x"2C11E627",
    x"2C11D3EB",
    x"2C11C1B2",
    x"2C11AF7B",
    x"2C119D46",
    x"2C118B14",
    x"2C1178E3",
    x"2C1166B6",
    x"2C11548A",
    x"2C114260",
    x"2C113039",
    x"2C111E14",
    x"2C110BF2",
    x"2C10F9D1",
    x"2C10E7B3",
    x"2C10D597",
    x"2C10C37E",
    x"2C10B167",
    x"2C109F51",
    x"2C108D3F",
    x"2C107B2E",
    x"2C106920",
    x"2C105714",
    x"2C10450A",
    x"2C103303",
    x"2C1020FD",
    x"2C100EFA",
    x"2C0FFCFA",
    x"2C0FEAFB",
    x"2C0FD8FF",
    x"2C0FC705",
    x"2C0FB50D",
    x"2C0FA318",
    x"2C0F9124",
    x"2C0F7F33",
    x"2C0F6D45",
    x"2C0F5B58",
    x"2C0F496E",
    x"2C0F3786",
    x"2C0F25A0",
    x"2C0F13BC",
    x"2C0F01DB",
    x"2C0EEFFC",
    x"2C0EDE1F",
    x"2C0ECC44",
    x"2C0EBA6C",
    x"2C0EA896",
    x"2C0E96C2",
    x"2C0E84F0",
    x"2C0E7320",
    x"2C0E6153",
    x"2C0E4F88",
    x"2C0E3DBF",
    x"2C0E2BF9",
    x"2C0E1A34",
    x"2C0E0872",
    x"2C0DF6B2",
    x"2C0DE4F4",
    x"2C0DD339",
    x"2C0DC180",
    x"2C0DAFC9",
    x"2C0D9E14",
    x"2C0D8C61",
    x"2C0D7AB1",
    x"2C0D6902",
    x"2C0D5756",
    x"2C0D45AD",
    x"2C0D3405",
    x"2C0D2260",
    x"2C0D10BC",
    x"2C0CFF1B",
    x"2C0CED7D",
    x"2C0CDBE0",
    x"2C0CCA46",
    x"2C0CB8AD",
    x"2C0CA717",
    x"2C0C9584",
    x"2C0C83F2",
    x"2C0C7263",
    x"2C0C60D5",
    x"2C0C4F4A",
    x"2C0C3DC2",
    x"2C0C2C3B",
    x"2C0C1AB7",
    x"2C0C0934",
    x"2C0BF7B4",
    x"2C0BE636",
    x"2C0BD4BB",
    x"2C0BC341",
    x"2C0BB1CA",
    x"2C0BA055",
    x"2C0B8EE2",
    x"2C0B7D71",
    x"2C0B6C02",
    x"2C0B5A96",
    x"2C0B492C",
    x"2C0B37C4",
    x"2C0B265E",
    x"2C0B14FA",
    x"2C0B0399",
    x"2C0AF239",
    x"2C0AE0DC",
    x"2C0ACF81",
    x"2C0ABE28",
    x"2C0AACD2",
    x"2C0A9B7D",
    x"2C0A8A2B",
    x"2C0A78DA",
    x"2C0A678C",
    x"2C0A5641",
    x"2C0A44F7",
    x"2C0A33AF",
    x"2C0A226A",
    x"2C0A1127",
    x"2C09FFE6",
    x"2C09EEA7",
    x"2C09DD6A",
    x"2C09CC2F",
    x"2C09BAF7",
    x"2C09A9C1",
    x"2C09988D",
    x"2C09875B",
    x"2C09762B",
    x"2C0964FD",
    x"2C0953D1",
    x"2C0942A8",
    x"2C093181",
    x"2C09205C",
    x"2C090F39",
    x"2C08FE18",
    x"2C08ECF9",
    x"2C08DBDD",
    x"2C08CAC2",
    x"2C08B9AA",
    x"2C08A894",
    x"2C089780",
    x"2C08866E",
    x"2C08755E",
    x"2C086451",
    x"2C085345",
    x"2C08423C",
    x"2C083135",
    x"2C08202F",
    x"2C080F2C",
    x"2C07FE2C",
    x"2C07ED2D",
    x"2C07DC30",
    x"2C07CB36",
    x"2C07BA3E",
    x"2C07A947",
    x"2C079853",
    x"2C078761",
    x"2C077671",
    x"2C076584",
    x"2C075498",
    x"2C0743AE",
    x"2C0732C7",
    x"2C0721E2",
    x"2C0710FF",
    x"2C07001E",
    x"2C06EF3F",
    x"2C06DE62",
    x"2C06CD87",
    x"2C06BCAE",
    x"2C06ABD8",
    x"2C069B03",
    x"2C068A31",
    x"2C067961",
    x"2C066893",
    x"2C0657C7",
    x"2C0646FD",
    x"2C063635",
    x"2C06256F",
    x"2C0614AC",
    x"2C0603EA",
    x"2C05F32B",
    x"2C05E26D",
    x"2C05D1B2",
    x"2C05C0F9",
    x"2C05B042",
    x"2C059F8D",
    x"2C058EDA",
    x"2C057E29",
    x"2C056D7A",
    x"2C055CCE",
    x"2C054C23",
    x"2C053B7B",
    x"2C052AD4",
    x"2C051A30",
    x"2C05098E",
    x"2C04F8EE",
    x"2C04E84F",
    x"2C04D7B3",
    x"2C04C71A",
    x"2C04B682",
    x"2C04A5EC",
    x"2C049558",
    x"2C0484C7",
    x"2C047437",
    x"2C0463AA",
    x"2C04531E",
    x"2C044295",
    x"2C04320D",
    x"2C042188",
    x"2C041105",
    x"2C040084",
    x"2C03F005",
    x"2C03DF88",
    x"2C03CF0D",
    x"2C03BE94",
    x"2C03AE1D",
    x"2C039DA9",
    x"2C038D36",
    x"2C037CC5",
    x"2C036C57",
    x"2C035BEA",
    x"2C034B80",
    x"2C033B17",
    x"2C032AB1",
    x"2C031A4D",
    x"2C0309EA",
    x"2C02F98A",
    x"2C02E92C",
    x"2C02D8D0",
    x"2C02C876",
    x"2C02B81E",
    x"2C02A7C8",
    x"2C029774",
    x"2C028722",
    x"2C0276D2",
    x"2C026684",
    x"2C025639",
    x"2C0245EF",
    x"2C0235A7",
    x"2C022561",
    x"2C02151E",
    x"2C0204DC",
    x"2C01F49C",
    x"2C01E45F",
    x"2C01D423",
    x"2C01C3EA",
    x"2C01B3B2",
    x"2C01A37D",
    x"2C01934A",
    x"2C018318",
    x"2C0172E9",
    x"2C0162BB",
    x"2C015290",
    x"2C014267",
    x"2C01323F",
    x"2C01221A",
    x"2C0111F7",
    x"2C0101D6",
    x"2C00F1B6",
    x"2C00E199",
    x"2C00D17E",
    x"2C00C165",
    x"2C00B14E",
    x"2C00A139",
    x"2C009125",
    x"2C008114",
    x"2C007105",
    x"2C0060F8",
    x"2C0050ED",
    x"2C0040E4",
    x"2C0030DD",
    x"2C0020D8",
    x"2C0010D4",
    x"2C0000D3",
    x"2BFFE1A9",
    x"2BFFC1AE",
    x"2BFFA1B8",
    x"2BFF81C6",
    x"2BFF61D8",
    x"2BFF41ED",
    x"2BFF2207",
    x"2BFF0225",
    x"2BFEE247",
    x"2BFEC26C",
    x"2BFEA296",
    x"2BFE82C4",
    x"2BFE62F5",
    x"2BFE432B",
    x"2BFE2365",
    x"2BFE03A2",
    x"2BFDE3E4",
    x"2BFDC429",
    x"2BFDA473",
    x"2BFD84C0",
    x"2BFD6511",
    x"2BFD4567",
    x"2BFD25C0",
    x"2BFD061D",
    x"2BFCE67F",
    x"2BFCC6E4",
    x"2BFCA74D",
    x"2BFC87BA",
    x"2BFC682B",
    x"2BFC48A0",
    x"2BFC2919",
    x"2BFC0996",
    x"2BFBEA16",
    x"2BFBCA9B",
    x"2BFBAB24",
    x"2BFB8BB0",
    x"2BFB6C41",
    x"2BFB4CD5",
    x"2BFB2D6E",
    x"2BFB0E0A",
    x"2BFAEEAA",
    x"2BFACF4E",
    x"2BFAAFF6",
    x"2BFA90A2",
    x"2BFA7152",
    x"2BFA5206",
    x"2BFA32BE",
    x"2BFA1379",
    x"2BF9F439",
    x"2BF9D4FC",
    x"2BF9B5C3",
    x"2BF9968F",
    x"2BF9775E",
    x"2BF95831",
    x"2BF93908",
    x"2BF919E3",
    x"2BF8FAC1",
    x"2BF8DBA4",
    x"2BF8BC8A",
    x"2BF89D75",
    x"2BF87E63",
    x"2BF85F55",
    x"2BF8404B",
    x"2BF82145",
    x"2BF80243",
    x"2BF7E345",
    x"2BF7C44A",
    x"2BF7A553",
    x"2BF78661",
    x"2BF76772",
    x"2BF74887",
    x"2BF729A0",
    x"2BF70ABC",
    x"2BF6EBDD",
    x"2BF6CD01",
    x"2BF6AE2A",
    x"2BF68F56",
    x"2BF67086",
    x"2BF651BA",
    x"2BF632F2",
    x"2BF6142D",
    x"2BF5F56C",
    x"2BF5D6B0",
    x"2BF5B7F7",
    x"2BF59942",
    x"2BF57A90",
    x"2BF55BE3",
    x"2BF53D3A",
    x"2BF51E94",
    x"2BF4FFF2",
    x"2BF4E154",
    x"2BF4C2BA",
    x"2BF4A423",
    x"2BF48590",
    x"2BF46702",
    x"2BF44877",
    x"2BF429F0",
    x"2BF40B6C",
    x"2BF3ECED",
    x"2BF3CE71",
    x"2BF3AFF9",
    x"2BF39185",
    x"2BF37315",
    x"2BF354A8",
    x"2BF33640",
    x"2BF317DB",
    x"2BF2F97A",
    x"2BF2DB1C",
    x"2BF2BCC3",
    x"2BF29E6D",
    x"2BF2801B",
    x"2BF261CD",
    x"2BF24383",
    x"2BF2253C",
    x"2BF206F9",
    x"2BF1E8BA",
    x"2BF1CA7F",
    x"2BF1AC48",
    x"2BF18E14",
    x"2BF16FE4",
    x"2BF151B8",
    x"2BF13390",
    x"2BF1156B",
    x"2BF0F74B",
    x"2BF0D92E",
    x"2BF0BB14",
    x"2BF09CFF",
    x"2BF07EED",
    x"2BF060DF",
    x"2BF042D5",
    x"2BF024CE",
    x"2BF006CC",
    x"2BEFE8CD",
    x"2BEFCAD1",
    x"2BEFACDA",
    x"2BEF8EE6",
    x"2BEF70F6",
    x"2BEF530A",
    x"2BEF3521",
    x"2BEF173D",
    x"2BEEF95C",
    x"2BEEDB7E",
    x"2BEEBDA5",
    x"2BEE9FCF",
    x"2BEE81FD",
    x"2BEE642E",
    x"2BEE4664",
    x"2BEE289D",
    x"2BEE0ADA",
    x"2BEDED1A",
    x"2BEDCF5E",
    x"2BEDB1A6",
    x"2BED93F2",
    x"2BED7641",
    x"2BED5894",
    x"2BED3AEB",
    x"2BED1D46",
    x"2BECFFA4",
    x"2BECE206",
    x"2BECC46B",
    x"2BECA6D5",
    x"2BEC8942",
    x"2BEC6BB2",
    x"2BEC4E27",
    x"2BEC309F",
    x"2BEC131B",
    x"2BEBF59A",
    x"2BEBD81D",
    x"2BEBBAA4",
    x"2BEB9D2E",
    x"2BEB7FBD",
    x"2BEB624F",
    x"2BEB44E4",
    x"2BEB277D",
    x"2BEB0A1A",
    x"2BEAECBB",
    x"2BEACF5F",
    x"2BEAB207",
    x"2BEA94B2",
    x"2BEA7762",
    x"2BEA5A15",
    x"2BEA3CCB",
    x"2BEA1F85",
    x"2BEA0243",
    x"2BE9E505",
    x"2BE9C7CA",
    x"2BE9AA93",
    x"2BE98D5F",
    x"2BE97030",
    x"2BE95303",
    x"2BE935DB",
    x"2BE918B6",
    x"2BE8FB95",
    x"2BE8DE77",
    x"2BE8C15D",
    x"2BE8A447",
    x"2BE88734",
    x"2BE86A25",
    x"2BE84D19",
    x"2BE83012",
    x"2BE8130D",
    x"2BE7F60D",
    x"2BE7D910",
    x"2BE7BC17",
    x"2BE79F21",
    x"2BE7822F",
    x"2BE76540",
    x"2BE74855",
    x"2BE72B6E",
    x"2BE70E8B",
    x"2BE6F1AB",
    x"2BE6D4CE",
    x"2BE6B7F5",
    x"2BE69B20",
    x"2BE67E4F",
    x"2BE66181",
    x"2BE644B6",
    x"2BE627EF",
    x"2BE60B2C",
    x"2BE5EE6D",
    x"2BE5D1B1",
    x"2BE5B4F8",
    x"2BE59843",
    x"2BE57B92",
    x"2BE55EE5",
    x"2BE5423A",
    x"2BE52594",
    x"2BE508F1",
    x"2BE4EC52",
    x"2BE4CFB6",
    x"2BE4B31E",
    x"2BE49689",
    x"2BE479F8",
    x"2BE45D6B",
    x"2BE440E1",
    x"2BE4245A",
    x"2BE407D8",
    x"2BE3EB59",
    x"2BE3CEDD",
    x"2BE3B265",
    x"2BE395F0",
    x"2BE3797F",
    x"2BE35D12",
    x"2BE340A8",
    x"2BE32442",
    x"2BE307DF",
    x"2BE2EB80",
    x"2BE2CF24",
    x"2BE2B2CC",
    x"2BE29677",
    x"2BE27A26",
    x"2BE25DD9",
    x"2BE2418F",
    x"2BE22548",
    x"2BE20906",
    x"2BE1ECC6",
    x"2BE1D08A",
    x"2BE1B452",
    x"2BE1981D",
    x"2BE17BEC",
    x"2BE15FBE",
    x"2BE14394",
    x"2BE1276D",
    x"2BE10B4A",
    x"2BE0EF2B",
    x"2BE0D30E",
    x"2BE0B6F6",
    x"2BE09AE1",
    x"2BE07ECF",
    x"2BE062C1",
    x"2BE046B6",
    x"2BE02AAF",
    x"2BE00EAC",
    x"2BDFF2AC",
    x"2BDFD6AF",
    x"2BDFBAB6",
    x"2BDF9EC0",
    x"2BDF82CE",
    x"2BDF66E0",
    x"2BDF4AF5",
    x"2BDF2F0D",
    x"2BDF1329",
    x"2BDEF748",
    x"2BDEDB6B",
    x"2BDEBF91",
    x"2BDEA3BB",
    x"2BDE87E8",
    x"2BDE6C19",
    x"2BDE504D",
    x"2BDE3485",
    x"2BDE18C0",
    x"2BDDFCFF",
    x"2BDDE141",
    x"2BDDC587",
    x"2BDDA9D0",
    x"2BDD8E1C",
    x"2BDD726C",
    x"2BDD56C0",
    x"2BDD3B16",
    x"2BDD1F71",
    x"2BDD03CF",
    x"2BDCE830",
    x"2BDCCC95",
    x"2BDCB0FD",
    x"2BDC9568",
    x"2BDC79D7",
    x"2BDC5E4A",
    x"2BDC42C0",
    x"2BDC2739",
    x"2BDC0BB6",
    x"2BDBF036",
    x"2BDBD4BA",
    x"2BDBB941",
    x"2BDB9DCC",
    x"2BDB825A",
    x"2BDB66EB",
    x"2BDB4B80",
    x"2BDB3018",
    x"2BDB14B4",
    x"2BDAF953",
    x"2BDADDF5",
    x"2BDAC29B",
    x"2BDAA745",
    x"2BDA8BF2",
    x"2BDA70A2",
    x"2BDA5555",
    x"2BDA3A0C",
    x"2BDA1EC7",
    x"2BDA0385",
    x"2BD9E846",
    x"2BD9CD0B",
    x"2BD9B1D3",
    x"2BD9969E",
    x"2BD97B6D",
    x"2BD9603F",
    x"2BD94515",
    x"2BD929EE",
    x"2BD90ECB",
    x"2BD8F3AA",
    x"2BD8D88E",
    x"2BD8BD74",
    x"2BD8A25E",
    x"2BD8874C",
    x"2BD86C3C",
    x"2BD85131",
    x"2BD83628",
    x"2BD81B23",
    x"2BD80021",
    x"2BD7E523",
    x"2BD7CA28",
    x"2BD7AF31",
    x"2BD7943C",
    x"2BD7794B",
    x"2BD75E5E",
    x"2BD74374",
    x"2BD7288D",
    x"2BD70DAA",
    x"2BD6F2CA",
    x"2BD6D7ED",
    x"2BD6BD14",
    x"2BD6A23E",
    x"2BD6876B",
    x"2BD66C9C",
    x"2BD651D0",
    x"2BD63707",
    x"2BD61C42",
    x"2BD60180",
    x"2BD5E6C2",
    x"2BD5CC07",
    x"2BD5B14F",
    x"2BD5969A",
    x"2BD57BE9",
    x"2BD5613B",
    x"2BD54691",
    x"2BD52BEA",
    x"2BD51146",
    x"2BD4F6A5",
    x"2BD4DC08",
    x"2BD4C16E",
    x"2BD4A6D8",
    x"2BD48C45",
    x"2BD471B5",
    x"2BD45728",
    x"2BD43C9F",
    x"2BD42219",
    x"2BD40797",
    x"2BD3ED17",
    x"2BD3D29B",
    x"2BD3B823",
    x"2BD39DAD",
    x"2BD3833B",
    x"2BD368CC",
    x"2BD34E61",
    x"2BD333F9",
    x"2BD31994",
    x"2BD2FF32",
    x"2BD2E4D4",
    x"2BD2CA79",
    x"2BD2B022",
    x"2BD295CD",
    x"2BD27B7C",
    x"2BD2612E",
    x"2BD246E4",
    x"2BD22C9D",
    x"2BD21259",
    x"2BD1F818",
    x"2BD1DDDB",
    x"2BD1C3A1",
    x"2BD1A96A",
    x"2BD18F36",
    x"2BD17506",
    x"2BD15AD9",
    x"2BD140AF",
    x"2BD12689",
    x"2BD10C66",
    x"2BD0F246",
    x"2BD0D829",
    x"2BD0BE10",
    x"2BD0A3F9",
    x"2BD089E7",
    x"2BD06FD7",
    x"2BD055CB",
    x"2BD03BC2",
    x"2BD021BC",
    x"2BD007B9",
    x"2BCFEDBA",
    x"2BCFD3BE",
    x"2BCFB9C5",
    x"2BCF9FCF",
    x"2BCF85DD",
    x"2BCF6BEE",
    x"2BCF5202",
    x"2BCF3819",
    x"2BCF1E34",
    x"2BCF0452",
    x"2BCEEA73",
    x"2BCED097",
    x"2BCEB6BF",
    x"2BCE9CE9",
    x"2BCE8317",
    x"2BCE6949",
    x"2BCE4F7D",
    x"2BCE35B5",
    x"2BCE1BF0",
    x"2BCE022E",
    x"2BCDE86F",
    x"2BCDCEB4",
    x"2BCDB4FB",
    x"2BCD9B46",
    x"2BCD8195",
    x"2BCD67E6",
    x"2BCD4E3B",
    x"2BCD3493",
    x"2BCD1AEE",
    x"2BCD014C",
    x"2BCCE7AD",
    x"2BCCCE12",
    x"2BCCB47A",
    x"2BCC9AE5",
    x"2BCC8153",
    x"2BCC67C4",
    x"2BCC4E39",
    x"2BCC34B1",
    x"2BCC1B2C",
    x"2BCC01AA",
    x"2BCBE82B",
    x"2BCBCEB0",
    x"2BCBB538",
    x"2BCB9BC3",
    x"2BCB8251",
    x"2BCB68E2",
    x"2BCB4F77",
    x"2BCB360E",
    x"2BCB1CA9",
    x"2BCB0347",
    x"2BCAE9E8",
    x"2BCAD08D",
    x"2BCAB734",
    x"2BCA9DDF",
    x"2BCA848D",
    x"2BCA6B3E",
    x"2BCA51F2",
    x"2BCA38A9",
    x"2BCA1F64",
    x"2BCA0621",
    x"2BC9ECE2",
    x"2BC9D3A6",
    x"2BC9BA6D",
    x"2BC9A138",
    x"2BC98805",
    x"2BC96ED6",
    x"2BC955A9",
    x"2BC93C80",
    x"2BC9235A",
    x"2BC90A37",
    x"2BC8F118",
    x"2BC8D7FB",
    x"2BC8BEE2",
    x"2BC8A5CB",
    x"2BC88CB8",
    x"2BC873A8",
    x"2BC85A9B",
    x"2BC84191",
    x"2BC8288B",
    x"2BC80F87",
    x"2BC7F687",
    x"2BC7DD8A",
    x"2BC7C490",
    x"2BC7AB99",
    x"2BC792A5",
    x"2BC779B4",
    x"2BC760C6",
    x"2BC747DC",
    x"2BC72EF4",
    x"2BC71610",
    x"2BC6FD2F",
    x"2BC6E451",
    x"2BC6CB76",
    x"2BC6B29E",
    x"2BC699C9",
    x"2BC680F7",
    x"2BC66829",
    x"2BC64F5D",
    x"2BC63695",
    x"2BC61DD0",
    x"2BC6050D",
    x"2BC5EC4E",
    x"2BC5D392",
    x"2BC5BAD9",
    x"2BC5A224",
    x"2BC58971",
    x"2BC570C1",
    x"2BC55815",
    x"2BC53F6B",
    x"2BC526C5",
    x"2BC50E22",
    x"2BC4F581",
    x"2BC4DCE4",
    x"2BC4C44A",
    x"2BC4ABB3",
    x"2BC4931F",
    x"2BC47A8E",
    x"2BC46201",
    x"2BC44976",
    x"2BC430EE",
    x"2BC4186A",
    x"2BC3FFE8",
    x"2BC3E76A",
    x"2BC3CEEE",
    x"2BC3B676",
    x"2BC39E01",
    x"2BC3858E",
    x"2BC36D1F",
    x"2BC354B3",
    x"2BC33C4A",
    x"2BC323E4",
    x"2BC30B81",
    x"2BC2F321",
    x"2BC2DAC4",
    x"2BC2C26A",
    x"2BC2AA14",
    x"2BC291C0",
    x"2BC2796F",
    x"2BC26122",
    x"2BC248D7",
    x"2BC2308F",
    x"2BC2184B",
    x"2BC20009",
    x"2BC1E7CB",
    x"2BC1CF8F",
    x"2BC1B757",
    x"2BC19F22",
    x"2BC186EF",
    x"2BC16EC0",
    x"2BC15693",
    x"2BC13E6A",
    x"2BC12644",
    x"2BC10E21",
    x"2BC0F600",
    x"2BC0DDE3",
    x"2BC0C5C9",
    x"2BC0ADB2",
    x"2BC0959D",
    x"2BC07D8C",
    x"2BC0657E",
    x"2BC04D73",
    x"2BC0356B",
    x"2BC01D66",
    x"2BC00563",
    x"2BBFED64",
    x"2BBFD568",
    x"2BBFBD6F",
    x"2BBFA579",
    x"2BBF8D85",
    x"2BBF7595",
    x"2BBF5DA8",
    x"2BBF45BE",
    x"2BBF2DD7",
    x"2BBF15F2",
    x"2BBEFE11",
    x"2BBEE633",
    x"2BBECE58",
    x"2BBEB67F",
    x"2BBE9EAA",
    x"2BBE86D8",
    x"2BBE6F08",
    x"2BBE573C",
    x"2BBE3F72",
    x"2BBE27AC",
    x"2BBE0FE9",
    x"2BBDF828",
    x"2BBDE06A",
    x"2BBDC8B0",
    x"2BBDB0F8",
    x"2BBD9944",
    x"2BBD8192",
    x"2BBD69E3",
    x"2BBD5238",
    x"2BBD3A8F",
    x"2BBD22E9",
    x"2BBD0B46",
    x"2BBCF3A6",
    x"2BBCDC09",
    x"2BBCC46F",
    x"2BBCACD8",
    x"2BBC9544",
    x"2BBC7DB3",
    x"2BBC6624",
    x"2BBC4E99",
    x"2BBC3711",
    x"2BBC1F8B",
    x"2BBC0809",
    x"2BBBF089",
    x"2BBBD90D",
    x"2BBBC193",
    x"2BBBAA1C",
    x"2BBB92A9",
    x"2BBB7B38",
    x"2BBB63CA",
    x"2BBB4C5F",
    x"2BBB34F7",
    x"2BBB1D91",
    x"2BBB062F",
    x"2BBAEED0",
    x"2BBAD774",
    x"2BBAC01A",
    x"2BBAA8C4",
    x"2BBA9170",
    x"2BBA7A1F",
    x"2BBA62D1",
    x"2BBA4B86",
    x"2BBA343E",
    x"2BBA1CF9",
    x"2BBA05B7",
    x"2BB9EE78",
    x"2BB9D73C",
    x"2BB9C002",
    x"2BB9A8CC",
    x"2BB99198",
    x"2BB97A67",
    x"2BB96339",
    x"2BB94C0E",
    x"2BB934E6",
    x"2BB91DC1",
    x"2BB9069F",
    x"2BB8EF80",
    x"2BB8D863",
    x"2BB8C149",
    x"2BB8AA33",
    x"2BB8931F",
    x"2BB87C0E",
    x"2BB86500",
    x"2BB84DF5",
    x"2BB836EC",
    x"2BB81FE7",
    x"2BB808E4",
    x"2BB7F1E5",
    x"2BB7DAE8",
    x"2BB7C3EE",
    x"2BB7ACF7",
    x"2BB79603",
    x"2BB77F11",
    x"2BB76823",
    x"2BB75137",
    x"2BB73A4F",
    x"2BB72369",
    x"2BB70C86",
    x"2BB6F5A6",
    x"2BB6DEC8",
    x"2BB6C7EE",
    x"2BB6B116",
    x"2BB69A42",
    x"2BB68370",
    x"2BB66CA1",
    x"2BB655D5",
    x"2BB63F0B",
    x"2BB62845",
    x"2BB61181",
    x"2BB5FAC1",
    x"2BB5E403",
    x"2BB5CD48",
    x"2BB5B68F",
    x"2BB59FDA",
    x"2BB58927",
    x"2BB57278",
    x"2BB55BCB",
    x"2BB54521",
    x"2BB52E79",
    x"2BB517D5",
    x"2BB50134",
    x"2BB4EA95",
    x"2BB4D3F9",
    x"2BB4BD60",
    x"2BB4A6CA",
    x"2BB49036",
    x"2BB479A5",
    x"2BB46318",
    x"2BB44C8D",
    x"2BB43605",
    x"2BB41F7F",
    x"2BB408FD",
    x"2BB3F27D",
    x"2BB3DC00",
    x"2BB3C586",
    x"2BB3AF0F",
    x"2BB3989A",
    x"2BB38229",
    x"2BB36BBA",
    x"2BB3554E",
    x"2BB33EE4",
    x"2BB3287E",
    x"2BB3121A",
    x"2BB2FBB9",
    x"2BB2E55B",
    x"2BB2CF00",
    x"2BB2B8A8",
    x"2BB2A252",
    x"2BB28BFF",
    x"2BB275AF",
    x"2BB25F62",
    x"2BB24917",
    x"2BB232CF",
    x"2BB21C8A",
    x"2BB20648",
    x"2BB1F009",
    x"2BB1D9CC",
    x"2BB1C392",
    x"2BB1AD5B",
    x"2BB19727",
    x"2BB180F5",
    x"2BB16AC7",
    x"2BB1549B",
    x"2BB13E72",
    x"2BB1284B",
    x"2BB11227",
    x"2BB0FC07",
    x"2BB0E5E8",
    x"2BB0CFCD",
    x"2BB0B9B4",
    x"2BB0A39F",
    x"2BB08D8C",
    x"2BB0777B",
    x"2BB0616E",
    x"2BB04B63",
    x"2BB0355B",
    x"2BB01F56",
    x"2BB00953",
    x"2BAFF353",
    x"2BAFDD56",
    x"2BAFC75C",
    x"2BAFB164",
    x"2BAF9B70",
    x"2BAF857E",
    x"2BAF6F8E",
    x"2BAF59A2",
    x"2BAF43B8",
    x"2BAF2DD1",
    x"2BAF17EC",
    x"2BAF020B",
    x"2BAEEC2C",
    x"2BAED650",
    x"2BAEC076",
    x"2BAEAAA0",
    x"2BAE94CC",
    x"2BAE7EFA",
    x"2BAE692C",
    x"2BAE5360",
    x"2BAE3D97",
    x"2BAE27D1",
    x"2BAE120D",
    x"2BADFC4C",
    x"2BADE68E",
    x"2BADD0D2",
    x"2BADBB1A",
    x"2BADA564",
    x"2BAD8FB0",
    x"2BAD7A00",
    x"2BAD6452",
    x"2BAD4EA7",
    x"2BAD38FE",
    x"2BAD2358",
    x"2BAD0DB5",
    x"2BACF815",
    x"2BACE277",
    x"2BACCCDC",
    x"2BACB744",
    x"2BACA1AF",
    x"2BAC8C1C",
    x"2BAC768C",
    x"2BAC60FE",
    x"2BAC4B73",
    x"2BAC35EB",
    x"2BAC2066",
    x"2BAC0AE3",
    x"2BABF563",
    x"2BABDFE6",
    x"2BABCA6B",
    x"2BABB4F3",
    x"2BAB9F7E",
    x"2BAB8A0B",
    x"2BAB749B",
    x"2BAB5F2E",
    x"2BAB49C4",
    x"2BAB345C",
    x"2BAB1EF7",
    x"2BAB0994",
    x"2BAAF434",
    x"2BAADED7",
    x"2BAAC97C",
    x"2BAAB425",
    x"2BAA9ECF",
    x"2BAA897D",
    x"2BAA742D",
    x"2BAA5EE0",
    x"2BAA4995",
    x"2BAA344D",
    x"2BAA1F08",
    x"2BAA09C6",
    x"2BA9F486",
    x"2BA9DF49",
    x"2BA9CA0E",
    x"2BA9B4D6",
    x"2BA99FA1",
    x"2BA98A6E",
    x"2BA9753E",
    x"2BA96011",
    x"2BA94AE6",
    x"2BA935BE",
    x"2BA92099",
    x"2BA90B76",
    x"2BA8F656",
    x"2BA8E138",
    x"2BA8CC1E",
    x"2BA8B705",
    x"2BA8A1F0",
    x"2BA88CDD",
    x"2BA877CD",
    x"2BA862BF",
    x"2BA84DB4",
    x"2BA838AB",
    x"2BA823A6",
    x"2BA80EA3",
    x"2BA7F9A2",
    x"2BA7E4A4",
    x"2BA7CFA9",
    x"2BA7BAB0",
    x"2BA7A5BA",
    x"2BA790C7",
    x"2BA77BD6",
    x"2BA766E8",
    x"2BA751FC",
    x"2BA73D13",
    x"2BA7282D",
    x"2BA71349",
    x"2BA6FE68",
    x"2BA6E98A",
    x"2BA6D4AE",
    x"2BA6BFD5",
    x"2BA6AAFE",
    x"2BA6962A",
    x"2BA68158",
    x"2BA66C89",
    x"2BA657BD",
    x"2BA642F3",
    x"2BA62E2C",
    x"2BA61968",
    x"2BA604A6",
    x"2BA5EFE7",
    x"2BA5DB2A",
    x"2BA5C670",
    x"2BA5B1B8",
    x"2BA59D04",
    x"2BA58851",
    x"2BA573A1",
    x"2BA55EF4",
    x"2BA54A4A",
    x"2BA535A2",
    x"2BA520FC",
    x"2BA50C5A",
    x"2BA4F7B9",
    x"2BA4E31C",
    x"2BA4CE80",
    x"2BA4B9E8",
    x"2BA4A552",
    x"2BA490BF",
    x"2BA47C2E",
    x"2BA467A0",
    x"2BA45314",
    x"2BA43E8B",
    x"2BA42A04",
    x"2BA41580",
    x"2BA400FF",
    x"2BA3EC80",
    x"2BA3D804",
    x"2BA3C38A",
    x"2BA3AF13",
    x"2BA39A9E",
    x"2BA3862C",
    x"2BA371BD",
    x"2BA35D50",
    x"2BA348E5",
    x"2BA3347E",
    x"2BA32018",
    x"2BA30BB6",
    x"2BA2F755",
    x"2BA2E2F8",
    x"2BA2CE9D",
    x"2BA2BA44",
    x"2BA2A5EE",
    x"2BA2919B",
    x"2BA27D4A",
    x"2BA268FB",
    x"2BA254AF",
    x"2BA24066",
    x"2BA22C1F",
    x"2BA217DB",
    x"2BA20399",
    x"2BA1EF5A",
    x"2BA1DB1D",
    x"2BA1C6E3",
    x"2BA1B2AC",
    x"2BA19E77",
    x"2BA18A44",
    x"2BA17614",
    x"2BA161E7",
    x"2BA14DBC",
    x"2BA13993",
    x"2BA1256D",
    x"2BA1114A",
    x"2BA0FD29",
    x"2BA0E90B",
    x"2BA0D4EF",
    x"2BA0C0D5",
    x"2BA0ACBE",
    x"2BA098AA",
    x"2BA08498",
    x"2BA07089",
    x"2BA05C7C",
    x"2BA04872",
    x"2BA0346A",
    x"2BA02065",
    x"2BA00C62",
    x"2B9FF862",
    x"2B9FE464",
    x"2B9FD069",
    x"2B9FBC70",
    x"2B9FA879",
    x"2B9F9486",
    x"2B9F8094",
    x"2B9F6CA5",
    x"2B9F58B9",
    x"2B9F44CF",
    x"2B9F30E8",
    x"2B9F1D03",
    x"2B9F0921",
    x"2B9EF541",
    x"2B9EE163",
    x"2B9ECD88",
    x"2B9EB9B0",
    x"2B9EA5DA",
    x"2B9E9207",
    x"2B9E7E36",
    x"2B9E6A67",
    x"2B9E569B",
    x"2B9E42D1",
    x"2B9E2F0A",
    x"2B9E1B46",
    x"2B9E0783",
    x"2B9DF3C4",
    x"2B9DE006",
    x"2B9DCC4C",
    x"2B9DB893",
    x"2B9DA4DE",
    x"2B9D912A",
    x"2B9D7D79",
    x"2B9D69CB",
    x"2B9D561F",
    x"2B9D4275",
    x"2B9D2ECE",
    x"2B9D1B2A",
    x"2B9D0787",
    x"2B9CF3E8",
    x"2B9CE04A",
    x"2B9CCCB0",
    x"2B9CB917",
    x"2B9CA581",
    x"2B9C91EE",
    x"2B9C7E5D",
    x"2B9C6ACE",
    x"2B9C5742",
    x"2B9C43B8",
    x"2B9C3031",
    x"2B9C1CAC",
    x"2B9C092A",
    x"2B9BF5AA",
    x"2B9BE22D",
    x"2B9BCEB2",
    x"2B9BBB39",
    x"2B9BA7C3",
    x"2B9B944F",
    x"2B9B80DE",
    x"2B9B6D6F",
    x"2B9B5A02",
    x"2B9B4698",
    x"2B9B3331",
    x"2B9B1FCC",
    x"2B9B0C69",
    x"2B9AF908",
    x"2B9AE5AA",
    x"2B9AD24F",
    x"2B9ABEF6",
    x"2B9AAB9F",
    x"2B9A984B",
    x"2B9A84F9",
    x"2B9A71AA",
    x"2B9A5E5D",
    x"2B9A4B12",
    x"2B9A37CA",
    x"2B9A2484",
    x"2B9A1141",
    x"2B99FE00",
    x"2B99EAC1",
    x"2B99D785",
    x"2B99C44B",
    x"2B99B114",
    x"2B999DDF",
    x"2B998AAD",
    x"2B99777D",
    x"2B99644F",
    x"2B995123",
    x"2B993DFB",
    x"2B992AD4",
    x"2B9917B0",
    x"2B99048E",
    x"2B98F16F",
    x"2B98DE52",
    x"2B98CB37",
    x"2B98B81F",
    x"2B98A509",
    x"2B9891F6",
    x"2B987EE5",
    x"2B986BD6",
    x"2B9858CA",
    x"2B9845C0",
    x"2B9832B8",
    x"2B981FB3",
    x"2B980CB0",
    x"2B97F9B0",
    x"2B97E6B2",
    x"2B97D3B6",
    x"2B97C0BD",
    x"2B97ADC6",
    x"2B979AD1",
    x"2B9787DF",
    x"2B9774EF",
    x"2B976202",
    x"2B974F17",
    x"2B973C2E",
    x"2B972948",
    x"2B971664",
    x"2B970382",
    x"2B96F0A3",
    x"2B96DDC6",
    x"2B96CAEC",
    x"2B96B813",
    x"2B96A53E",
    x"2B96926A",
    x"2B967F99",
    x"2B966CCA",
    x"2B9659FE",
    x"2B964734",
    x"2B96346C",
    x"2B9621A7",
    x"2B960EE4",
    x"2B95FC23",
    x"2B95E965",
    x"2B95D6A9",
    x"2B95C3EF",
    x"2B95B138",
    x"2B959E83",
    x"2B958BD0",
    x"2B957920",
    x"2B956672",
    x"2B9553C6",
    x"2B95411D",
    x"2B952E76",
    x"2B951BD1",
    x"2B95092F",
    x"2B94F68F",
    x"2B94E3F1",
    x"2B94D156",
    x"2B94BEBD",
    x"2B94AC26",
    x"2B949992",
    x"2B948700",
    x"2B947470",
    x"2B9461E3",
    x"2B944F58",
    x"2B943CCF",
    x"2B942A48",
    x"2B9417C4",
    x"2B940542",
    x"2B93F2C3",
    x"2B93E046",
    x"2B93CDCB",
    x"2B93BB52",
    x"2B93A8DC",
    x"2B939668",
    x"2B9383F6",
    x"2B937187",
    x"2B935F1A",
    x"2B934CAF",
    x"2B933A47",
    x"2B9327E1",
    x"2B93157D",
    x"2B93031B",
    x"2B92F0BC",
    x"2B92DE5F",
    x"2B92CC05",
    x"2B92B9AC",
    x"2B92A756",
    x"2B929502",
    x"2B9282B1",
    x"2B927062",
    x"2B925E15",
    x"2B924BCA",
    x"2B923982",
    x"2B92273C",
    x"2B9214F8",
    x"2B9202B7",
    x"2B91F077",
    x"2B91DE3A",
    x"2B91CC00",
    x"2B91B9C7",
    x"2B91A791",
    x"2B91955E",
    x"2B91832C",
    x"2B9170FD",
    x"2B915ED0",
    x"2B914CA5",
    x"2B913A7D",
    x"2B912856",
    x"2B911632",
    x"2B910411",
    x"2B90F1F1",
    x"2B90DFD4",
    x"2B90CDBA",
    x"2B90BBA1",
    x"2B90A98B",
    x"2B909777",
    x"2B908565",
    x"2B907355",
    x"2B906148",
    x"2B904F3D",
    x"2B903D34",
    x"2B902B2E",
    x"2B901929",
    x"2B900727",
    x"2B8FF528",
    x"2B8FE32A",
    x"2B8FD12F",
    x"2B8FBF36",
    x"2B8FAD3F",
    x"2B8F9B4A",
    x"2B8F8958",
    x"2B8F7768",
    x"2B8F657A",
    x"2B8F538F",
    x"2B8F41A5",
    x"2B8F2FBE",
    x"2B8F1DD9",
    x"2B8F0BF7",
    x"2B8EFA16",
    x"2B8EE838",
    x"2B8ED65C",
    x"2B8EC483",
    x"2B8EB2AB",
    x"2B8EA0D6",
    x"2B8E8F03",
    x"2B8E7D32",
    x"2B8E6B64",
    x"2B8E5997",
    x"2B8E47CD",
    x"2B8E3605",
    x"2B8E2440",
    x"2B8E127C",
    x"2B8E00BB",
    x"2B8DEEFC",
    x"2B8DDD3F",
    x"2B8DCB85",
    x"2B8DB9CD",
    x"2B8DA816",
    x"2B8D9663",
    x"2B8D84B1",
    x"2B8D7301",
    x"2B8D6154",
    x"2B8D4FA9",
    x"2B8D3E00",
    x"2B8D2C5A",
    x"2B8D1AB5",
    x"2B8D0913",
    x"2B8CF773",
    x"2B8CE5D5",
    x"2B8CD439",
    x"2B8CC2A0",
    x"2B8CB109",
    x"2B8C9F74",
    x"2B8C8DE1",
    x"2B8C7C50",
    x"2B8C6AC2",
    x"2B8C5936",
    x"2B8C47AB",
    x"2B8C3624",
    x"2B8C249E",
    x"2B8C131A",
    x"2B8C0199",
    x"2B8BF01A",
    x"2B8BDE9D",
    x"2B8BCD22",
    x"2B8BBBAA",
    x"2B8BAA33",
    x"2B8B98BF",
    x"2B8B874D",
    x"2B8B75DD",
    x"2B8B6470",
    x"2B8B5304",
    x"2B8B419B",
    x"2B8B3034",
    x"2B8B1ECF",
    x"2B8B0D6C",
    x"2B8AFC0C",
    x"2B8AEAAD",
    x"2B8AD951",
    x"2B8AC7F7",
    x"2B8AB69F",
    x"2B8AA549",
    x"2B8A93F6",
    x"2B8A82A4",
    x"2B8A7155",
    x"2B8A6008",
    x"2B8A4EBD",
    x"2B8A3D74",
    x"2B8A2C2E",
    x"2B8A1AE9",
    x"2B8A09A7",
    x"2B89F867",
    x"2B89E729",
    x"2B89D5ED",
    x"2B89C4B3",
    x"2B89B37C",
    x"2B89A246",
    x"2B899113",
    x"2B897FE2",
    x"2B896EB3",
    x"2B895D87",
    x"2B894C5C",
    x"2B893B33",
    x"2B892A0D",
    x"2B8918E9",
    x"2B8907C7",
    x"2B88F6A7",
    x"2B88E589",
    x"2B88D46E",
    x"2B88C354",
    x"2B88B23D",
    x"2B88A128",
    x"2B889014",
    x"2B887F04",
    x"2B886DF5",
    x"2B885CE8",
    x"2B884BDE",
    x"2B883AD5",
    x"2B8829CF",
    x"2B8818CB",
    x"2B8807C9",
    x"2B87F6C9",
    x"2B87E5CB",
    x"2B87D4CF",
    x"2B87C3D6",
    x"2B87B2DE",
    x"2B87A1E9",
    x"2B8790F6",
    x"2B878005",
    x"2B876F16",
    x"2B875E29",
    x"2B874D3E",
    x"2B873C56",
    x"2B872B6F",
    x"2B871A8B",
    x"2B8709A9",
    x"2B86F8C8",
    x"2B86E7EA",
    x"2B86D70E",
    x"2B86C635",
    x"2B86B55D",
    x"2B86A487",
    x"2B8693B4",
    x"2B8682E2",
    x"2B867213",
    x"2B866146",
    x"2B86507B",
    x"2B863FB2",
    x"2B862EEB",
    x"2B861E26",
    x"2B860D63",
    x"2B85FCA3",
    x"2B85EBE4",
    x"2B85DB28",
    x"2B85CA6D",
    x"2B85B9B5",
    x"2B85A8FF",
    x"2B85984B",
    x"2B858799",
    x"2B8576E9",
    x"2B85663B",
    x"2B85558F",
    x"2B8544E6",
    x"2B85343E",
    x"2B852399",
    x"2B8512F5",
    x"2B850254",
    x"2B84F1B5",
    x"2B84E117",
    x"2B84D07C",
    x"2B84BFE3",
    x"2B84AF4C",
    x"2B849EB7",
    x"2B848E25",
    x"2B847D94",
    x"2B846D05",
    x"2B845C79",
    x"2B844BEE",
    x"2B843B66",
    x"2B842ADF",
    x"2B841A5B",
    x"2B8409D9",
    x"2B83F959",
    x"2B83E8DA",
    x"2B83D85E",
    x"2B83C7E4",
    x"2B83B76C",
    x"2B83A6F6",
    x"2B839683",
    x"2B838611",
    x"2B8375A1",
    x"2B836533",
    x"2B8354C8",
    x"2B83445E",
    x"2B8333F7",
    x"2B832391",
    x"2B83132E",
    x"2B8302CC",
    x"2B82F26D",
    x"2B82E210",
    x"2B82D1B5",
    x"2B82C15B",
    x"2B82B104",
    x"2B82A0AF",
    x"2B82905C",
    x"2B82800B",
    x"2B826FBC",
    x"2B825F6F",
    x"2B824F24",
    x"2B823EDB",
    x"2B822E94",
    x"2B821E50",
    x"2B820E0D",
    x"2B81FDCC",
    x"2B81ED8D",
    x"2B81DD51",
    x"2B81CD16",
    x"2B81BCDE",
    x"2B81ACA7",
    x"2B819C72",
    x"2B818C40",
    x"2B817C0F",
    x"2B816BE1",
    x"2B815BB4",
    x"2B814B8A",
    x"2B813B61",
    x"2B812B3B",
    x"2B811B17",
    x"2B810AF4",
    x"2B80FAD4",
    x"2B80EAB6",
    x"2B80DA99",
    x"2B80CA7F",
    x"2B80BA67",
    x"2B80AA50",
    x"2B809A3C",
    x"2B808A2A",
    x"2B807A19",
    x"2B806A0B",
    x"2B8059FF",
    x"2B8049F5",
    x"2B8039EC",
    x"2B8029E6",
    x"2B8019E2",
    x"2B8009E0",
    x"2B7FF3BF",
    x"2B7FD3C3",
    x"2B7FB3CA",
    x"2B7F93D6",
    x"2B7F73E5",
    x"2B7F53F9",
    x"2B7F3410",
    x"2B7F142C",
    x"2B7EF44B",
    x"2B7ED46F",
    x"2B7EB496",
    x"2B7E94C1",
    x"2B7E74F1",
    x"2B7E5524",
    x"2B7E355B",
    x"2B7E1597",
    x"2B7DF5D6",
    x"2B7DD619",
    x"2B7DB661",
    x"2B7D96AC",
    x"2B7D76FB",
    x"2B7D574E",
    x"2B7D37A5",
    x"2B7D1800",
    x"2B7CF85F",
    x"2B7CD8C2",
    x"2B7CB929",
    x"2B7C9994",
    x"2B7C7A02",
    x"2B7C5A75",
    x"2B7C3AEC",
    x"2B7C1B66",
    x"2B7BFBE5",
    x"2B7BDC68",
    x"2B7BBCEE",
    x"2B7B9D78",
    x"2B7B7E07",
    x"2B7B5E99",
    x"2B7B3F2F",
    x"2B7B1FC9",
    x"2B7B0067",
    x"2B7AE109",
    x"2B7AC1AF",
    x"2B7AA258",
    x"2B7A8306",
    x"2B7A63B8",
    x"2B7A446D",
    x"2B7A2527",
    x"2B7A05E4",
    x"2B79E6A5",
    x"2B79C76A",
    x"2B79A833",
    x"2B798900",
    x"2B7969D1",
    x"2B794AA6",
    x"2B792B7E",
    x"2B790C5B",
    x"2B78ED3B",
    x"2B78CE20",
    x"2B78AF08",
    x"2B788FF4",
    x"2B7870E4",
    x"2B7851D8",
    x"2B7832CF",
    x"2B7813CB",
    x"2B77F4CA",
    x"2B77D5CE",
    x"2B77B6D5",
    x"2B7797E0",
    x"2B7778EF",
    x"2B775A02",
    x"2B773B18",
    x"2B771C33",
    x"2B76FD51",
    x"2B76DE74",
    x"2B76BF9A",
    x"2B76A0C4",
    x"2B7681F2",
    x"2B766323",
    x"2B764459",
    x"2B762592",
    x"2B7606CF",
    x"2B75E810",
    x"2B75C955",
    x"2B75AA9E",
    x"2B758BEB",
    x"2B756D3B",
    x"2B754E8F",
    x"2B752FE7",
    x"2B751143",
    x"2B74F2A3",
    x"2B74D407",
    x"2B74B56E",
    x"2B7496D9",
    x"2B747848",
    x"2B7459BB",
    x"2B743B32",
    x"2B741CAD",
    x"2B73FE2B",
    x"2B73DFAD",
    x"2B73C133",
    x"2B73A2BD",
    x"2B73844A",
    x"2B7365DC",
    x"2B734771",
    x"2B73290A",
    x"2B730AA7",
    x"2B72EC47",
    x"2B72CDEB",
    x"2B72AF94",
    x"2B729140",
    x"2B7272EF",
    x"2B7254A3",
    x"2B72365A",
    x"2B721815",
    x"2B71F9D4",
    x"2B71DB97",
    x"2B71BD5D",
    x"2B719F27",
    x"2B7180F5",
    x"2B7162C7",
    x"2B71449D",
    x"2B712676",
    x"2B710853",
    x"2B70EA34",
    x"2B70CC19",
    x"2B70AE01",
    x"2B708FED",
    x"2B7071DD",
    x"2B7053D1",
    x"2B7035C8",
    x"2B7017C3",
    x"2B6FF9C2",
    x"2B6FDBC5",
    x"2B6FBDCB",
    x"2B6F9FD5",
    x"2B6F81E3",
    x"2B6F63F5",
    x"2B6F460A",
    x"2B6F2823",
    x"2B6F0A40",
    x"2B6EEC61",
    x"2B6ECE85",
    x"2B6EB0AD",
    x"2B6E92D9",
    x"2B6E7508",
    x"2B6E573C",
    x"2B6E3973",
    x"2B6E1BAD",
    x"2B6DFDEC",
    x"2B6DE02E",
    x"2B6DC274",
    x"2B6DA4BD",
    x"2B6D870A",
    x"2B6D695B",
    x"2B6D4BB0",
    x"2B6D2E08",
    x"2B6D1065",
    x"2B6CF2C4",
    x"2B6CD528",
    x"2B6CB78F",
    x"2B6C99FA",
    x"2B6C7C69",
    x"2B6C5EDB",
    x"2B6C4151",
    x"2B6C23CB",
    x"2B6C0648",
    x"2B6BE8C9",
    x"2B6BCB4E",
    x"2B6BADD6",
    x"2B6B9062",
    x"2B6B72F2",
    x"2B6B5586",
    x"2B6B381D",
    x"2B6B1AB7",
    x"2B6AFD56",
    x"2B6ADFF8",
    x"2B6AC29E",
    x"2B6AA548",
    x"2B6A87F5",
    x"2B6A6AA6",
    x"2B6A4D5A",
    x"2B6A3012",
    x"2B6A12CE",
    x"2B69F58D",
    x"2B69D851",
    x"2B69BB17",
    x"2B699DE2",
    x"2B6980B0",
    x"2B696382",
    x"2B694657",
    x"2B692930",
    x"2B690C0D",
    x"2B68EEED",
    x"2B68D1D1",
    x"2B68B4B9",
    x"2B6897A4",
    x"2B687A93",
    x"2B685D85",
    x"2B68407B",
    x"2B682375",
    x"2B680672",
    x"2B67E973",
    x"2B67CC78",
    x"2B67AF80",
    x"2B67928C",
    x"2B67759C",
    x"2B6758AF",
    x"2B673BC6",
    x"2B671EE0",
    x"2B6701FE",
    x"2B66E51F",
    x"2B66C845",
    x"2B66AB6D",
    x"2B668E9A",
    x"2B6671CA",
    x"2B6654FD",
    x"2B663834",
    x"2B661B6F",
    x"2B65FEAE",
    x"2B65E1F0",
    x"2B65C535",
    x"2B65A87E",
    x"2B658BCB",
    x"2B656F1B",
    x"2B65526F",
    x"2B6535C7",
    x"2B651922",
    x"2B64FC80",
    x"2B64DFE3",
    x"2B64C348",
    x"2B64A6B2",
    x"2B648A1F",
    x"2B646D8F",
    x"2B645103",
    x"2B64347B",
    x"2B6417F6",
    x"2B63FB75",
    x"2B63DEF7",
    x"2B63C27D",
    x"2B63A607",
    x"2B638994",
    x"2B636D24",
    x"2B6350B8",
    x"2B633450",
    x"2B6317EB",
    x"2B62FB8A",
    x"2B62DF2C",
    x"2B62C2D2",
    x"2B62A67C",
    x"2B628A29",
    x"2B626DD9",
    x"2B62518D",
    x"2B623545",
    x"2B621900",
    x"2B61FCBF",
    x"2B61E081",
    x"2B61C446",
    x"2B61A810",
    x"2B618BDC",
    x"2B616FAD",
    x"2B615381",
    x"2B613758",
    x"2B611B33",
    x"2B60FF11",
    x"2B60E2F3",
    x"2B60C6D8",
    x"2B60AAC1",
    x"2B608EAE",
    x"2B60729E",
    x"2B605691",
    x"2B603A88",
    x"2B601E82",
    x"2B600280",
    x"2B5FE682",
    x"2B5FCA87",
    x"2B5FAE8F",
    x"2B5F929B",
    x"2B5F76AA",
    x"2B5F5ABD",
    x"2B5F3ED4",
    x"2B5F22EE",
    x"2B5F070B",
    x"2B5EEB2C",
    x"2B5ECF50",
    x"2B5EB378",
    x"2B5E97A3",
    x"2B5E7BD2",
    x"2B5E6004",
    x"2B5E443A",
    x"2B5E2873",
    x"2B5E0CB0",
    x"2B5DF0F0",
    x"2B5DD534",
    x"2B5DB97B",
    x"2B5D9DC5",
    x"2B5D8213",
    x"2B5D6665",
    x"2B5D4ABA",
    x"2B5D2F12",
    x"2B5D136E",
    x"2B5CF7CD",
    x"2B5CDC30",
    x"2B5CC096",
    x"2B5CA500",
    x"2B5C896D",
    x"2B5C6DDE",
    x"2B5C5252",
    x"2B5C36C9",
    x"2B5C1B44",
    x"2B5BFFC2",
    x"2B5BE444",
    x"2B5BC8C9",
    x"2B5BAD52",
    x"2B5B91DE",
    x"2B5B766D",
    x"2B5B5B00",
    x"2B5B3F97",
    x"2B5B2430",
    x"2B5B08CD",
    x"2B5AED6E",
    x"2B5AD212",
    x"2B5AB6BA",
    x"2B5A9B64",
    x"2B5A8013",
    x"2B5A64C4",
    x"2B5A497A",
    x"2B5A2E32",
    x"2B5A12EE",
    x"2B59F7AD",
    x"2B59DC70",
    x"2B59C136",
    x"2B59A600",
    x"2B598ACD",
    x"2B596F9D",
    x"2B595471",
    x"2B593948",
    x"2B591E22",
    x"2B590300",
    x"2B58E7E2",
    x"2B58CCC6",
    x"2B58B1AF",
    x"2B58969A",
    x"2B587B89",
    x"2B58607B",
    x"2B584571",
    x"2B582A6A",
    x"2B580F66",
    x"2B57F466",
    x"2B57D969",
    x"2B57BE70",
    x"2B57A379",
    x"2B578887",
    x"2B576D97",
    x"2B5752AB",
    x"2B5737C3",
    x"2B571CDD",
    x"2B5701FB",
    x"2B56E71D",
    x"2B56CC42",
    x"2B56B16A",
    x"2B569695",
    x"2B567BC4",
    x"2B5660F6",
    x"2B56462C",
    x"2B562B65",
    x"2B5610A1",
    x"2B55F5E1",
    x"2B55DB24",
    x"2B55C06A",
    x"2B55A5B4",
    x"2B558B00",
    x"2B557051",
    x"2B5555A4",
    x"2B553AFB",
    x"2B552056",
    x"2B5505B3",
    x"2B54EB14",
    x"2B54D078",
    x"2B54B5E0",
    x"2B549B4B",
    x"2B5480B9",
    x"2B54662B",
    x"2B544BA0",
    x"2B543118",
    x"2B541693",
    x"2B53FC12",
    x"2B53E194",
    x"2B53C71A",
    x"2B53ACA3",
    x"2B53922F",
    x"2B5377BE",
    x"2B535D51",
    x"2B5342E7",
    x"2B532880",
    x"2B530E1D",
    x"2B52F3BD",
    x"2B52D960",
    x"2B52BF06",
    x"2B52A4B0",
    x"2B528A5D",
    x"2B52700D",
    x"2B5255C1",
    x"2B523B78",
    x"2B522132",
    x"2B5206F0",
    x"2B51ECB0",
    x"2B51D274",
    x"2B51B83C",
    x"2B519E06",
    x"2B5183D4",
    x"2B5169A5",
    x"2B514F7A",
    x"2B513552",
    x"2B511B2D",
    x"2B51010B",
    x"2B50E6EC",
    x"2B50CCD1",
    x"2B50B2B9",
    x"2B5098A4",
    x"2B507E93",
    x"2B506485",
    x"2B504A7A",
    x"2B503072",
    x"2B50166E",
    x"2B4FFC6D",
    x"2B4FE26F",
    x"2B4FC874",
    x"2B4FAE7C",
    x"2B4F9488",
    x"2B4F7A97",
    x"2B4F60AA",
    x"2B4F46BF",
    x"2B4F2CD8",
    x"2B4F12F4",
    x"2B4EF913",
    x"2B4EDF36",
    x"2B4EC55B",
    x"2B4EAB84",
    x"2B4E91B1",
    x"2B4E77E0",
    x"2B4E5E13",
    x"2B4E4448",
    x"2B4E2A81",
    x"2B4E10BE",
    x"2B4DF6FD",
    x"2B4DDD40",
    x"2B4DC386",
    x"2B4DA9CF",
    x"2B4D901C",
    x"2B4D766B",
    x"2B4D5CBE",
    x"2B4D4314",
    x"2B4D296D",
    x"2B4D0FCA",
    x"2B4CF629",
    x"2B4CDC8C",
    x"2B4CC2F2",
    x"2B4CA95B",
    x"2B4C8FC8",
    x"2B4C7637",
    x"2B4C5CAA",
    x"2B4C4320",
    x"2B4C2999",
    x"2B4C1016",
    x"2B4BF695",
    x"2B4BDD18",
    x"2B4BC39E",
    x"2B4BAA27",
    x"2B4B90B4",
    x"2B4B7743",
    x"2B4B5DD6",
    x"2B4B446C",
    x"2B4B2B05",
    x"2B4B11A1",
    x"2B4AF840",
    x"2B4ADEE3",
    x"2B4AC589",
    x"2B4AAC31",
    x"2B4A92DD",
    x"2B4A798D",
    x"2B4A603F",
    x"2B4A46F5",
    x"2B4A2DAD",
    x"2B4A1469",
    x"2B49FB28",
    x"2B49E1EA",
    x"2B49C8B0",
    x"2B49AF78",
    x"2B499644",
    x"2B497D13",
    x"2B4963E5",
    x"2B494ABA",
    x"2B493192",
    x"2B49186D",
    x"2B48FF4C",
    x"2B48E62D",
    x"2B48CD12",
    x"2B48B3FA",
    x"2B489AE5",
    x"2B4881D3",
    x"2B4868C5",
    x"2B484FB9",
    x"2B4836B1",
    x"2B481DAC",
    x"2B4804A9",
    x"2B47EBAA",
    x"2B47D2AF",
    x"2B47B9B6",
    x"2B47A0C0",
    x"2B4787CE",
    x"2B476EDE",
    x"2B4755F2",
    x"2B473D09",
    x"2B472423",
    x"2B470B40",
    x"2B46F260",
    x"2B46D983",
    x"2B46C0A9",
    x"2B46A7D3",
    x"2B468EFF",
    x"2B46762F",
    x"2B465D62",
    x"2B464498",
    x"2B462BD1",
    x"2B46130D",
    x"2B45FA4C",
    x"2B45E18E",
    x"2B45C8D4",
    x"2B45B01C",
    x"2B459768",
    x"2B457EB6",
    x"2B456608",
    x"2B454D5D",
    x"2B4534B5",
    x"2B451C10",
    x"2B45036E",
    x"2B44EACF",
    x"2B44D233",
    x"2B44B99A",
    x"2B44A104",
    x"2B448872",
    x"2B446FE2",
    x"2B445756",
    x"2B443ECD",
    x"2B442646",
    x"2B440DC3",
    x"2B43F543",
    x"2B43DCC6",
    x"2B43C44C",
    x"2B43ABD5",
    x"2B439361",
    x"2B437AF0",
    x"2B436282",
    x"2B434A17",
    x"2B4331AF",
    x"2B43194B",
    x"2B4300E9",
    x"2B42E88A",
    x"2B42D02F",
    x"2B42B7D6",
    x"2B429F81",
    x"2B42872F",
    x"2B426EDF",
    x"2B425693",
    x"2B423E49",
    x"2B422603",
    x"2B420DC0",
    x"2B41F580",
    x"2B41DD43",
    x"2B41C508",
    x"2B41ACD1",
    x"2B41949D",
    x"2B417C6C",
    x"2B41643E",
    x"2B414C13",
    x"2B4133EB",
    x"2B411BC6",
    x"2B4103A4",
    x"2B40EB85",
    x"2B40D369",
    x"2B40BB50",
    x"2B40A33A",
    x"2B408B28",
    x"2B407318",
    x"2B405B0B",
    x"2B404301",
    x"2B402AFA",
    x"2B4012F6",
    x"2B3FFAF5",
    x"2B3FE2F7",
    x"2B3FCAFD",
    x"2B3FB305",
    x"2B3F9B10",
    x"2B3F831E",
    x"2B3F6B2F",
    x"2B3F5343",
    x"2B3F3B5A",
    x"2B3F2374",
    x"2B3F0B91",
    x"2B3EF3B1",
    x"2B3EDBD4",
    x"2B3EC3FA",
    x"2B3EAC23",
    x"2B3E944F",
    x"2B3E7C7E",
    x"2B3E64B0",
    x"2B3E4CE5",
    x"2B3E351D",
    x"2B3E1D58",
    x"2B3E0596",
    x"2B3DEDD7",
    x"2B3DD61A",
    x"2B3DBE61",
    x"2B3DA6AB",
    x"2B3D8EF7",
    x"2B3D7747",
    x"2B3D5F99",
    x"2B3D47EF",
    x"2B3D3048",
    x"2B3D18A3",
    x"2B3D0101",
    x"2B3CE963",
    x"2B3CD1C7",
    x"2B3CBA2E",
    x"2B3CA298",
    x"2B3C8B06",
    x"2B3C7376",
    x"2B3C5BE9",
    x"2B3C445F",
    x"2B3C2CD8",
    x"2B3C1554",
    x"2B3BFDD2",
    x"2B3BE654",
    x"2B3BCED9",
    x"2B3BB760",
    x"2B3B9FEB",
    x"2B3B8878",
    x"2B3B7109",
    x"2B3B599C",
    x"2B3B4232",
    x"2B3B2ACC",
    x"2B3B1368",
    x"2B3AFC07",
    x"2B3AE4A9",
    x"2B3ACD4E",
    x"2B3AB5F5",
    x"2B3A9EA0",
    x"2B3A874E",
    x"2B3A6FFE",
    x"2B3A58B2",
    x"2B3A4168",
    x"2B3A2A21",
    x"2B3A12DE",
    x"2B39FB9D",
    x"2B39E45F",
    x"2B39CD24",
    x"2B39B5EB",
    x"2B399EB6",
    x"2B398784",
    x"2B397054",
    x"2B395928",
    x"2B3941FE",
    x"2B392AD7",
    x"2B3913B3",
    x"2B38FC92",
    x"2B38E574",
    x"2B38CE59",
    x"2B38B740",
    x"2B38A02B",
    x"2B388918",
    x"2B387209",
    x"2B385AFC",
    x"2B3843F2",
    x"2B382CEB",
    x"2B3815E7",
    x"2B37FEE5",
    x"2B37E7E7",
    x"2B37D0EB",
    x"2B37B9F3",
    x"2B37A2FD",
    x"2B378C0A",
    x"2B37751A",
    x"2B375E2D",
    x"2B374742",
    x"2B37305B",
    x"2B371976",
    x"2B370295",
    x"2B36EBB6",
    x"2B36D4DA",
    x"2B36BE00",
    x"2B36A72A",
    x"2B369057",
    x"2B367986",
    x"2B3662B8",
    x"2B364BED",
    x"2B363525",
    x"2B361E60",
    x"2B36079E",
    x"2B35F0DE",
    x"2B35DA21",
    x"2B35C368",
    x"2B35ACB1",
    x"2B3595FC",
    x"2B357F4B",
    x"2B35689D",
    x"2B3551F1",
    x"2B353B48",
    x"2B3524A2",
    x"2B350DFF",
    x"2B34F75F",
    x"2B34E0C1",
    x"2B34CA26",
    x"2B34B38F",
    x"2B349CFA",
    x"2B348667",
    x"2B346FD8",
    x"2B34594B",
    x"2B3442C2",
    x"2B342C3B",
    x"2B3415B7",
    x"2B33FF35",
    x"2B33E8B7",
    x"2B33D23B",
    x"2B33BBC2",
    x"2B33A54C",
    x"2B338ED9",
    x"2B337868",
    x"2B3361FB",
    x"2B334B90",
    x"2B333528",
    x"2B331EC3",
    x"2B330860",
    x"2B32F201",
    x"2B32DBA4",
    x"2B32C54A",
    x"2B32AEF2",
    x"2B32989E",
    x"2B32824C",
    x"2B326BFD",
    x"2B3255B1",
    x"2B323F68",
    x"2B322921",
    x"2B3212DE",
    x"2B31FC9D",
    x"2B31E65E",
    x"2B31D023",
    x"2B31B9EA",
    x"2B31A3B5",
    x"2B318D82",
    x"2B317751",
    x"2B316124",
    x"2B314AF9",
    x"2B3134D1",
    x"2B311EAC",
    x"2B310889",
    x"2B30F26A",
    x"2B30DC4D",
    x"2B30C633",
    x"2B30B01B",
    x"2B309A07",
    x"2B3083F5",
    x"2B306DE6",
    x"2B3057D9",
    x"2B3041D0",
    x"2B302BC9",
    x"2B3015C5",
    x"2B2FFFC3",
    x"2B2FE9C5",
    x"2B2FD3C9",
    x"2B2FBDD0",
    x"2B2FA7D9",
    x"2B2F91E6",
    x"2B2F7BF5",
    x"2B2F6607",
    x"2B2F501B",
    x"2B2F3A33",
    x"2B2F244D",
    x"2B2F0E6A",
    x"2B2EF889",
    x"2B2EE2AC",
    x"2B2ECCD1",
    x"2B2EB6F8",
    x"2B2EA123",
    x"2B2E8B50",
    x"2B2E7580",
    x"2B2E5FB3",
    x"2B2E49E8",
    x"2B2E3420",
    x"2B2E1E5B",
    x"2B2E0899",
    x"2B2DF2D9",
    x"2B2DDD1C",
    x"2B2DC762",
    x"2B2DB1AA",
    x"2B2D9BF5",
    x"2B2D8643",
    x"2B2D7094",
    x"2B2D5AE7",
    x"2B2D453D",
    x"2B2D2F96",
    x"2B2D19F1",
    x"2B2D044F",
    x"2B2CEEB0",
    x"2B2CD913",
    x"2B2CC37A",
    x"2B2CADE3",
    x"2B2C984E",
    x"2B2C82BC",
    x"2B2C6D2E",
    x"2B2C57A1",
    x"2B2C4218",
    x"2B2C2C91",
    x"2B2C170C",
    x"2B2C018B",
    x"2B2BEC0C",
    x"2B2BD690",
    x"2B2BC116",
    x"2B2BABA0",
    x"2B2B962C",
    x"2B2B80BA",
    x"2B2B6B4B",
    x"2B2B55DF",
    x"2B2B4076",
    x"2B2B2B0F",
    x"2B2B15AB",
    x"2B2B004A",
    x"2B2AEAEB",
    x"2B2AD58F",
    x"2B2AC036",
    x"2B2AAADF",
    x"2B2A958B",
    x"2B2A803A",
    x"2B2A6AEB",
    x"2B2A559F",
    x"2B2A4055",
    x"2B2A2B0F",
    x"2B2A15CB",
    x"2B2A0089",
    x"2B29EB4B",
    x"2B29D60E",
    x"2B29C0D5",
    x"2B29AB9E",
    x"2B29966A",
    x"2B298139",
    x"2B296C0A",
    x"2B2956DE",
    x"2B2941B4",
    x"2B292C8D",
    x"2B291769",
    x"2B290247",
    x"2B28ED28",
    x"2B28D80C",
    x"2B28C2F2",
    x"2B28ADDB",
    x"2B2898C7",
    x"2B2883B5",
    x"2B286EA6",
    x"2B285999",
    x"2B284490",
    x"2B282F88",
    x"2B281A84",
    x"2B280582",
    x"2B27F082",
    x"2B27DB86",
    x"2B27C68B",
    x"2B27B194",
    x"2B279C9F",
    x"2B2787AD",
    x"2B2772BD",
    x"2B275DD0",
    x"2B2748E6",
    x"2B2733FE",
    x"2B271F19",
    x"2B270A36",
    x"2B26F556",
    x"2B26E079",
    x"2B26CB9E",
    x"2B26B6C6",
    x"2B26A1F0",
    x"2B268D1D",
    x"2B26784D",
    x"2B26637F",
    x"2B264EB4",
    x"2B2639EC",
    x"2B262526",
    x"2B261062",
    x"2B25FBA2",
    x"2B25E6E3",
    x"2B25D228",
    x"2B25BD6F",
    x"2B25A8B9",
    x"2B259405",
    x"2B257F54",
    x"2B256AA5",
    x"2B2555F9",
    x"2B25414F",
    x"2B252CA9",
    x"2B251804",
    x"2B250363",
    x"2B24EEC3",
    x"2B24DA27",
    x"2B24C58D",
    x"2B24B0F5",
    x"2B249C61",
    x"2B2487CE",
    x"2B24733F",
    x"2B245EB2",
    x"2B244A27",
    x"2B24359F",
    x"2B24211A",
    x"2B240C97",
    x"2B23F816",
    x"2B23E399",
    x"2B23CF1E",
    x"2B23BAA5",
    x"2B23A62F",
    x"2B2391BB",
    x"2B237D4A",
    x"2B2368DC",
    x"2B235470",
    x"2B234007",
    x"2B232BA0",
    x"2B23173C",
    x"2B2302DA",
    x"2B22EE7B",
    x"2B22DA1F",
    x"2B22C5C5",
    x"2B22B16D",
    x"2B229D18",
    x"2B2288C6",
    x"2B227476",
    x"2B226029",
    x"2B224BDE",
    x"2B223796",
    x"2B222350",
    x"2B220F0D",
    x"2B21FACD",
    x"2B21E68E",
    x"2B21D253",
    x"2B21BE1A",
    x"2B21A9E3",
    x"2B2195AF",
    x"2B21817E",
    x"2B216D4F",
    x"2B215923",
    x"2B2144F9",
    x"2B2130D1",
    x"2B211CAD",
    x"2B21088A",
    x"2B20F46A",
    x"2B20E04D",
    x"2B20CC32",
    x"2B20B81A",
    x"2B20A404",
    x"2B208FF1",
    x"2B207BE0",
    x"2B2067D2",
    x"2B2053C6",
    x"2B203FBD",
    x"2B202BB6",
    x"2B2017B2",
    x"2B2003B0",
    x"2B1FEFB1",
    x"2B1FDBB5",
    x"2B1FC7BA",
    x"2B1FB3C3",
    x"2B1F9FCD",
    x"2B1F8BDB",
    x"2B1F77EA",
    x"2B1F63FD",
    x"2B1F5011",
    x"2B1F3C29",
    x"2B1F2842",
    x"2B1F145F",
    x"2B1F007D",
    x"2B1EEC9F",
    x"2B1ED8C2",
    x"2B1EC4E8",
    x"2B1EB111",
    x"2B1E9D3C",
    x"2B1E896A",
    x"2B1E759A",
    x"2B1E61CC",
    x"2B1E4E01",
    x"2B1E3A39",
    x"2B1E2673",
    x"2B1E12AF",
    x"2B1DFEEE",
    x"2B1DEB2F",
    x"2B1DD773",
    x"2B1DC3BA",
    x"2B1DB002",
    x"2B1D9C4E",
    x"2B1D889B",
    x"2B1D74EB",
    x"2B1D613E",
    x"2B1D4D93",
    x"2B1D39EB",
    x"2B1D2645",
    x"2B1D12A1",
    x"2B1CFF00",
    x"2B1CEB61",
    x"2B1CD7C5",
    x"2B1CC42B",
    x"2B1CB094",
    x"2B1C9CFF",
    x"2B1C896D",
    x"2B1C75DD",
    x"2B1C624F",
    x"2B1C4EC4",
    x"2B1C3B3C",
    x"2B1C27B5",
    x"2B1C1432",
    x"2B1C00B0",
    x"2B1BED32",
    x"2B1BD9B5",
    x"2B1BC63B",
    x"2B1BB2C4",
    x"2B1B9F4E",
    x"2B1B8BDC",
    x"2B1B786B",
    x"2B1B64FE",
    x"2B1B5192",
    x"2B1B3E29",
    x"2B1B2AC3",
    x"2B1B175F",
    x"2B1B03FD",
    x"2B1AF09E",
    x"2B1ADD41",
    x"2B1AC9E6",
    x"2B1AB68E",
    x"2B1AA339",
    x"2B1A8FE5",
    x"2B1A7C95",
    x"2B1A6946",
    x"2B1A55FA",
    x"2B1A42B1",
    x"2B1A2F6A",
    x"2B1A1C25",
    x"2B1A08E3",
    x"2B19F5A3",
    x"2B19E265",
    x"2B19CF2A",
    x"2B19BBF1",
    x"2B19A8BB",
    x"2B199587",
    x"2B198256",
    x"2B196F27",
    x"2B195BFA",
    x"2B1948D0",
    x"2B1935A8",
    x"2B192282",
    x"2B190F5F",
    x"2B18FC3E",
    x"2B18E920",
    x"2B18D604",
    x"2B18C2EB",
    x"2B18AFD3",
    x"2B189CBF",
    x"2B1889AC",
    x"2B18769C",
    x"2B18638E",
    x"2B185083",
    x"2B183D7A",
    x"2B182A74",
    x"2B181770",
    x"2B18046E",
    x"2B17F16F",
    x"2B17DE72",
    x"2B17CB77",
    x"2B17B87F",
    x"2B17A589",
    x"2B179295",
    x"2B177FA4",
    x"2B176CB5",
    x"2B1759C9",
    x"2B1746DF",
    x"2B1733F7",
    x"2B172112",
    x"2B170E2F",
    x"2B16FB4F",
    x"2B16E870",
    x"2B16D594",
    x"2B16C2BB",
    x"2B16AFE4",
    x"2B169D0F",
    x"2B168A3C",
    x"2B16776C",
    x"2B16649F",
    x"2B1651D3",
    x"2B163F0A",
    x"2B162C43",
    x"2B16197F",
    x"2B1606BD",
    x"2B15F3FD",
    x"2B15E140",
    x"2B15CE85",
    x"2B15BBCC",
    x"2B15A916",
    x"2B159662",
    x"2B1583B1",
    x"2B157101",
    x"2B155E54",
    x"2B154BAA",
    x"2B153901",
    x"2B15265B",
    x"2B1513B8",
    x"2B150116",
    x"2B14EE77",
    x"2B14DBDB",
    x"2B14C941",
    x"2B14B6A9",
    x"2B14A413",
    x"2B149180",
    x"2B147EEE",
    x"2B146C60",
    x"2B1459D3",
    x"2B144749",
    x"2B1434C2",
    x"2B14223C",
    x"2B140FB9",
    x"2B13FD38",
    x"2B13EABA",
    x"2B13D83E",
    x"2B13C5C4",
    x"2B13B34C",
    x"2B13A0D7",
    x"2B138E64",
    x"2B137BF3",
    x"2B136985",
    x"2B135719",
    x"2B1344AF",
    x"2B133248",
    x"2B131FE3",
    x"2B130D80",
    x"2B12FB1F",
    x"2B12E8C1",
    x"2B12D665",
    x"2B12C40B",
    x"2B12B1B4",
    x"2B129F5F",
    x"2B128D0C",
    x"2B127ABC",
    x"2B12686D",
    x"2B125622",
    x"2B1243D8",
    x"2B123191",
    x"2B121F4C",
    x"2B120D09",
    x"2B11FAC8",
    x"2B11E88A",
    x"2B11D64E",
    x"2B11C414",
    x"2B11B1DD",
    x"2B119FA8",
    x"2B118D75",
    x"2B117B45",
    x"2B116916",
    x"2B1156EA",
    x"2B1144C1",
    x"2B113299",
    x"2B112074",
    x"2B110E51",
    x"2B10FC30",
    x"2B10EA12",
    x"2B10D7F6",
    x"2B10C5DC",
    x"2B10B3C4",
    x"2B10A1AF",
    x"2B108F9C",
    x"2B107D8B",
    x"2B106B7D",
    x"2B105970",
    x"2B104766",
    x"2B10355E",
    x"2B102359",
    x"2B101156",
    x"2B0FFF55",
    x"2B0FED56",
    x"2B0FDB59",
    x"2B0FC95F",
    x"2B0FB767",
    x"2B0FA571",
    x"2B0F937E",
    x"2B0F818C",
    x"2B0F6F9D",
    x"2B0F5DB0",
    x"2B0F4BC6",
    x"2B0F39DD",
    x"2B0F27F7",
    x"2B0F1613",
    x"2B0F0432",
    x"2B0EF252",
    x"2B0EE075",
    x"2B0ECE9A",
    x"2B0EBCC2",
    x"2B0EAAEB",
    x"2B0E9917",
    x"2B0E8745",
    x"2B0E7575",
    x"2B0E63A7",
    x"2B0E51DC",
    x"2B0E4013",
    x"2B0E2E4C",
    x"2B0E1C87",
    x"2B0E0AC5",
    x"2B0DF905",
    x"2B0DE747",
    x"2B0DD58B",
    x"2B0DC3D1",
    x"2B0DB21A",
    x"2B0DA065",
    x"2B0D8EB2",
    x"2B0D7D01",
    x"2B0D6B53",
    x"2B0D59A6",
    x"2B0D47FC",
    x"2B0D3654",
    x"2B0D24AF",
    x"2B0D130B",
    x"2B0D016A",
    x"2B0CEFCB",
    x"2B0CDE2E",
    x"2B0CCC93",
    x"2B0CBAFB",
    x"2B0CA964",
    x"2B0C97D0",
    x"2B0C863E",
    x"2B0C74AF",
    x"2B0C6321",
    x"2B0C5196",
    x"2B0C400D",
    x"2B0C2E86",
    x"2B0C1D01",
    x"2B0C0B7F",
    x"2B0BF9FE",
    x"2B0BE880",
    x"2B0BD704",
    x"2B0BC58A",
    x"2B0BB413",
    x"2B0BA29D",
    x"2B0B912A",
    x"2B0B7FB9",
    x"2B0B6E4A",
    x"2B0B5CDE",
    x"2B0B4B73",
    x"2B0B3A0B",
    x"2B0B28A5",
    x"2B0B1741",
    x"2B0B05DF",
    x"2B0AF47F",
    x"2B0AE322",
    x"2B0AD1C6",
    x"2B0AC06D",
    x"2B0AAF16",
    x"2B0A9DC1",
    x"2B0A8C6F",
    x"2B0A7B1E",
    x"2B0A69D0",
    x"2B0A5884",
    x"2B0A473A",
    x"2B0A35F2",
    x"2B0A24AC",
    x"2B0A1369",
    x"2B0A0228",
    x"2B09F0E8",
    x"2B09DFAB",
    x"2B09CE70",
    x"2B09BD38",
    x"2B09AC01",
    x"2B099ACD",
    x"2B09899A",
    x"2B09786A",
    x"2B09673C",
    x"2B095610",
    x"2B0944E7",
    x"2B0933BF",
    x"2B09229A",
    x"2B091177",
    x"2B090055",
    x"2B08EF37",
    x"2B08DE1A",
    x"2B08CCFF",
    x"2B08BBE6",
    x"2B08AAD0",
    x"2B0899BC",
    x"2B0888AA",
    x"2B08779A",
    x"2B08668C",
    x"2B085580",
    x"2B084476",
    x"2B08336F",
    x"2B082269",
    x"2B081166",
    x"2B080065",
    x"2B07EF66",
    x"2B07DE69",
    x"2B07CD6F",
    x"2B07BC76",
    x"2B07AB7F",
    x"2B079A8B",
    x"2B078999",
    x"2B0778A9",
    x"2B0767BB",
    x"2B0756CF",
    x"2B0745E5",
    x"2B0734FD",
    x"2B072418",
    x"2B071334",
    x"2B070253",
    x"2B06F174",
    x"2B06E096",
    x"2B06CFBB",
    x"2B06BEE3",
    x"2B06AE0C",
    x"2B069D37",
    x"2B068C64",
    x"2B067B94",
    x"2B066AC6",
    x"2B0659F9",
    x"2B06492F",
    x"2B063867",
    x"2B0627A1",
    x"2B0616DD",
    x"2B06061B",
    x"2B05F55C",
    x"2B05E49E",
    x"2B05D3E2",
    x"2B05C329",
    x"2B05B272",
    x"2B05A1BC",
    x"2B059109",
    x"2B058058",
    x"2B056FA9",
    x"2B055EFC",
    x"2B054E51",
    x"2B053DA9",
    x"2B052D02",
    x"2B051C5D",
    x"2B050BBB",
    x"2B04FB1A",
    x"2B04EA7C",
    x"2B04D9E0",
    x"2B04C946",
    x"2B04B8AD",
    x"2B04A817",
    x"2B049783",
    x"2B0486F2",
    x"2B047662",
    x"2B0465D4",
    x"2B045548",
    x"2B0444BF",
    x"2B043437",
    x"2B0423B2",
    x"2B04132E",
    x"2B0402AD",
    x"2B03F22D",
    x"2B03E1B0",
    x"2B03D135",
    x"2B03C0BC",
    x"2B03B045",
    x"2B039FD0",
    x"2B038F5D",
    x"2B037EEC",
    x"2B036E7D",
    x"2B035E10",
    x"2B034DA6",
    x"2B033D3D",
    x"2B032CD6",
    x"2B031C72",
    x"2B030C0F",
    x"2B02FBAF",
    x"2B02EB50",
    x"2B02DAF4",
    x"2B02CA9A",
    x"2B02BA41",
    x"2B02A9EB",
    x"2B029997",
    x"2B028945",
    x"2B0278F4",
    x"2B0268A6",
    x"2B02585A",
    x"2B024810",
    x"2B0237C8",
    x"2B022782",
    x"2B02173E",
    x"2B0206FD",
    x"2B01F6BD",
    x"2B01E67F",
    x"2B01D643",
    x"2B01C609",
    x"2B01B5D2",
    x"2B01A59C",
    x"2B019568",
    x"2B018536",
    x"2B017507",
    x"2B0164D9",
    x"2B0154AE",
    x"2B014484",
    x"2B01345C",
    x"2B012437",
    x"2B011413",
    x"2B0103F2",
    x"2B00F3D2",
    x"2B00E3B5",
    x"2B00D399",
    x"2B00C380",
    x"2B00B369",
    x"2B00A353",
    x"2B009340",
    x"2B00832E",
    x"2B00731F",
    x"2B006312",
    x"2B005306",
    x"2B0042FD",
    x"2B0032F5",
    x"2B0022F0",
    x"2B0012ED",
    x"2B0002EB",
    x"2AFFE5D8",
    x"2AFFC5DD",
    x"2AFFA5E7",
    x"2AFF85F4",
    x"2AFF6605",
    x"2AFF461A",
    x"2AFF2634",
    x"2AFF0651",
    x"2AFEE672",
    x"2AFEC697",
    x"2AFEA6C0",
    x"2AFE86ED",
    x"2AFE671F",
    x"2AFE4754",
    x"2AFE278D",
    x"2AFE07CA",
    x"2AFDE80B",
    x"2AFDC850",
    x"2AFDA899",
    x"2AFD88E6",
    x"2AFD6937",
    x"2AFD498B",
    x"2AFD29E4",
    x"2AFD0A41",
    x"2AFCEAA2",
    x"2AFCCB06",
    x"2AFCAB6F",
    x"2AFC8BDB",
    x"2AFC6C4C",
    x"2AFC4CC0",
    x"2AFC2D39",
    x"2AFC0DB5",
    x"2AFBEE35",
    x"2AFBCEB9",
    x"2AFBAF42",
    x"2AFB8FCE",
    x"2AFB705E",
    x"2AFB50F1",
    x"2AFB3189",
    x"2AFB1225",
    x"2AFAF2C5",
    x"2AFAD368",
    x"2AFAB410",
    x"2AFA94BB",
    x"2AFA756B",
    x"2AFA561E",
    x"2AFA36D5",
    x"2AFA1790",
    x"2AF9F84F",
    x"2AF9D912",
    x"2AF9B9D9",
    x"2AF99AA4",
    x"2AF97B72",
    x"2AF95C45",
    x"2AF93D1B",
    x"2AF91DF6",
    x"2AF8FED4",
    x"2AF8DFB6",
    x"2AF8C09C",
    x"2AF8A186",
    x"2AF88274",
    x"2AF86365",
    x"2AF8445B",
    x"2AF82554",
    x"2AF80651",
    x"2AF7E753",
    x"2AF7C858",
    x"2AF7A960",
    x"2AF78A6D",
    x"2AF76B7E",
    x"2AF74C92",
    x"2AF72DAB",
    x"2AF70EC7",
    x"2AF6EFE7",
    x"2AF6D10B",
    x"2AF6B233",
    x"2AF6935E",
    x"2AF6748E",
    x"2AF655C1",
    x"2AF636F8",
    x"2AF61833",
    x"2AF5F972",
    x"2AF5DAB5",
    x"2AF5BBFC",
    x"2AF59D46",
    x"2AF57E94",
    x"2AF55FE6",
    x"2AF5413C",
    x"2AF52296",
    x"2AF503F4",
    x"2AF4E555",
    x"2AF4C6BA",
    x"2AF4A824",
    x"2AF48990",
    x"2AF46B01",
    x"2AF44C76",
    x"2AF42DEE",
    x"2AF40F6A",
    x"2AF3F0EA",
    x"2AF3D26E",
    x"2AF3B3F6",
    x"2AF39581",
    x"2AF37710",
    x"2AF358A3",
    x"2AF33A3A",
    x"2AF31BD5",
    x"2AF2FD73",
    x"2AF2DF15",
    x"2AF2C0BB",
    x"2AF2A265",
    x"2AF28413",
    x"2AF265C4",
    x"2AF24779",
    x"2AF22932",
    x"2AF20AEF",
    x"2AF1ECAF",
    x"2AF1CE74",
    x"2AF1B03C",
    x"2AF19208",
    x"2AF173D7",
    x"2AF155AB",
    x"2AF13782",
    x"2AF1195D",
    x"2AF0FB3C",
    x"2AF0DD1E",
    x"2AF0BF04",
    x"2AF0A0EE",
    x"2AF082DC",
    x"2AF064CE",
    x"2AF046C3",
    x"2AF028BC",
    x"2AF00AB9",
    x"2AEFECB9",
    x"2AEFCEBD",
    x"2AEFB0C6",
    x"2AEF92D1",
    x"2AEF74E1",
    x"2AEF56F4",
    x"2AEF390B",
    x"2AEF1B26",
    x"2AEEFD44",
    x"2AEEDF67",
    x"2AEEC18C",
    x"2AEEA3B6",
    x"2AEE85E4",
    x"2AEE6815",
    x"2AEE4A49",
    x"2AEE2C82",
    x"2AEE0EBE",
    x"2AEDF0FE",
    x"2AEDD342",
    x"2AEDB58A",
    x"2AED97D5",
    x"2AED7A24",
    x"2AED5C76",
    x"2AED3ECC",
    x"2AED2126",
    x"2AED0384",
    x"2AECE5E6",
    x"2AECC84B",
    x"2AECAAB4",
    x"2AEC8D20",
    x"2AEC6F90",
    x"2AEC5204",
    x"2AEC347C",
    x"2AEC16F7",
    x"2AEBF976",
    x"2AEBDBF9",
    x"2AEBBE7F",
    x"2AEBA109",
    x"2AEB8397",
    x"2AEB6628",
    x"2AEB48BD",
    x"2AEB2B56",
    x"2AEB0DF2",
    x"2AEAF092",
    x"2AEAD336",
    x"2AEAB5DE",
    x"2AEA9889",
    x"2AEA7B38",
    x"2AEA5DEA",
    x"2AEA40A0",
    x"2AEA235A",
    x"2AEA0617",
    x"2AE9E8D8",
    x"2AE9CB9D",
    x"2AE9AE65",
    x"2AE99131",
    x"2AE97401",
    x"2AE956D4",
    x"2AE939AB",
    x"2AE91C86",
    x"2AE8FF64",
    x"2AE8E246",
    x"2AE8C52C",
    x"2AE8A815",
    x"2AE88B02",
    x"2AE86DF2",
    x"2AE850E6",
    x"2AE833DE",
    x"2AE816D9",
    x"2AE7F9D8",
    x"2AE7DCDB",
    x"2AE7BFE1",
    x"2AE7A2EB",
    x"2AE785F8",
    x"2AE76909",
    x"2AE74C1E",
    x"2AE72F36",
    x"2AE71252",
    x"2AE6F572",
    x"2AE6D895",
    x"2AE6BBBC",
    x"2AE69EE6",
    x"2AE68214",
    x"2AE66545",
    x"2AE6487A",
    x"2AE62BB3",
    x"2AE60EF0",
    x"2AE5F22F",
    x"2AE5D573",
    x"2AE5B8BA",
    x"2AE59C05",
    x"2AE57F53",
    x"2AE562A5",
    x"2AE545FA",
    x"2AE52953",
    x"2AE50CB0",
    x"2AE4F010",
    x"2AE4D374",
    x"2AE4B6DB",
    x"2AE49A46",
    x"2AE47DB5",
    x"2AE46127",
    x"2AE4449D",
    x"2AE42816",
    x"2AE40B93",
    x"2AE3EF13",
    x"2AE3D297",
    x"2AE3B61E",
    x"2AE399A9",
    x"2AE37D38",
    x"2AE360CA",
    x"2AE34460",
    x"2AE327F9",
    x"2AE30B96",
    x"2AE2EF36",
    x"2AE2D2DA",
    x"2AE2B681",
    x"2AE29A2C",
    x"2AE27DDB",
    x"2AE2618D",
    x"2AE24542",
    x"2AE228FB",
    x"2AE20CB8",
    x"2AE1F078",
    x"2AE1D43C",
    x"2AE1B803",
    x"2AE19BCE",
    x"2AE17F9C",
    x"2AE1636E",
    x"2AE14743",
    x"2AE12B1C",
    x"2AE10EF9",
    x"2AE0F2D9",
    x"2AE0D6BC",
    x"2AE0BAA3",
    x"2AE09E8D",
    x"2AE0827B",
    x"2AE0666D",
    x"2AE04A62",
    x"2AE02E5A",
    x"2AE01256",
    x"2ADFF655",
    x"2ADFDA58",
    x"2ADFBE5F",
    x"2ADFA269",
    x"2ADF8676",
    x"2ADF6A87",
    x"2ADF4E9C",
    x"2ADF32B4",
    x"2ADF16CF",
    x"2ADEFAEE",
    x"2ADEDF10",
    x"2ADEC336",
    x"2ADEA75F",
    x"2ADE8B8C",
    x"2ADE6FBD",
    x"2ADE53F0",
    x"2ADE3828",
    x"2ADE1C62",
    x"2ADE00A0",
    x"2ADDE4E2",
    x"2ADDC927",
    x"2ADDAD70",
    x"2ADD91BC",
    x"2ADD760B",
    x"2ADD5A5E",
    x"2ADD3EB5",
    x"2ADD230F",
    x"2ADD076C",
    x"2ADCEBCD",
    x"2ADCD031",
    x"2ADCB499",
    x"2ADC9904",
    x"2ADC7D73",
    x"2ADC61E5",
    x"2ADC465A",
    x"2ADC2AD3",
    x"2ADC0F4F",
    x"2ADBF3CF",
    x"2ADBD852",
    x"2ADBBCD9",
    x"2ADBA163",
    x"2ADB85F1",
    x"2ADB6A82",
    x"2ADB4F16",
    x"2ADB33AE",
    x"2ADB1849",
    x"2ADAFCE8",
    x"2ADAE18A",
    x"2ADAC62F",
    x"2ADAAAD8",
    x"2ADA8F85",
    x"2ADA7435",
    x"2ADA58E8",
    x"2ADA3D9E",
    x"2ADA2258",
    x"2ADA0716",
    x"2AD9EBD7",
    x"2AD9D09B",
    x"2AD9B562",
    x"2AD99A2D",
    x"2AD97EFC",
    x"2AD963CE",
    x"2AD948A3",
    x"2AD92D7B",
    x"2AD91257",
    x"2AD8F737",
    x"2AD8DC1A",
    x"2AD8C100",
    x"2AD8A5E9",
    x"2AD88AD6",
    x"2AD86FC7",
    x"2AD854BA",
    x"2AD839B2",
    x"2AD81EAC",
    x"2AD803AA",
    x"2AD7E8AB",
    x"2AD7CDB0",
    x"2AD7B2B8",
    x"2AD797C3",
    x"2AD77CD2",
    x"2AD761E4",
    x"2AD746F9",
    x"2AD72C12",
    x"2AD7112E",
    x"2AD6F64E",
    x"2AD6DB71",
    x"2AD6C097",
    x"2AD6A5C1",
    x"2AD68AED",
    x"2AD6701E",
    x"2AD65551",
    x"2AD63A88",
    x"2AD61FC3",
    x"2AD60501",
    x"2AD5EA42",
    x"2AD5CF86",
    x"2AD5B4CE",
    x"2AD59A19",
    x"2AD57F67",
    x"2AD564B9",
    x"2AD54A0E",
    x"2AD52F66",
    x"2AD514C2",
    x"2AD4FA21",
    x"2AD4DF84",
    x"2AD4C4E9",
    x"2AD4AA52",
    x"2AD48FBF",
    x"2AD4752E",
    x"2AD45AA1",
    x"2AD44018",
    x"2AD42591",
    x"2AD40B0E",
    x"2AD3F08F",
    x"2AD3D612",
    x"2AD3BB99",
    x"2AD3A123",
    x"2AD386B1",
    x"2AD36C42",
    x"2AD351D6",
    x"2AD3376D",
    x"2AD31D08",
    x"2AD302A6",
    x"2AD2E847",
    x"2AD2CDEC",
    x"2AD2B394",
    x"2AD2993F",
    x"2AD27EED",
    x"2AD2649F",
    x"2AD24A54",
    x"2AD2300D",
    x"2AD215C8",
    x"2AD1FB87",
    x"2AD1E149",
    x"2AD1C70F",
    x"2AD1ACD8",
    x"2AD192A4",
    x"2AD17873",
    x"2AD15E46",
    x"2AD1441B",
    x"2AD129F5",
    x"2AD10FD1",
    x"2AD0F5B1",
    x"2AD0DB94",
    x"2AD0C17A",
    x"2AD0A763",
    x"2AD08D50",
    x"2AD07340",
    x"2AD05933",
    x"2AD03F2A",
    x"2AD02523",
    x"2AD00B20",
    x"2ACFF120",
    x"2ACFD724",
    x"2ACFBD2B",
    x"2ACFA335",
    x"2ACF8942",
    x"2ACF6F52",
    x"2ACF5566",
    x"2ACF3B7D",
    x"2ACF2197",
    x"2ACF07B5",
    x"2ACEEDD5",
    x"2ACED3F9",
    x"2ACEBA20",
    x"2ACEA04B",
    x"2ACE8678",
    x"2ACE6CA9",
    x"2ACE52DD",
    x"2ACE3914",
    x"2ACE1F4F",
    x"2ACE058C",
    x"2ACDEBCD",
    x"2ACDD212",
    x"2ACDB859",
    x"2ACD9EA3",
    x"2ACD84F1",
    x"2ACD6B42",
    x"2ACD5196",
    x"2ACD37EE",
    x"2ACD1E48",
    x"2ACD04A6",
    x"2ACCEB07",
    x"2ACCD16B",
    x"2ACCB7D3",
    x"2ACC9E3D",
    x"2ACC84AB",
    x"2ACC6B1C",
    x"2ACC5191",
    x"2ACC3808",
    x"2ACC1E83",
    x"2ACC0500",
    x"2ACBEB81",
    x"2ACBD205",
    x"2ACBB88D",
    x"2ACB9F17",
    x"2ACB85A5",
    x"2ACB6C36",
    x"2ACB52CA",
    x"2ACB3961",
    x"2ACB1FFC",
    x"2ACB0699",
    x"2ACAED3A",
    x"2ACAD3DE",
    x"2ACABA85",
    x"2ACAA12F",
    x"2ACA87DD",
    x"2ACA6E8D",
    x"2ACA5541",
    x"2ACA3BF8",
    x"2ACA22B2",
    x"2ACA096F",
    x"2AC9F030",
    x"2AC9D6F3",
    x"2AC9BDBA",
    x"2AC9A484",
    x"2AC98B51",
    x"2AC97221",
    x"2AC958F4",
    x"2AC93FCB",
    x"2AC926A4",
    x"2AC90D81",
    x"2AC8F461",
    x"2AC8DB44",
    x"2AC8C22A",
    x"2AC8A913",
    x"2AC89000",
    x"2AC876EF",
    x"2AC85DE2",
    x"2AC844D8",
    x"2AC82BD1",
    x"2AC812CD",
    x"2AC7F9CC",
    x"2AC7E0CF",
    x"2AC7C7D4",
    x"2AC7AEDD",
    x"2AC795E8",
    x"2AC77CF7",
    x"2AC76409",
    x"2AC74B1E",
    x"2AC73236",
    x"2AC71952",
    x"2AC70070",
    x"2AC6E791",
    x"2AC6CEB6",
    x"2AC6B5DE",
    x"2AC69D09",
    x"2AC68437",
    x"2AC66B68",
    x"2AC6529C",
    x"2AC639D3",
    x"2AC6210D",
    x"2AC6084B",
    x"2AC5EF8B",
    x"2AC5D6CF",
    x"2AC5BE15",
    x"2AC5A55F",
    x"2AC58CAC",
    x"2AC573FC",
    x"2AC55B4F",
    x"2AC542A5",
    x"2AC529FE",
    x"2AC5115B",
    x"2AC4F8BA",
    x"2AC4E01D",
    x"2AC4C782",
    x"2AC4AEEB",
    x"2AC49656",
    x"2AC47DC5",
    x"2AC46537",
    x"2AC44CAC",
    x"2AC43424",
    x"2AC41B9F",
    x"2AC4031D",
    x"2AC3EA9E",
    x"2AC3D222",
    x"2AC3B9A9",
    x"2AC3A134",
    x"2AC388C1",
    x"2AC37052",
    x"2AC357E5",
    x"2AC33F7C",
    x"2AC32715",
    x"2AC30EB2",
    x"2AC2F652",
    x"2AC2DDF4",
    x"2AC2C59A",
    x"2AC2AD43",
    x"2AC294EF",
    x"2AC27C9E",
    x"2AC26450",
    x"2AC24C05",
    x"2AC233BD",
    x"2AC21B78",
    x"2AC20336",
    x"2AC1EAF7",
    x"2AC1D2BB",
    x"2AC1BA82",
    x"2AC1A24C",
    x"2AC18A1A",
    x"2AC171EA",
    x"2AC159BD",
    x"2AC14193",
    x"2AC1296D",
    x"2AC11149",
    x"2AC0F928",
    x"2AC0E10B",
    x"2AC0C8F0",
    x"2AC0B0D8",
    x"2AC098C4",
    x"2AC080B2",
    x"2AC068A4",
    x"2AC05098",
    x"2AC03890",
    x"2AC0208A",
    x"2AC00887",
    x"2ABFF088",
    x"2ABFD88B",
    x"2ABFC092",
    x"2ABFA89B",
    x"2ABF90A8",
    x"2ABF78B7",
    x"2ABF60C9",
    x"2ABF48DF",
    x"2ABF30F7",
    x"2ABF1913",
    x"2ABF0131",
    x"2ABEE952",
    x"2ABED177",
    x"2ABEB99E",
    x"2ABEA1C8",
    x"2ABE89F5",
    x"2ABE7226",
    x"2ABE5A59",
    x"2ABE428F",
    x"2ABE2AC8",
    x"2ABE1304",
    x"2ABDFB43",
    x"2ABDE386",
    x"2ABDCBCB",
    x"2ABDB413",
    x"2ABD9C5E",
    x"2ABD84AC",
    x"2ABD6CFC",
    x"2ABD5550",
    x"2ABD3DA7",
    x"2ABD2601",
    x"2ABD0E5E",
    x"2ABCF6BD",
    x"2ABCDF20",
    x"2ABCC785",
    x"2ABCAFEE",
    x"2ABC985A",
    x"2ABC80C8",
    x"2ABC6939",
    x"2ABC51AE",
    x"2ABC3A25",
    x"2ABC229F",
    x"2ABC0B1C",
    x"2ABBF39C",
    x"2ABBDC1F",
    x"2ABBC4A5",
    x"2ABBAD2E",
    x"2ABB95BA",
    x"2ABB7E49",
    x"2ABB66DA",
    x"2ABB4F6F",
    x"2ABB3807",
    x"2ABB20A1",
    x"2ABB093E",
    x"2ABAF1DF",
    x"2ABADA82",
    x"2ABAC328",
    x"2ABAABD1",
    x"2ABA947D",
    x"2ABA7D2C",
    x"2ABA65DE",
    x"2ABA4E93",
    x"2ABA374A",
    x"2ABA2005",
    x"2ABA08C2",
    x"2AB9F183",
    x"2AB9DA46",
    x"2AB9C30C",
    x"2AB9ABD5",
    x"2AB994A1",
    x"2AB97D70",
    x"2AB96642",
    x"2AB94F16",
    x"2AB937EE",
    x"2AB920C8",
    x"2AB909A6",
    x"2AB8F286",
    x"2AB8DB69",
    x"2AB8C44F",
    x"2AB8AD38",
    x"2AB89624",
    x"2AB87F12",
    x"2AB86804",
    x"2AB850F8",
    x"2AB839F0",
    x"2AB822EA",
    x"2AB80BE7",
    x"2AB7F4E7",
    x"2AB7DDEA",
    x"2AB7C6EF",
    x"2AB7AFF8",
    x"2AB79904",
    x"2AB78212",
    x"2AB76B23",
    x"2AB75437",
    x"2AB73D4E",
    x"2AB72668",
    x"2AB70F84",
    x"2AB6F8A4",
    x"2AB6E1C6",
    x"2AB6CAEB",
    x"2AB6B413",
    x"2AB69D3E",
    x"2AB6866C",
    x"2AB66F9D",
    x"2AB658D0",
    x"2AB64207",
    x"2AB62B40",
    x"2AB6147C",
    x"2AB5FDBB",
    x"2AB5E6FC",
    x"2AB5D041",
    x"2AB5B988",
    x"2AB5A2D2",
    x"2AB58C20",
    x"2AB5756F",
    x"2AB55EC2",
    x"2AB54818",
    x"2AB53170",
    x"2AB51ACB",
    x"2AB50429",
    x"2AB4ED8A",
    x"2AB4D6EE",
    x"2AB4C055",
    x"2AB4A9BE",
    x"2AB4932A",
    x"2AB47C99",
    x"2AB4660B",
    x"2AB44F80",
    x"2AB438F7",
    x"2AB42271",
    x"2AB40BEF",
    x"2AB3F56E",
    x"2AB3DEF1",
    x"2AB3C877",
    x"2AB3B1FF",
    x"2AB39B8A",
    x"2AB38518",
    x"2AB36EA9",
    x"2AB3583D",
    x"2AB341D3",
    x"2AB32B6C",
    x"2AB31508",
    x"2AB2FEA7",
    x"2AB2E848",
    x"2AB2D1ED",
    x"2AB2BB94",
    x"2AB2A53E",
    x"2AB28EEB",
    x"2AB2789A",
    x"2AB2624C",
    x"2AB24C02",
    x"2AB235B9",
    x"2AB21F74",
    x"2AB20932",
    x"2AB1F2F2",
    x"2AB1DCB5",
    x"2AB1C67B",
    x"2AB1B043",
    x"2AB19A0F",
    x"2AB183DD",
    x"2AB16DAE",
    x"2AB15781",
    x"2AB14158",
    x"2AB12B31",
    x"2AB1150D",
    x"2AB0FEEC",
    x"2AB0E8CD",
    x"2AB0D2B1",
    x"2AB0BC99",
    x"2AB0A682",
    x"2AB0906F",
    x"2AB07A5E",
    x"2AB06450",
    x"2AB04E45",
    x"2AB0383D",
    x"2AB02237",
    x"2AB00C34",
    x"2AAFF634",
    x"2AAFE037",
    x"2AAFCA3C",
    x"2AAFB444",
    x"2AAF9E4F",
    x"2AAF885C",
    x"2AAF726D",
    x"2AAF5C80",
    x"2AAF4696",
    x"2AAF30AE",
    x"2AAF1ACA",
    x"2AAF04E8",
    x"2AAEEF08",
    x"2AAED92C",
    x"2AAEC352",
    x"2AAEAD7B",
    x"2AAE97A7",
    x"2AAE81D5",
    x"2AAE6C06",
    x"2AAE563A",
    x"2AAE4071",
    x"2AAE2AAA",
    x"2AAE14E6",
    x"2AADFF25",
    x"2AADE966",
    x"2AADD3AA",
    x"2AADBDF1",
    x"2AADA83B",
    x"2AAD9287",
    x"2AAD7CD6",
    x"2AAD6728",
    x"2AAD517C",
    x"2AAD3BD4",
    x"2AAD262D",
    x"2AAD108A",
    x"2AACFAE9",
    x"2AACE54B",
    x"2AACCFB0",
    x"2AACBA17",
    x"2AACA481",
    x"2AAC8EEE",
    x"2AAC795E",
    x"2AAC63D0",
    x"2AAC4E45",
    x"2AAC38BC",
    x"2AAC2337",
    x"2AAC0DB4",
    x"2AABF833",
    x"2AABE2B6",
    x"2AABCD3B",
    x"2AABB7C2",
    x"2AABA24D",
    x"2AAB8CDA",
    x"2AAB7769",
    x"2AAB61FC",
    x"2AAB4C91",
    x"2AAB3729",
    x"2AAB21C3",
    x"2AAB0C60",
    x"2AAAF700",
    x"2AAAE1A2",
    x"2AAACC48",
    x"2AAAB6EF",
    x"2AAAA19A",
    x"2AAA8C47",
    x"2AAA76F7",
    x"2AAA61A9",
    x"2AAA4C5E",
    x"2AAA3716",
    x"2AAA21D1",
    x"2AAA0C8E",
    x"2AA9F74D",
    x"2AA9E210",
    x"2AA9CCD5",
    x"2AA9B79D",
    x"2AA9A267",
    x"2AA98D34",
    x"2AA97804",
    x"2AA962D6",
    x"2AA94DAB",
    x"2AA93883",
    x"2AA9235D",
    x"2AA90E3A",
    x"2AA8F919",
    x"2AA8E3FC",
    x"2AA8CEE0",
    x"2AA8B9C8",
    x"2AA8A4B2",
    x"2AA88F9F",
    x"2AA87A8E",
    x"2AA86580",
    x"2AA85075",
    x"2AA83B6C",
    x"2AA82666",
    x"2AA81162",
    x"2AA7FC61",
    x"2AA7E763",
    x"2AA7D268",
    x"2AA7BD6F",
    x"2AA7A878",
    x"2AA79384",
    x"2AA77E93",
    x"2AA769A5",
    x"2AA754B9",
    x"2AA73FD0",
    x"2AA72AE9",
    x"2AA71605",
    x"2AA70123",
    x"2AA6EC45",
    x"2AA6D768",
    x"2AA6C28F",
    x"2AA6ADB8",
    x"2AA698E3",
    x"2AA68412",
    x"2AA66F42",
    x"2AA65A76",
    x"2AA645AC",
    x"2AA630E4",
    x"2AA61C1F",
    x"2AA6075D",
    x"2AA5F29E",
    x"2AA5DDE1",
    x"2AA5C926",
    x"2AA5B46E",
    x"2AA59FB9",
    x"2AA58B06",
    x"2AA57656",
    x"2AA561A9",
    x"2AA54CFE",
    x"2AA53856",
    x"2AA523B0",
    x"2AA50F0D",
    x"2AA4FA6C",
    x"2AA4E5CE",
    x"2AA4D133",
    x"2AA4BC9A",
    x"2AA4A803",
    x"2AA49370",
    x"2AA47EDF",
    x"2AA46A50",
    x"2AA455C4",
    x"2AA4413B",
    x"2AA42CB4",
    x"2AA4182F",
    x"2AA403AE",
    x"2AA3EF2E",
    x"2AA3DAB2",
    x"2AA3C638",
    x"2AA3B1C0",
    x"2AA39D4B",
    x"2AA388D9",
    x"2AA37469",
    x"2AA35FFC",
    x"2AA34B91",
    x"2AA33729",
    x"2AA322C3",
    x"2AA30E60",
    x"2AA2FA00",
    x"2AA2E5A2",
    x"2AA2D146",
    x"2AA2BCED",
    x"2AA2A897",
    x"2AA29443",
    x"2AA27FF2",
    x"2AA26BA3",
    x"2AA25757",
    x"2AA2430D",
    x"2AA22EC6",
    x"2AA21A82",
    x"2AA20640",
    x"2AA1F200",
    x"2AA1DDC3",
    x"2AA1C989",
    x"2AA1B551",
    x"2AA1A11B",
    x"2AA18CE9",
    x"2AA178B8",
    x"2AA1648A",
    x"2AA1505F",
    x"2AA13C36",
    x"2AA12810",
    x"2AA113EC",
    x"2AA0FFCB",
    x"2AA0EBAC",
    x"2AA0D790",
    x"2AA0C376",
    x"2AA0AF5F",
    x"2AA09B4B",
    x"2AA08738",
    x"2AA07329",
    x"2AA05F1C",
    x"2AA04B11",
    x"2AA03709",
    x"2AA02303",
    x"2AA00F00",
    x"2A9FFB00",
    x"2A9FE701",
    x"2A9FD306",
    x"2A9FBF0D",
    x"2A9FAB16",
    x"2A9F9722",
    x"2A9F8330",
    x"2A9F6F41",
    x"2A9F5B54",
    x"2A9F476A",
    x"2A9F3383",
    x"2A9F1F9D",
    x"2A9F0BBB",
    x"2A9EF7DA",
    x"2A9EE3FD",
    x"2A9ED021",
    x"2A9EBC49",
    x"2A9EA872",
    x"2A9E949F",
    x"2A9E80CD",
    x"2A9E6CFE",
    x"2A9E5932",
    x"2A9E4568",
    x"2A9E31A1",
    x"2A9E1DDC",
    x"2A9E0A19",
    x"2A9DF659",
    x"2A9DE29C",
    x"2A9DCEE0",
    x"2A9DBB28",
    x"2A9DA772",
    x"2A9D93BE",
    x"2A9D800D",
    x"2A9D6C5E",
    x"2A9D58B2",
    x"2A9D4508",
    x"2A9D3160",
    x"2A9D1DBB",
    x"2A9D0A19",
    x"2A9CF679",
    x"2A9CE2DB",
    x"2A9CCF40",
    x"2A9CBBA8",
    x"2A9CA811",
    x"2A9C947D",
    x"2A9C80EC",
    x"2A9C6D5D",
    x"2A9C59D1",
    x"2A9C4647",
    x"2A9C32BF",
    x"2A9C1F3A",
    x"2A9C0BB7",
    x"2A9BF837",
    x"2A9BE4B9",
    x"2A9BD13E",
    x"2A9BBDC5",
    x"2A9BAA4F",
    x"2A9B96DA",
    x"2A9B8369",
    x"2A9B6FFA",
    x"2A9B5C8D",
    x"2A9B4923",
    x"2A9B35BB",
    x"2A9B2255",
    x"2A9B0EF2",
    x"2A9AFB91",
    x"2A9AE833",
    x"2A9AD4D7",
    x"2A9AC17E",
    x"2A9AAE27",
    x"2A9A9AD2",
    x"2A9A8780",
    x"2A9A7430",
    x"2A9A60E3",
    x"2A9A4D98",
    x"2A9A3A50",
    x"2A9A270A",
    x"2A9A13C6",
    x"2A9A0085",
    x"2A99ED46",
    x"2A99DA09",
    x"2A99C6CF",
    x"2A99B398",
    x"2A99A062",
    x"2A998D30",
    x"2A9979FF",
    x"2A9966D1",
    x"2A9953A5",
    x"2A99407C",
    x"2A992D55",
    x"2A991A31",
    x"2A99070F",
    x"2A98F3EF",
    x"2A98E0D2",
    x"2A98CDB7",
    x"2A98BA9E",
    x"2A98A788",
    x"2A989474",
    x"2A988163",
    x"2A986E54",
    x"2A985B48",
    x"2A98483D",
    x"2A983535",
    x"2A982230",
    x"2A980F2D",
    x"2A97FC2C",
    x"2A97E92E",
    x"2A97D632",
    x"2A97C338",
    x"2A97B041",
    x"2A979D4C",
    x"2A978A5A",
    x"2A97776A",
    x"2A97647C",
    x"2A975191",
    x"2A973EA8",
    x"2A972BC1",
    x"2A9718DD",
    x"2A9705FB",
    x"2A96F31B",
    x"2A96E03E",
    x"2A96CD63",
    x"2A96BA8B",
    x"2A96A7B4",
    x"2A9694E1",
    x"2A96820F",
    x"2A966F40",
    x"2A965C73",
    x"2A9649A9",
    x"2A9636E1",
    x"2A96241B",
    x"2A961158",
    x"2A95FE97",
    x"2A95EBD8",
    x"2A95D91C",
    x"2A95C662",
    x"2A95B3AA",
    x"2A95A0F5",
    x"2A958E42",
    x"2A957B92",
    x"2A9568E3",
    x"2A955637",
    x"2A95438E",
    x"2A9530E6",
    x"2A951E41",
    x"2A950B9F",
    x"2A94F8FF",
    x"2A94E661",
    x"2A94D3C5",
    x"2A94C12C",
    x"2A94AE95",
    x"2A949C00",
    x"2A94896E",
    x"2A9476DE",
    x"2A946450",
    x"2A9451C5",
    x"2A943F3C",
    x"2A942CB5",
    x"2A941A30",
    x"2A9407AE",
    x"2A93F52E",
    x"2A93E2B1",
    x"2A93D036",
    x"2A93BDBD",
    x"2A93AB46",
    x"2A9398D2",
    x"2A938660",
    x"2A9373F0",
    x"2A936183",
    x"2A934F18",
    x"2A933CAF",
    x"2A932A49",
    x"2A9317E5",
    x"2A930583",
    x"2A92F323",
    x"2A92E0C6",
    x"2A92CE6B",
    x"2A92BC13",
    x"2A92A9BC",
    x"2A929768",
    x"2A928516",
    x"2A9272C7",
    x"2A92607A",
    x"2A924E2F",
    x"2A923BE6",
    x"2A9229A0",
    x"2A92175C",
    x"2A92051A",
    x"2A91F2DA",
    x"2A91E09D",
    x"2A91CE62",
    x"2A91BC2A",
    x"2A91A9F3",
    x"2A9197BF",
    x"2A91858D",
    x"2A91735E",
    x"2A916130",
    x"2A914F05",
    x"2A913CDD",
    x"2A912AB6",
    x"2A911892",
    x"2A910670",
    x"2A90F450",
    x"2A90E233",
    x"2A90D018",
    x"2A90BDFF",
    x"2A90ABE8",
    x"2A9099D4",
    x"2A9087C2",
    x"2A9075B2",
    x"2A9063A4",
    x"2A905199",
    x"2A903F90",
    x"2A902D89",
    x"2A901B85",
    x"2A900982",
    x"2A8FF782",
    x"2A8FE585",
    x"2A8FD389",
    x"2A8FC190",
    x"2A8FAF99",
    x"2A8F9DA4",
    x"2A8F8BB1",
    x"2A8F79C1",
    x"2A8F67D3",
    x"2A8F55E7",
    x"2A8F43FD",
    x"2A8F3216",
    x"2A8F2031",
    x"2A8F0E4E",
    x"2A8EFC6D",
    x"2A8EEA8F",
    x"2A8ED8B2",
    x"2A8EC6D9",
    x"2A8EB501",
    x"2A8EA32B",
    x"2A8E9158",
    x"2A8E7F87",
    x"2A8E6DB8",
    x"2A8E5BEB",
    x"2A8E4A21",
    x"2A8E3859",
    x"2A8E2693",
    x"2A8E14CF",
    x"2A8E030E",
    x"2A8DF14F",
    x"2A8DDF91",
    x"2A8DCDD7",
    x"2A8DBC1E",
    x"2A8DAA68",
    x"2A8D98B3",
    x"2A8D8701",
    x"2A8D7552",
    x"2A8D63A4",
    x"2A8D51F9",
    x"2A8D4050",
    x"2A8D2EA9",
    x"2A8D1D04",
    x"2A8D0B61",
    x"2A8CF9C1",
    x"2A8CE823",
    x"2A8CD687",
    x"2A8CC4ED",
    x"2A8CB356",
    x"2A8CA1C1",
    x"2A8C902D",
    x"2A8C7E9C",
    x"2A8C6D0E",
    x"2A8C5B81",
    x"2A8C49F7",
    x"2A8C386F",
    x"2A8C26E9",
    x"2A8C1565",
    x"2A8C03E3",
    x"2A8BF264",
    x"2A8BE0E7",
    x"2A8BCF6C",
    x"2A8BBDF3",
    x"2A8BAC7C",
    x"2A8B9B08",
    x"2A8B8996",
    x"2A8B7825",
    x"2A8B66B8",
    x"2A8B554C",
    x"2A8B43E2",
    x"2A8B327B",
    x"2A8B2116",
    x"2A8B0FB3",
    x"2A8AFE52",
    x"2A8AECF3",
    x"2A8ADB96",
    x"2A8ACA3C",
    x"2A8AB8E4",
    x"2A8AA78E",
    x"2A8A963A",
    x"2A8A84E8",
    x"2A8A7399",
    x"2A8A624B",
    x"2A8A5100",
    x"2A8A3FB7",
    x"2A8A2E70",
    x"2A8A1D2C",
    x"2A8A0BE9",
    x"2A89FAA9",
    x"2A89E96A",
    x"2A89D82E",
    x"2A89C6F4",
    x"2A89B5BC",
    x"2A89A487",
    x"2A899353",
    x"2A898222",
    x"2A8970F3",
    x"2A895FC6",
    x"2A894E9B",
    x"2A893D72",
    x"2A892C4B",
    x"2A891B27",
    x"2A890A05",
    x"2A88F8E5",
    x"2A88E7C6",
    x"2A88D6AB",
    x"2A88C591",
    x"2A88B479",
    x"2A88A364",
    x"2A889250",
    x"2A88813F",
    x"2A887030",
    x"2A885F23",
    x"2A884E18",
    x"2A883D10",
    x"2A882C09",
    x"2A881B05",
    x"2A880A02",
    x"2A87F902",
    x"2A87E804",
    x"2A87D708",
    x"2A87C60E",
    x"2A87B516",
    x"2A87A421",
    x"2A87932D",
    x"2A87823C",
    x"2A87714D",
    x"2A876060",
    x"2A874F75",
    x"2A873E8C",
    x"2A872DA5",
    x"2A871CC1",
    x"2A870BDE",
    x"2A86FAFE",
    x"2A86EA1F",
    x"2A86D943",
    x"2A86C869",
    x"2A86B791",
    x"2A86A6BB",
    x"2A8695E7",
    x"2A868516",
    x"2A867446",
    x"2A866378",
    x"2A8652AD",
    x"2A8641E4",
    x"2A86311D",
    x"2A862058",
    x"2A860F95",
    x"2A85FED4",
    x"2A85EE15",
    x"2A85DD58",
    x"2A85CC9E",
    x"2A85BBE5",
    x"2A85AB2F",
    x"2A859A7A",
    x"2A8589C8",
    x"2A857918",
    x"2A85686A",
    x"2A8557BE",
    x"2A854714",
    x"2A85366C",
    x"2A8525C6",
    x"2A851522",
    x"2A850481",
    x"2A84F3E1",
    x"2A84E344",
    x"2A84D2A8",
    x"2A84C20F",
    x"2A84B178",
    x"2A84A0E3",
    x"2A849050",
    x"2A847FBF",
    x"2A846F30",
    x"2A845EA3",
    x"2A844E18",
    x"2A843D8F",
    x"2A842D09",
    x"2A841C84",
    x"2A840C02",
    x"2A83FB81",
    x"2A83EB03",
    x"2A83DA86",
    x"2A83CA0C",
    x"2A83B994",
    x"2A83A91E",
    x"2A8398AA",
    x"2A838838",
    x"2A8377C8",
    x"2A83675A",
    x"2A8356EE",
    x"2A834684",
    x"2A83361C",
    x"2A8325B6",
    x"2A831553",
    x"2A8304F1",
    x"2A82F491",
    x"2A82E434",
    x"2A82D3D8",
    x"2A82C37F",
    x"2A82B327",
    x"2A82A2D2",
    x"2A82927F",
    x"2A82822D",
    x"2A8271DE",
    x"2A826191",
    x"2A825146",
    x"2A8240FD",
    x"2A8230B6",
    x"2A822071",
    x"2A82102D",
    x"2A81FFEC",
    x"2A81EFAE",
    x"2A81DF71",
    x"2A81CF36",
    x"2A81BEFD",
    x"2A81AEC6",
    x"2A819E91",
    x"2A818E5E",
    x"2A817E2D",
    x"2A816DFF",
    x"2A815DD2",
    x"2A814DA7",
    x"2A813D7F",
    x"2A812D58",
    x"2A811D33",
    x"2A810D11",
    x"2A80FCF0",
    x"2A80ECD1",
    x"2A80DCB5",
    x"2A80CC9A",
    x"2A80BC82",
    x"2A80AC6B",
    x"2A809C57",
    x"2A808C44",
    x"2A807C33",
    x"2A806C25",
    x"2A805C18",
    x"2A804C0E",
    x"2A803C05",
    x"2A802BFF",
    x"2A801BFA",
    x"2A800BF8",
    x"2A7FF7EF",
    x"2A7FD7F2",
    x"2A7FB7F9",
    x"2A7F9804",
    x"2A7F7813",
    x"2A7F5826",
    x"2A7F383D",
    x"2A7F1858",
    x"2A7EF877",
    x"2A7ED89A",
    x"2A7EB8C1",
    x"2A7E98EB",
    x"2A7E791A",
    x"2A7E594D",
    x"2A7E3984",
    x"2A7E19BF",
    x"2A7DF9FE",
    x"2A7DDA40",
    x"2A7DBA87",
    x"2A7D9AD2",
    x"2A7D7B20",
    x"2A7D5B73",
    x"2A7D3BC9",
    x"2A7D1C24",
    x"2A7CFC82",
    x"2A7CDCE5",
    x"2A7CBD4B",
    x"2A7C9DB5",
    x"2A7C7E24",
    x"2A7C5E96",
    x"2A7C3F0C",
    x"2A7C1F86",
    x"2A7C0004",
    x"2A7BE086",
    x"2A7BC10C",
    x"2A7BA196",
    x"2A7B8224",
    x"2A7B62B5",
    x"2A7B434B",
    x"2A7B23E5",
    x"2A7B0482",
    x"2A7AE523",
    x"2A7AC5C9",
    x"2A7AA672",
    x"2A7A871F",
    x"2A7A67D0",
    x"2A7A4885",
    x"2A7A293E",
    x"2A7A09FB",
    x"2A79EABC",
    x"2A79CB80",
    x"2A79AC49",
    x"2A798D15",
    x"2A796DE5",
    x"2A794EBA",
    x"2A792F92",
    x"2A79106E",
    x"2A78F14E",
    x"2A78D231",
    x"2A78B319",
    x"2A789405",
    x"2A7874F4",
    x"2A7855E7",
    x"2A7836DF",
    x"2A7817DA",
    x"2A77F8D9",
    x"2A77D9DB",
    x"2A77BAE2",
    x"2A779BED",
    x"2A777CFB",
    x"2A775E0D",
    x"2A773F24",
    x"2A77203E",
    x"2A77015C",
    x"2A76E27D",
    x"2A76C3A3",
    x"2A76A4CC",
    x"2A7685FA",
    x"2A76672B",
    x"2A764860",
    x"2A762999",
    x"2A760AD6",
    x"2A75EC16",
    x"2A75CD5B",
    x"2A75AEA3",
    x"2A758FEF",
    x"2A75713F",
    x"2A755293",
    x"2A7533EA",
    x"2A751546",
    x"2A74F6A5",
    x"2A74D808",
    x"2A74B96F",
    x"2A749ADA",
    x"2A747C48",
    x"2A745DBB",
    x"2A743F31",
    x"2A7420AB",
    x"2A740229",
    x"2A73E3AA",
    x"2A73C530",
    x"2A73A6B9",
    x"2A738846",
    x"2A7369D7",
    x"2A734B6B",
    x"2A732D04",
    x"2A730EA0",
    x"2A72F040",
    x"2A72D1E4",
    x"2A72B38C",
    x"2A729537",
    x"2A7276E7",
    x"2A72589A",
    x"2A723A50",
    x"2A721C0B",
    x"2A71FDC9",
    x"2A71DF8C",
    x"2A71C151",
    x"2A71A31B",
    x"2A7184E9",
    x"2A7166BA",
    x"2A71488F",
    x"2A712A68",
    x"2A710C44",
    x"2A70EE25",
    x"2A70D009",
    x"2A70B1F1",
    x"2A7093DC",
    x"2A7075CC",
    x"2A7057BF",
    x"2A7039B6",
    x"2A701BB1",
    x"2A6FFDAF",
    x"2A6FDFB1",
    x"2A6FC1B7",
    x"2A6FA3C1",
    x"2A6F85CE",
    x"2A6F67DF",
    x"2A6F49F4",
    x"2A6F2C0D",
    x"2A6F0E29",
    x"2A6EF049",
    x"2A6ED26D",
    x"2A6EB495",
    x"2A6E96C0",
    x"2A6E78EF",
    x"2A6E5B22",
    x"2A6E3D58",
    x"2A6E1F92",
    x"2A6E01D0",
    x"2A6DE412",
    x"2A6DC657",
    x"2A6DA8A0",
    x"2A6D8AED",
    x"2A6D6D3E",
    x"2A6D4F92",
    x"2A6D31EA",
    x"2A6D1445",
    x"2A6CF6A5",
    x"2A6CD908",
    x"2A6CBB6E",
    x"2A6C9DD9",
    x"2A6C8047",
    x"2A6C62B9",
    x"2A6C452E",
    x"2A6C27A7",
    x"2A6C0A24",
    x"2A6BECA5",
    x"2A6BCF29",
    x"2A6BB1B1",
    x"2A6B943D",
    x"2A6B76CC",
    x"2A6B595F",
    x"2A6B3BF6",
    x"2A6B1E90",
    x"2A6B012E",
    x"2A6AE3D0",
    x"2A6AC675",
    x"2A6AA91E",
    x"2A6A8BCB",
    x"2A6A6E7B",
    x"2A6A512F",
    x"2A6A33E7",
    x"2A6A16A2",
    x"2A69F961",
    x"2A69DC24",
    x"2A69BEEA",
    x"2A69A1B4",
    x"2A698482",
    x"2A696753",
    x"2A694A28",
    x"2A692D00",
    x"2A690FDD",
    x"2A68F2BC",
    x"2A68D5A0",
    x"2A68B887",
    x"2A689B72",
    x"2A687E60",
    x"2A686152",
    x"2A684448",
    x"2A682741",
    x"2A680A3E",
    x"2A67ED3F",
    x"2A67D043",
    x"2A67B34A",
    x"2A679656",
    x"2A677965",
    x"2A675C78",
    x"2A673F8E",
    x"2A6722A8",
    x"2A6705C5",
    x"2A66E8E6",
    x"2A66CC0B",
    x"2A66AF33",
    x"2A66925F",
    x"2A66758F",
    x"2A6658C2",
    x"2A663BF8",
    x"2A661F33",
    x"2A660271",
    x"2A65E5B2",
    x"2A65C8F7",
    x"2A65AC40",
    x"2A658F8C",
    x"2A6572DC",
    x"2A65562F",
    x"2A653986",
    x"2A651CE1",
    x"2A65003F",
    x"2A64E3A1",
    x"2A64C706",
    x"2A64AA6F",
    x"2A648DDC",
    x"2A64714C",
    x"2A6454BF",
    x"2A643837",
    x"2A641BB1",
    x"2A63FF30",
    x"2A63E2B2",
    x"2A63C637",
    x"2A63A9C0",
    x"2A638D4D",
    x"2A6370DD",
    x"2A635470",
    x"2A633808",
    x"2A631BA2",
    x"2A62FF41",
    x"2A62E2E2",
    x"2A62C688",
    x"2A62AA31",
    x"2A628DDD",
    x"2A62718D",
    x"2A625541",
    x"2A6238F8",
    x"2A621CB3",
    x"2A620071",
    x"2A61E433",
    x"2A61C7F8",
    x"2A61ABC1",
    x"2A618F8D",
    x"2A61735D",
    x"2A615730",
    x"2A613B07",
    x"2A611EE1",
    x"2A6102BF",
    x"2A60E6A1",
    x"2A60CA86",
    x"2A60AE6E",
    x"2A60925A",
    x"2A607649",
    x"2A605A3C",
    x"2A603E33",
    x"2A60222D",
    x"2A60062A",
    x"2A5FEA2B",
    x"2A5FCE30",
    x"2A5FB238",
    x"2A5F9643",
    x"2A5F7A52",
    x"2A5F5E65",
    x"2A5F427B",
    x"2A5F2694",
    x"2A5F0AB1",
    x"2A5EEED1",
    x"2A5ED2F5",
    x"2A5EB71D",
    x"2A5E9B47",
    x"2A5E7F76",
    x"2A5E63A8",
    x"2A5E47DD",
    x"2A5E2C16",
    x"2A5E1052",
    x"2A5DF492",
    x"2A5DD8D5",
    x"2A5DBD1B",
    x"2A5DA165",
    x"2A5D85B3",
    x"2A5D6A04",
    x"2A5D4E58",
    x"2A5D32B0",
    x"2A5D170C",
    x"2A5CFB6B",
    x"2A5CDFCD",
    x"2A5CC433",
    x"2A5CA89C",
    x"2A5C8D09",
    x"2A5C7179",
    x"2A5C55EC",
    x"2A5C3A63",
    x"2A5C1EDE",
    x"2A5C035B",
    x"2A5BE7DD",
    x"2A5BCC61",
    x"2A5BB0EA",
    x"2A5B9575",
    x"2A5B7A04",
    x"2A5B5E97",
    x"2A5B432D",
    x"2A5B27C6",
    x"2A5B0C63",
    x"2A5AF103",
    x"2A5AD5A6",
    x"2A5ABA4D",
    x"2A5A9EF8",
    x"2A5A83A6",
    x"2A5A6857",
    x"2A5A4D0C",
    x"2A5A31C4",
    x"2A5A167F",
    x"2A59FB3E",
    x"2A59E000",
    x"2A59C4C6",
    x"2A59A98F",
    x"2A598E5C",
    x"2A59732C",
    x"2A5957FF",
    x"2A593CD6",
    x"2A5921B0",
    x"2A59068D",
    x"2A58EB6E",
    x"2A58D052",
    x"2A58B53A",
    x"2A589A25",
    x"2A587F13",
    x"2A586405",
    x"2A5848FA",
    x"2A582DF3",
    x"2A5812EF",
    x"2A57F7EE",
    x"2A57DCF1",
    x"2A57C1F7",
    x"2A57A700",
    x"2A578C0D",
    x"2A57711D",
    x"2A575631",
    x"2A573B48",
    x"2A572062",
    x"2A570580",
    x"2A56EAA1",
    x"2A56CFC5",
    x"2A56B4ED",
    x"2A569A18",
    x"2A567F46",
    x"2A566478",
    x"2A5649AD",
    x"2A562EE6",
    x"2A561421",
    x"2A55F961",
    x"2A55DEA3",
    x"2A55C3E9",
    x"2A55A932",
    x"2A558E7F",
    x"2A5573CF",
    x"2A555922",
    x"2A553E78",
    x"2A5523D2",
    x"2A55092F",
    x"2A54EE90",
    x"2A54D3F4",
    x"2A54B95B",
    x"2A549EC5",
    x"2A548433",
    x"2A5469A4",
    x"2A544F19",
    x"2A543490",
    x"2A541A0C",
    x"2A53FF8A",
    x"2A53E50C",
    x"2A53CA91",
    x"2A53B019",
    x"2A5395A5",
    x"2A537B34",
    x"2A5360C6",
    x"2A53465B",
    x"2A532BF4",
    x"2A531190",
    x"2A52F730",
    x"2A52DCD3",
    x"2A52C279",
    x"2A52A822",
    x"2A528DCF",
    x"2A52737F",
    x"2A525932",
    x"2A523EE8",
    x"2A5224A2",
    x"2A520A5F",
    x"2A51F01F",
    x"2A51D5E3",
    x"2A51BBAA",
    x"2A51A174",
    x"2A518742",
    x"2A516D12",
    x"2A5152E6",
    x"2A5138BE",
    x"2A511E98",
    x"2A510476",
    x"2A50EA57",
    x"2A50D03B",
    x"2A50B623",
    x"2A509C0E",
    x"2A5081FC",
    x"2A5067ED",
    x"2A504DE2",
    x"2A5033DA",
    x"2A5019D5",
    x"2A4FFFD3",
    x"2A4FE5D5",
    x"2A4FCBDA",
    x"2A4FB1E2",
    x"2A4F97ED",
    x"2A4F7DFC",
    x"2A4F640E",
    x"2A4F4A23",
    x"2A4F303B",
    x"2A4F1657",
    x"2A4EFC76",
    x"2A4EE298",
    x"2A4EC8BD",
    x"2A4EAEE6",
    x"2A4E9511",
    x"2A4E7B40",
    x"2A4E6173",
    x"2A4E47A8",
    x"2A4E2DE1",
    x"2A4E141D",
    x"2A4DFA5C",
    x"2A4DE09E",
    x"2A4DC6E4",
    x"2A4DAD2C",
    x"2A4D9378",
    x"2A4D79C7",
    x"2A4D601A",
    x"2A4D466F",
    x"2A4D2CC8",
    x"2A4D1324",
    x"2A4CF983",
    x"2A4CDFE6",
    x"2A4CC64B",
    x"2A4CACB4",
    x"2A4C9320",
    x"2A4C7990",
    x"2A4C6002",
    x"2A4C4678",
    x"2A4C2CF0",
    x"2A4C136C",
    x"2A4BF9EB",
    x"2A4BE06E",
    x"2A4BC6F3",
    x"2A4BAD7C",
    x"2A4B9408",
    x"2A4B7A97",
    x"2A4B6129",
    x"2A4B47BF",
    x"2A4B2E57",
    x"2A4B14F3",
    x"2A4AFB92",
    x"2A4AE234",
    x"2A4AC8DA",
    x"2A4AAF82",
    x"2A4A962E",
    x"2A4A7CDD",
    x"2A4A638E",
    x"2A4A4A44",
    x"2A4A30FC",
    x"2A4A17B7",
    x"2A49FE76",
    x"2A49E538",
    x"2A49CBFD",
    x"2A49B2C5",
    x"2A499990",
    x"2A49805E",
    x"2A496730",
    x"2A494E05",
    x"2A4934DC",
    x"2A491BB7",
    x"2A490295",
    x"2A48E977",
    x"2A48D05B",
    x"2A48B743",
    x"2A489E2D",
    x"2A48851B",
    x"2A486C0C",
    x"2A485300",
    x"2A4839F7",
    x"2A4820F2",
    x"2A4807EF",
    x"2A47EEF0",
    x"2A47D5F3",
    x"2A47BCFA",
    x"2A47A404",
    x"2A478B11",
    x"2A477221",
    x"2A475935",
    x"2A47404B",
    x"2A472764",
    x"2A470E81",
    x"2A46F5A1",
    x"2A46DCC4",
    x"2A46C3EA",
    x"2A46AB13",
    x"2A46923F",
    x"2A46796E",
    x"2A4660A1",
    x"2A4647D6",
    x"2A462F0F",
    x"2A46164A",
    x"2A45FD89",
    x"2A45E4CB",
    x"2A45CC10",
    x"2A45B358",
    x"2A459AA3",
    x"2A4581F1",
    x"2A456942",
    x"2A455097",
    x"2A4537EE",
    x"2A451F49",
    x"2A4506A7",
    x"2A44EE07",
    x"2A44D56B",
    x"2A44BCD2",
    x"2A44A43C",
    x"2A448BA9",
    x"2A447319",
    x"2A445A8C",
    x"2A444202",
    x"2A44297C",
    x"2A4410F8",
    x"2A43F877",
    x"2A43DFFA",
    x"2A43C77F",
    x"2A43AF08",
    x"2A439694",
    x"2A437E22",
    x"2A4365B4",
    x"2A434D49",
    x"2A4334E1",
    x"2A431C7C",
    x"2A43041A",
    x"2A42EBBB",
    x"2A42D35F",
    x"2A42BB06",
    x"2A42A2B0",
    x"2A428A5D",
    x"2A42720D",
    x"2A4259C1",
    x"2A424177",
    x"2A422930",
    x"2A4210ED",
    x"2A41F8AC",
    x"2A41E06E",
    x"2A41C834",
    x"2A41AFFC",
    x"2A4197C8",
    x"2A417F96",
    x"2A416768",
    x"2A414F3D",
    x"2A413714",
    x"2A411EEF",
    x"2A4106CC",
    x"2A40EEAD",
    x"2A40D691",
    x"2A40BE77",
    x"2A40A661",
    x"2A408E4E",
    x"2A40763E",
    x"2A405E30",
    x"2A404626",
    x"2A402E1F",
    x"2A40161A",
    x"2A3FFE19",
    x"2A3FE61B",
    x"2A3FCE20",
    x"2A3FB627",
    x"2A3F9E32",
    x"2A3F8640",
    x"2A3F6E51",
    x"2A3F5664",
    x"2A3F3E7B",
    x"2A3F2695",
    x"2A3F0EB1",
    x"2A3EF6D1",
    x"2A3EDEF4",
    x"2A3EC719",
    x"2A3EAF42",
    x"2A3E976D",
    x"2A3E7F9C",
    x"2A3E67CE",
    x"2A3E5002",
    x"2A3E383A",
    x"2A3E2074",
    x"2A3E08B1",
    x"2A3DF0F2",
    x"2A3DD935",
    x"2A3DC17C",
    x"2A3DA9C5",
    x"2A3D9211",
    x"2A3D7A60",
    x"2A3D62B2",
    x"2A3D4B08",
    x"2A3D3360",
    x"2A3D1BBB",
    x"2A3D0419",
    x"2A3CEC7A",
    x"2A3CD4DE",
    x"2A3CBD45",
    x"2A3CA5AE",
    x"2A3C8E1B",
    x"2A3C768B",
    x"2A3C5EFD",
    x"2A3C4773",
    x"2A3C2FEC",
    x"2A3C1867",
    x"2A3C00E6",
    x"2A3BE967",
    x"2A3BD1EB",
    x"2A3BBA72",
    x"2A3BA2FD",
    x"2A3B8B8A",
    x"2A3B741A",
    x"2A3B5CAD",
    x"2A3B4542",
    x"2A3B2DDB",
    x"2A3B1677",
    x"2A3AFF16",
    x"2A3AE7B7",
    x"2A3AD05C",
    x"2A3AB903",
    x"2A3AA1AD",
    x"2A3A8A5B",
    x"2A3A730B",
    x"2A3A5BBE",
    x"2A3A4474",
    x"2A3A2D2D",
    x"2A3A15E9",
    x"2A39FEA7",
    x"2A39E769",
    x"2A39D02E",
    x"2A39B8F5",
    x"2A39A1BF",
    x"2A398A8D",
    x"2A39735D",
    x"2A395C30",
    x"2A394506",
    x"2A392DDE",
    x"2A3916BA",
    x"2A38FF99",
    x"2A38E87A",
    x"2A38D15F",
    x"2A38BA46",
    x"2A38A330",
    x"2A388C1D",
    x"2A38750D",
    x"2A385E00",
    x"2A3846F6",
    x"2A382FEE",
    x"2A3818EA",
    x"2A3801E8",
    x"2A37EAE9",
    x"2A37D3ED",
    x"2A37BCF4",
    x"2A37A5FE",
    x"2A378F0B",
    x"2A37781A",
    x"2A37612D",
    x"2A374A42",
    x"2A37335A",
    x"2A371C75",
    x"2A370593",
    x"2A36EEB4",
    x"2A36D7D7",
    x"2A36C0FE",
    x"2A36AA27",
    x"2A369353",
    x"2A367C82",
    x"2A3665B4",
    x"2A364EE9",
    x"2A363820",
    x"2A36215B",
    x"2A360A98",
    x"2A35F3D8",
    x"2A35DD1B",
    x"2A35C661",
    x"2A35AFA9",
    x"2A3598F5",
    x"2A358243",
    x"2A356B94",
    x"2A3554E8",
    x"2A353E3F",
    x"2A352799",
    x"2A3510F5",
    x"2A34FA54",
    x"2A34E3B7",
    x"2A34CD1C",
    x"2A34B683",
    x"2A349FEE",
    x"2A34895B",
    x"2A3472CC",
    x"2A345C3F",
    x"2A3445B4",
    x"2A342F2D",
    x"2A3418A9",
    x"2A340227",
    x"2A33EBA8",
    x"2A33D52C",
    x"2A33BEB3",
    x"2A33A83C",
    x"2A3391C9",
    x"2A337B58",
    x"2A3364EA",
    x"2A334E7F",
    x"2A333816",
    x"2A3321B1",
    x"2A330B4E",
    x"2A32F4EE",
    x"2A32DE91",
    x"2A32C836",
    x"2A32B1DF",
    x"2A329B8A",
    x"2A328538",
    x"2A326EE8",
    x"2A32589C",
    x"2A324252",
    x"2A322C0B",
    x"2A3215C7",
    x"2A31FF86",
    x"2A31E947",
    x"2A31D30C",
    x"2A31BCD3",
    x"2A31A69C",
    x"2A319069",
    x"2A317A38",
    x"2A31640A",
    x"2A314DDF",
    x"2A3137B7",
    x"2A312191",
    x"2A310B6F",
    x"2A30F54F",
    x"2A30DF31",
    x"2A30C917",
    x"2A30B2FF",
    x"2A309CEA",
    x"2A3086D8",
    x"2A3070C8",
    x"2A305ABC",
    x"2A3044B2",
    x"2A302EAA",
    x"2A3018A6",
    x"2A3002A4",
    x"2A2FECA5",
    x"2A2FD6A9",
    x"2A2FC0B0",
    x"2A2FAAB9",
    x"2A2F94C5",
    x"2A2F7ED4",
    x"2A2F68E5",
    x"2A2F52F9",
    x"2A2F3D10",
    x"2A2F272A",
    x"2A2F1147",
    x"2A2EFB66",
    x"2A2EE588",
    x"2A2ECFAD",
    x"2A2EB9D4",
    x"2A2EA3FE",
    x"2A2E8E2B",
    x"2A2E785B",
    x"2A2E628D",
    x"2A2E4CC2",
    x"2A2E36FA",
    x"2A2E2134",
    x"2A2E0B71",
    x"2A2DF5B1",
    x"2A2DDFF4",
    x"2A2DCA39",
    x"2A2DB481",
    x"2A2D9ECC",
    x"2A2D891A",
    x"2A2D736A",
    x"2A2D5DBD",
    x"2A2D4812",
    x"2A2D326B",
    x"2A2D1CC6",
    x"2A2D0724",
    x"2A2CF184",
    x"2A2CDBE7",
    x"2A2CC64D",
    x"2A2CB0B6",
    x"2A2C9B21",
    x"2A2C858F",
    x"2A2C7000",
    x"2A2C5A73",
    x"2A2C44E9",
    x"2A2C2F62",
    x"2A2C19DD",
    x"2A2C045B",
    x"2A2BEEDC",
    x"2A2BD95F",
    x"2A2BC3E6",
    x"2A2BAE6E",
    x"2A2B98FA",
    x"2A2B8388",
    x"2A2B6E19",
    x"2A2B58AD",
    x"2A2B4343",
    x"2A2B2DDC",
    x"2A2B1877",
    x"2A2B0316",
    x"2A2AEDB7",
    x"2A2AD85A",
    x"2A2AC301",
    x"2A2AADAA",
    x"2A2A9855",
    x"2A2A8304",
    x"2A2A6DB4",
    x"2A2A5868",
    x"2A2A431E",
    x"2A2A2DD7",
    x"2A2A1893",
    x"2A2A0351",
    x"2A29EE12",
    x"2A29D8D6",
    x"2A29C39C",
    x"2A29AE65",
    x"2A299930",
    x"2A2983FE",
    x"2A296ECF",
    x"2A2959A3",
    x"2A294479",
    x"2A292F52",
    x"2A291A2D",
    x"2A29050B",
    x"2A28EFEC",
    x"2A28DACF",
    x"2A28C5B5",
    x"2A28B09E",
    x"2A289B89",
    x"2A288677",
    x"2A287167",
    x"2A285C5A",
    x"2A284750",
    x"2A283249",
    x"2A281D44",
    x"2A280841",
    x"2A27F342",
    x"2A27DE44",
    x"2A27C94A",
    x"2A27B452",
    x"2A279F5D",
    x"2A278A6A",
    x"2A27757A",
    x"2A27608D",
    x"2A274BA2",
    x"2A2736BA",
    x"2A2721D4",
    x"2A270CF2",
    x"2A26F811",
    x"2A26E334",
    x"2A26CE58",
    x"2A26B980",
    x"2A26A4AA",
    x"2A268FD7",
    x"2A267B06",
    x"2A266638",
    x"2A26516D",
    x"2A263CA4",
    x"2A2627DD",
    x"2A26131A",
    x"2A25FE59",
    x"2A25E99A",
    x"2A25D4DE",
    x"2A25C025",
    x"2A25AB6E",
    x"2A2596BA",
    x"2A258209",
    x"2A256D5A",
    x"2A2558AD",
    x"2A254403",
    x"2A252F5C",
    x"2A251AB8",
    x"2A250615",
    x"2A24F176",
    x"2A24DCD9",
    x"2A24C83F",
    x"2A24B3A7",
    x"2A249F12",
    x"2A248A7F",
    x"2A2475EF",
    x"2A246162",
    x"2A244CD7",
    x"2A24384F",
    x"2A2423C9",
    x"2A240F46",
    x"2A23FAC5",
    x"2A23E647",
    x"2A23D1CB",
    x"2A23BD53",
    x"2A23A8DC",
    x"2A239468",
    x"2A237FF7",
    x"2A236B88",
    x"2A23571C",
    x"2A2342B3",
    x"2A232E4B",
    x"2A2319E7",
    x"2A230585",
    x"2A22F126",
    x"2A22DCC9",
    x"2A22C86E",
    x"2A22B417",
    x"2A229FC1",
    x"2A228B6F",
    x"2A22771E",
    x"2A2262D1",
    x"2A224E86",
    x"2A223A3D",
    x"2A2225F7",
    x"2A2211B4",
    x"2A21FD73",
    x"2A21E934",
    x"2A21D4F9",
    x"2A21C0BF",
    x"2A21AC88",
    x"2A219854",
    x"2A218422",
    x"2A216FF3",
    x"2A215BC6",
    x"2A21479C",
    x"2A213374",
    x"2A211F4F",
    x"2A210B2D",
    x"2A20F70C",
    x"2A20E2EF",
    x"2A20CED4",
    x"2A20BABB",
    x"2A20A6A5",
    x"2A209291",
    x"2A207E80",
    x"2A206A72",
    x"2A205666",
    x"2A20425C",
    x"2A202E55",
    x"2A201A51",
    x"2A20064F",
    x"2A1FF24F",
    x"2A1FDE52",
    x"2A1FCA57",
    x"2A1FB65F",
    x"2A1FA26A",
    x"2A1F8E77",
    x"2A1F7A86",
    x"2A1F6698",
    x"2A1F52AD",
    x"2A1F3EC3",
    x"2A1F2ADD",
    x"2A1F16F9",
    x"2A1F0317",
    x"2A1EEF38",
    x"2A1EDB5B",
    x"2A1EC781",
    x"2A1EB3A9",
    x"2A1E9FD4",
    x"2A1E8C01",
    x"2A1E7831",
    x"2A1E6463",
    x"2A1E5098",
    x"2A1E3CCF",
    x"2A1E2909",
    x"2A1E1545",
    x"2A1E0184",
    x"2A1DEDC5",
    x"2A1DDA08",
    x"2A1DC64E",
    x"2A1DB297",
    x"2A1D9EE1",
    x"2A1D8B2F",
    x"2A1D777F",
    x"2A1D63D1",
    x"2A1D5026",
    x"2A1D3C7D",
    x"2A1D28D7",
    x"2A1D1533",
    x"2A1D0191",
    x"2A1CEDF2",
    x"2A1CDA56",
    x"2A1CC6BC",
    x"2A1CB324",
    x"2A1C9F8F",
    x"2A1C8BFC",
    x"2A1C786C",
    x"2A1C64DE",
    x"2A1C5153",
    x"2A1C3DCA",
    x"2A1C2A43",
    x"2A1C16BF",
    x"2A1C033E",
    x"2A1BEFBE",
    x"2A1BDC42",
    x"2A1BC8C7",
    x"2A1BB550",
    x"2A1BA1DA",
    x"2A1B8E67",
    x"2A1B7AF6",
    x"2A1B6788",
    x"2A1B541D",
    x"2A1B40B3",
    x"2A1B2D4C",
    x"2A1B19E8",
    x"2A1B0686",
    x"2A1AF326",
    x"2A1ADFC9",
    x"2A1ACC6E",
    x"2A1AB916",
    x"2A1AA5C0",
    x"2A1A926D",
    x"2A1A7F1B",
    x"2A1A6BCD",
    x"2A1A5881",
    x"2A1A4537",
    x"2A1A31EF",
    x"2A1A1EAA",
    x"2A1A0B68",
    x"2A19F827",
    x"2A19E4EA",
    x"2A19D1AE",
    x"2A19BE75",
    x"2A19AB3F",
    x"2A19980A",
    x"2A1984D8",
    x"2A1971A9",
    x"2A195E7C",
    x"2A194B51",
    x"2A193829",
    x"2A192503",
    x"2A1911E0",
    x"2A18FEBF",
    x"2A18EBA0",
    x"2A18D884",
    x"2A18C56A",
    x"2A18B253",
    x"2A189F3E",
    x"2A188C2B",
    x"2A18791B",
    x"2A18660D",
    x"2A185301",
    x"2A183FF8",
    x"2A182CF1",
    x"2A1819ED",
    x"2A1806EB",
    x"2A17F3EB",
    x"2A17E0EE",
    x"2A17CDF3",
    x"2A17BAFA",
    x"2A17A804",
    x"2A179510",
    x"2A17821F",
    x"2A176F30",
    x"2A175C43",
    x"2A174959",
    x"2A173671",
    x"2A17238B",
    x"2A1710A8",
    x"2A16FDC7",
    x"2A16EAE8",
    x"2A16D80C",
    x"2A16C532",
    x"2A16B25B",
    x"2A169F86",
    x"2A168CB3",
    x"2A1679E2",
    x"2A166714",
    x"2A165449",
    x"2A16417F",
    x"2A162EB8",
    x"2A161BF4",
    x"2A160931",
    x"2A15F671",
    x"2A15E3B4",
    x"2A15D0F8",
    x"2A15BE3F",
    x"2A15AB89",
    x"2A1598D5",
    x"2A158623",
    x"2A157373",
    x"2A1560C6",
    x"2A154E1B",
    x"2A153B72",
    x"2A1528CC",
    x"2A151628",
    x"2A150386",
    x"2A14F0E7",
    x"2A14DE4A",
    x"2A14CBB0",
    x"2A14B917",
    x"2A14A681",
    x"2A1493EE",
    x"2A14815C",
    x"2A146ECD",
    x"2A145C41",
    x"2A1449B6",
    x"2A14372E",
    x"2A1424A8",
    x"2A141225",
    x"2A13FFA4",
    x"2A13ED25",
    x"2A13DAA9",
    x"2A13C82E",
    x"2A13B5B7",
    x"2A13A341",
    x"2A1390CE",
    x"2A137E5D",
    x"2A136BEE",
    x"2A135982",
    x"2A134718",
    x"2A1334B0",
    x"2A13224B",
    x"2A130FE7",
    x"2A12FD87",
    x"2A12EB28",
    x"2A12D8CC",
    x"2A12C672",
    x"2A12B41A",
    x"2A12A1C5",
    x"2A128F72",
    x"2A127D21",
    x"2A126AD3",
    x"2A125886",
    x"2A12463C",
    x"2A1233F5",
    x"2A1221AF",
    x"2A120F6C",
    x"2A11FD2C",
    x"2A11EAED",
    x"2A11D8B1",
    x"2A11C677",
    x"2A11B43F",
    x"2A11A20A",
    x"2A118FD7",
    x"2A117DA6",
    x"2A116B77",
    x"2A11594B",
    x"2A114721",
    x"2A1134F9",
    x"2A1122D4",
    x"2A1110B0",
    x"2A10FE90",
    x"2A10EC71",
    x"2A10DA54",
    x"2A10C83A",
    x"2A10B622",
    x"2A10A40D",
    x"2A1091F9",
    x"2A107FE8",
    x"2A106DD9",
    x"2A105BCD",
    x"2A1049C2",
    x"2A1037BA",
    x"2A1025B4",
    x"2A1013B1",
    x"2A1001B0",
    x"2A0FEFB0",
    x"2A0FDDB4",
    x"2A0FCBB9",
    x"2A0FB9C1",
    x"2A0FA7CB",
    x"2A0F95D7",
    x"2A0F83E5",
    x"2A0F71F6",
    x"2A0F6009",
    x"2A0F4E1E",
    x"2A0F3C35",
    x"2A0F2A4F",
    x"2A0F186B",
    x"2A0F0689",
    x"2A0EF4A9",
    x"2A0EE2CB",
    x"2A0ED0F0",
    x"2A0EBF17",
    x"2A0EAD40",
    x"2A0E9B6C",
    x"2A0E899A",
    x"2A0E77CA",
    x"2A0E65FC",
    x"2A0E5430",
    x"2A0E4267",
    x"2A0E309F",
    x"2A0E1EDA",
    x"2A0E0D18",
    x"2A0DFB57",
    x"2A0DE999",
    x"2A0DD7DD",
    x"2A0DC623",
    x"2A0DB46B",
    x"2A0DA2B6",
    x"2A0D9103",
    x"2A0D7F52",
    x"2A0D6DA3",
    x"2A0D5BF6",
    x"2A0D4A4C",
    x"2A0D38A4",
    x"2A0D26FE",
    x"2A0D155A",
    x"2A0D03B8",
    x"2A0CF219",
    x"2A0CE07C",
    x"2A0CCEE1",
    x"2A0CBD48",
    x"2A0CABB1",
    x"2A0C9A1D",
    x"2A0C888B",
    x"2A0C76FB",
    x"2A0C656D",
    x"2A0C53E2",
    x"2A0C4258",
    x"2A0C30D1",
    x"2A0C1F4C",
    x"2A0C0DC9",
    x"2A0BFC49",
    x"2A0BEACA",
    x"2A0BD94E",
    x"2A0BC7D4",
    x"2A0BB65C",
    x"2A0BA4E6",
    x"2A0B9373",
    x"2A0B8201",
    x"2A0B7092",
    x"2A0B5F25",
    x"2A0B4DBA",
    x"2A0B3C52",
    x"2A0B2AEB",
    x"2A0B1987",
    x"2A0B0825",
    x"2A0AF6C5",
    x"2A0AE567",
    x"2A0AD40C",
    x"2A0AC2B2",
    x"2A0AB15B",
    x"2A0AA006",
    x"2A0A8EB3",
    x"2A0A7D62",
    x"2A0A6C14",
    x"2A0A5AC7",
    x"2A0A497D",
    x"2A0A3835",
    x"2A0A26EF",
    x"2A0A15AB",
    x"2A0A0469",
    x"2A09F32A",
    x"2A09E1ED",
    x"2A09D0B1",
    x"2A09BF78",
    x"2A09AE42",
    x"2A099D0D",
    x"2A098BDA",
    x"2A097AAA",
    x"2A09697C",
    x"2A095850",
    x"2A094726",
    x"2A0935FE",
    x"2A0924D8",
    x"2A0913B5",
    x"2A090293",
    x"2A08F174",
    x"2A08E057",
    x"2A08CF3C",
    x"2A08BE23",
    x"2A08AD0C",
    x"2A089BF8",
    x"2A088AE5",
    x"2A0879D5",
    x"2A0868C7",
    x"2A0857BB",
    x"2A0846B1",
    x"2A0835A9",
    x"2A0824A4",
    x"2A0813A0",
    x"2A08029F",
    x"2A07F19F",
    x"2A07E0A2",
    x"2A07CFA7",
    x"2A07BEAE",
    x"2A07ADB8",
    x"2A079CC3",
    x"2A078BD0",
    x"2A077AE0",
    x"2A0769F2",
    x"2A075905",
    x"2A07481B",
    x"2A073733",
    x"2A07264E",
    x"2A07156A",
    x"2A070488",
    x"2A06F3A9",
    x"2A06E2CB",
    x"2A06D1F0",
    x"2A06C117",
    x"2A06B040",
    x"2A069F6B",
    x"2A068E98",
    x"2A067DC7",
    x"2A066CF8",
    x"2A065C2C",
    x"2A064B61",
    x"2A063A99",
    x"2A0629D3",
    x"2A06190F",
    x"2A06084C",
    x"2A05F78C",
    x"2A05E6CF",
    x"2A05D613",
    x"2A05C559",
    x"2A05B4A1",
    x"2A05A3EC",
    x"2A059338",
    x"2A058287",
    x"2A0571D8",
    x"2A05612B",
    x"2A055080",
    x"2A053FD6",
    x"2A052F30",
    x"2A051E8B",
    x"2A050DE8",
    x"2A04FD47",
    x"2A04ECA9",
    x"2A04DC0C",
    x"2A04CB72",
    x"2A04BAD9",
    x"2A04AA43",
    x"2A0499AF",
    x"2A04891C",
    x"2A04788C",
    x"2A0467FE",
    x"2A045772",
    x"2A0446E8",
    x"2A043661",
    x"2A0425DB",
    x"2A041557",
    x"2A0404D6",
    x"2A03F456",
    x"2A03E3D8",
    x"2A03D35D",
    x"2A03C2E4",
    x"2A03B26C",
    x"2A03A1F7",
    x"2A039184",
    x"2A038113",
    x"2A0370A3",
    x"2A036036",
    x"2A034FCB",
    x"2A033F62",
    x"2A032EFC",
    x"2A031E97",
    x"2A030E34",
    x"2A02FDD3",
    x"2A02ED74",
    x"2A02DD18",
    x"2A02CCBD",
    x"2A02BC65",
    x"2A02AC0E",
    x"2A029BBA",
    x"2A028B67",
    x"2A027B17",
    x"2A026AC8",
    x"2A025A7C",
    x"2A024A32",
    x"2A0239EA",
    x"2A0229A3",
    x"2A02195F",
    x"2A02091D",
    x"2A01F8DD",
    x"2A01E89F",
    x"2A01D863",
    x"2A01C829",
    x"2A01B7F1",
    x"2A01A7BB",
    x"2A019787",
    x"2A018755",
    x"2A017725",
    x"2A0166F7",
    x"2A0156CB",
    x"2A0146A1",
    x"2A013679",
    x"2A012654",
    x"2A011630",
    x"2A01060E",
    x"2A00F5EE",
    x"2A00E5D1",
    x"2A00D5B5",
    x"2A00C59B",
    x"2A00B584",
    x"2A00A56E",
    x"2A00955A",
    x"2A008549",
    x"2A007539",
    x"2A00652B",
    x"2A005520",
    x"2A004516",
    x"2A00350E",
    x"2A002509",
    x"2A001505",
    x"2A000503",
    x"29FFEA08",
    x"29FFCA0C",
    x"29FFAA15",
    x"29FF8A22",
    x"29FF6A33",
    x"29FF4A47",
    x"29FF2A60",
    x"29FF0A7D",
    x"29FEEA9D",
    x"29FECAC2",
    x"29FEAAEB",
    x"29FE8B17",
    x"29FE6B48",
    x"29FE4B7C",
    x"29FE2BB5",
    x"29FE0BF2",
    x"29FDEC32",
    x"29FDCC76",
    x"29FDACBF",
    x"29FD8D0B",
    x"29FD6D5C",
    x"29FD4DB0",
    x"29FD2E08",
    x"29FD0E64",
    x"29FCEEC5",
    x"29FCCF29",
    x"29FCAF91",
    x"29FC8FFD",
    x"29FC706D",
    x"29FC50E1",
    x"29FC3159",
    x"29FC11D4",
    x"29FBF254",
    x"29FBD2D8",
    x"29FBB35F",
    x"29FB93EB",
    x"29FB747A",
    x"29FB550E",
    x"29FB35A5",
    x"29FB1640",
    x"29FAF6E0",
    x"29FAD783",
    x"29FAB82A",
    x"29FA98D5",
    x"29FA7984",
    x"29FA5A36",
    x"29FA3AED",
    x"29FA1BA8",
    x"29F9FC66",
    x"29F9DD28",
    x"29F9BDEF",
    x"29F99EB9",
    x"29F97F87",
    x"29F96059",
    x"29F9412F",
    x"29F92209",
    x"29F902E7",
    x"29F8E3C8",
    x"29F8C4AE",
    x"29F8A597",
    x"29F88684",
    x"29F86775",
    x"29F8486A",
    x"29F82963",
    x"29F80A60",
    x"29F7EB61",
    x"29F7CC65",
    x"29F7AD6D",
    x"29F78E7A",
    x"29F76F8A",
    x"29F7509E",
    x"29F731B6",
    x"29F712D1",
    x"29F6F3F1",
    x"29F6D514",
    x"29F6B63C",
    x"29F69767",
    x"29F67896",
    x"29F659C9",
    x"29F63AFF",
    x"29F61C3A",
    x"29F5FD78",
    x"29F5DEBB",
    x"29F5C001",
    x"29F5A14B",
    x"29F58298",
    x"29F563EA",
    x"29F5453F",
    x"29F52699",
    x"29F507F6",
    x"29F4E957",
    x"29F4CABB",
    x"29F4AC24",
    x"29F48D90",
    x"29F46F01",
    x"29F45075",
    x"29F431EC",
    x"29F41368",
    x"29F3F4E8",
    x"29F3D66B",
    x"29F3B7F2",
    x"29F3997D",
    x"29F37B0C",
    x"29F35C9E",
    x"29F33E34",
    x"29F31FCF",
    x"29F3016D",
    x"29F2E30E",
    x"29F2C4B4",
    x"29F2A65D",
    x"29F2880A",
    x"29F269BB",
    x"29F24B70",
    x"29F22D28",
    x"29F20EE4",
    x"29F1F0A4",
    x"29F1D268",
    x"29F1B430",
    x"29F195FB",
    x"29F177CA",
    x"29F1599D",
    x"29F13B74",
    x"29F11D4E",
    x"29F0FF2D",
    x"29F0E10F",
    x"29F0C2F4",
    x"29F0A4DE",
    x"29F086CB",
    x"29F068BC",
    x"29F04AB1",
    x"29F02CAA",
    x"29F00EA6",
    x"29EFF0A6",
    x"29EFD2AA",
    x"29EFB4B1",
    x"29EF96BC",
    x"29EF78CC",
    x"29EF5ADE",
    x"29EF3CF5",
    x"29EF1F0F",
    x"29EF012D",
    x"29EEE34F",
    x"29EEC574",
    x"29EEA79D",
    x"29EE89CA",
    x"29EE6BFB",
    x"29EE4E2F",
    x"29EE3067",
    x"29EE12A3",
    x"29EDF4E3",
    x"29EDD726",
    x"29EDB96D",
    x"29ED9BB8",
    x"29ED7E06",
    x"29ED6058",
    x"29ED42AE",
    x"29ED2507",
    x"29ED0765",
    x"29ECE9C6",
    x"29ECCC2A",
    x"29ECAE93",
    x"29EC90FF",
    x"29EC736E",
    x"29EC55E2",
    x"29EC3859",
    x"29EC1AD4",
    x"29EBFD52",
    x"29EBDFD4",
    x"29EBC25A",
    x"29EBA4E4",
    x"29EB8771",
    x"29EB6A02",
    x"29EB4C96",
    x"29EB2F2F",
    x"29EB11CB",
    x"29EAF46A",
    x"29EAD70E",
    x"29EAB9B4",
    x"29EA9C5F",
    x"29EA7F0D",
    x"29EA61BF",
    x"29EA4475",
    x"29EA272E",
    x"29EA09EB",
    x"29E9ECAC",
    x"29E9CF70",
    x"29E9B238",
    x"29E99503",
    x"29E977D3",
    x"29E95AA5",
    x"29E93D7C",
    x"29E92056",
    x"29E90334",
    x"29E8E615",
    x"29E8C8FA",
    x"29E8ABE3",
    x"29E88ECF",
    x"29E871BF",
    x"29E854B3",
    x"29E837AA",
    x"29E81AA5",
    x"29E7FDA4",
    x"29E7E0A6",
    x"29E7C3AB",
    x"29E7A6B5",
    x"29E789C2",
    x"29E76CD2",
    x"29E74FE6",
    x"29E732FE",
    x"29E7161A",
    x"29E6F939",
    x"29E6DC5B",
    x"29E6BF82",
    x"29E6A2AC",
    x"29E685D9",
    x"29E6690A",
    x"29E64C3F",
    x"29E62F77",
    x"29E612B3",
    x"29E5F5F2",
    x"29E5D935",
    x"29E5BC7C",
    x"29E59FC6",
    x"29E58314",
    x"29E56666",
    x"29E549BB",
    x"29E52D13",
    x"29E5106F",
    x"29E4F3CF",
    x"29E4D732",
    x"29E4BA99",
    x"29E49E04",
    x"29E48172",
    x"29E464E3",
    x"29E44858",
    x"29E42BD1",
    x"29E40F4D",
    x"29E3F2CD",
    x"29E3D651",
    x"29E3B9D8",
    x"29E39D62",
    x"29E380F0",
    x"29E36482",
    x"29E34817",
    x"29E32BB0",
    x"29E30F4C",
    x"29E2F2EC",
    x"29E2D690",
    x"29E2BA37",
    x"29E29DE1",
    x"29E2818F",
    x"29E26541",
    x"29E248F6",
    x"29E22CAE",
    x"29E2106B",
    x"29E1F42A",
    x"29E1D7EE",
    x"29E1BBB4",
    x"29E19F7F",
    x"29E1834D",
    x"29E1671E",
    x"29E14AF3",
    x"29E12ECB",
    x"29E112A7",
    x"29E0F686",
    x"29E0DA69",
    x"29E0BE50",
    x"29E0A23A",
    x"29E08627",
    x"29E06A18",
    x"29E04E0D",
    x"29E03205",
    x"29E01600",
    x"29DFF9FF",
    x"29DFDE02",
    x"29DFC208",
    x"29DFA611",
    x"29DF8A1E",
    x"29DF6E2F",
    x"29DF5243",
    x"29DF365A",
    x"29DF1A75",
    x"29DEFE94",
    x"29DEE2B5",
    x"29DEC6DB",
    x"29DEAB04",
    x"29DE8F30",
    x"29DE7360",
    x"29DE5793",
    x"29DE3BCA",
    x"29DE2004",
    x"29DE0442",
    x"29DDE883",
    x"29DDCCC8",
    x"29DDB110",
    x"29DD955C",
    x"29DD79AB",
    x"29DD5DFD",
    x"29DD4253",
    x"29DD26AD",
    x"29DD0B0A",
    x"29DCEF6A",
    x"29DCD3CE",
    x"29DCB835",
    x"29DC9CA0",
    x"29DC810E",
    x"29DC657F",
    x"29DC49F4",
    x"29DC2E6D",
    x"29DC12E9",
    x"29DBF768",
    x"29DBDBEB",
    x"29DBC071",
    x"29DBA4FB",
    x"29DB8988",
    x"29DB6E18",
    x"29DB52AC",
    x"29DB3744",
    x"29DB1BDF",
    x"29DB007D",
    x"29DAE51E",
    x"29DAC9C4",
    x"29DAAE6C",
    x"29DA9318",
    x"29DA77C7",
    x"29DA5C7A",
    x"29DA4130",
    x"29DA25EA",
    x"29DA0AA7",
    x"29D9EF67",
    x"29D9D42B",
    x"29D9B8F2",
    x"29D99DBD",
    x"29D9828B",
    x"29D9675C",
    x"29D94C31",
    x"29D93109",
    x"29D915E4",
    x"29D8FAC3",
    x"29D8DFA6",
    x"29D8C48C",
    x"29D8A975",
    x"29D88E61",
    x"29D87351",
    x"29D85844",
    x"29D83D3B",
    x"29D82235",
    x"29D80732",
    x"29D7EC33",
    x"29D7D137",
    x"29D7B63F",
    x"29D79B4A",
    x"29D78058",
    x"29D7656A",
    x"29D74A7F",
    x"29D72F97",
    x"29D714B3",
    x"29D6F9D2",
    x"29D6DEF4",
    x"29D6C41A",
    x"29D6A943",
    x"29D68E70",
    x"29D673A0",
    x"29D658D3",
    x"29D63E0A",
    x"29D62343",
    x"29D60881",
    x"29D5EDC1",
    x"29D5D305",
    x"29D5B84D",
    x"29D59D97",
    x"29D582E5",
    x"29D56836",
    x"29D54D8B",
    x"29D532E3",
    x"29D5183E",
    x"29D4FD9D",
    x"29D4E2FF",
    x"29D4C864",
    x"29D4ADCD",
    x"29D49339",
    x"29D478A8",
    x"29D45E1B",
    x"29D44391",
    x"29D4290A",
    x"29D40E86",
    x"29D3F406",
    x"29D3D989",
    x"29D3BF10",
    x"29D3A49A",
    x"29D38A27",
    x"29D36FB7",
    x"29D3554B",
    x"29D33AE2",
    x"29D3207C",
    x"29D3061A",
    x"29D2EBBA",
    x"29D2D15F",
    x"29D2B706",
    x"29D29CB1",
    x"29D2825F",
    x"29D26810",
    x"29D24DC5",
    x"29D2337D",
    x"29D21938",
    x"29D1FEF7",
    x"29D1E4B8",
    x"29D1CA7D",
    x"29D1B046",
    x"29D19611",
    x"29D17BE0",
    x"29D161B2",
    x"29D14788",
    x"29D12D60",
    x"29D1133C",
    x"29D0F91C",
    x"29D0DEFE",
    x"29D0C4E4",
    x"29D0AACD",
    x"29D090B9",
    x"29D076A9",
    x"29D05C9B",
    x"29D04292",
    x"29D0288B",
    x"29D00E87",
    x"29CFF487",
    x"29CFDA8A",
    x"29CFC091",
    x"29CFA69A",
    x"29CF8CA7",
    x"29CF72B7",
    x"29CF58CA",
    x"29CF3EE1",
    x"29CF24FB",
    x"29CF0B18",
    x"29CEF138",
    x"29CED75B",
    x"29CEBD82",
    x"29CEA3AC",
    x"29CE89D9",
    x"29CE7009",
    x"29CE563D",
    x"29CE3C74",
    x"29CE22AE",
    x"29CE08EB",
    x"29CDEF2C",
    x"29CDD56F",
    x"29CDBBB6",
    x"29CDA200",
    x"29CD884E",
    x"29CD6E9E",
    x"29CD54F2",
    x"29CD3B49",
    x"29CD21A3",
    x"29CD0801",
    x"29CCEE61",
    x"29CCD4C5",
    x"29CCBB2C",
    x"29CCA196",
    x"29CC8804",
    x"29CC6E74",
    x"29CC54E8",
    x"29CC3B5F",
    x"29CC21D9",
    x"29CC0857",
    x"29CBEED7",
    x"29CBD55B",
    x"29CBBBE2",
    x"29CBA26C",
    x"29CB88F9",
    x"29CB6F8A",
    x"29CB561D",
    x"29CB3CB4",
    x"29CB234E",
    x"29CB09EB",
    x"29CAF08C",
    x"29CAD72F",
    x"29CABDD6",
    x"29CAA480",
    x"29CA8B2D",
    x"29CA71DD",
    x"29CA5890",
    x"29CA3F47",
    x"29CA2600",
    x"29CA0CBD",
    x"29C9F37D",
    x"29C9DA40",
    x"29C9C107",
    x"29C9A7D0",
    x"29C98E9D",
    x"29C9756D",
    x"29C95C3F",
    x"29C94315",
    x"29C929EF",
    x"29C910CB",
    x"29C8F7AA",
    x"29C8DE8D",
    x"29C8C573",
    x"29C8AC5C",
    x"29C89348",
    x"29C87A37",
    x"29C86129",
    x"29C8481F",
    x"29C82F17",
    x"29C81613",
    x"29C7FD12",
    x"29C7E414",
    x"29C7CB19",
    x"29C7B221",
    x"29C7992C",
    x"29C7803A",
    x"29C7674C",
    x"29C74E61",
    x"29C73578",
    x"29C71C93",
    x"29C703B1",
    x"29C6EAD2",
    x"29C6D1F7",
    x"29C6B91E",
    x"29C6A048",
    x"29C68776",
    x"29C66EA6",
    x"29C655DA",
    x"29C63D11",
    x"29C6244B",
    x"29C60B88",
    x"29C5F2C8",
    x"29C5DA0B",
    x"29C5C151",
    x"29C5A89B",
    x"29C58FE7",
    x"29C57737",
    x"29C55E8A",
    x"29C545DF",
    x"29C52D38",
    x"29C51494",
    x"29C4FBF3",
    x"29C4E355",
    x"29C4CABA",
    x"29C4B222",
    x"29C4998E",
    x"29C480FC",
    x"29C4686D",
    x"29C44FE2",
    x"29C43759",
    x"29C41ED4",
    x"29C40652",
    x"29C3EDD2",
    x"29C3D556",
    x"29C3BCDD",
    x"29C3A467",
    x"29C38BF4",
    x"29C37384",
    x"29C35B17",
    x"29C342AD",
    x"29C32A46",
    x"29C311E3",
    x"29C2F982",
    x"29C2E124",
    x"29C2C8CA",
    x"29C2B072",
    x"29C2981D",
    x"29C27FCC",
    x"29C2677E",
    x"29C24F32",
    x"29C236EA",
    x"29C21EA4",
    x"29C20662",
    x"29C1EE23",
    x"29C1D5E7",
    x"29C1BDAD",
    x"29C1A577",
    x"29C18D44",
    x"29C17514",
    x"29C15CE7",
    x"29C144BD",
    x"29C12C96",
    x"29C11471",
    x"29C0FC50",
    x"29C0E432",
    x"29C0CC17",
    x"29C0B3FF",
    x"29C09BEA",
    x"29C083D8",
    x"29C06BC9",
    x"29C053BD",
    x"29C03BB4",
    x"29C023AE",
    x"29C00BAC",
    x"29BFF3AC",
    x"29BFDBAF",
    x"29BFC3B5",
    x"29BFABBE",
    x"29BF93CA",
    x"29BF7BD9",
    x"29BF63EB",
    x"29BF4C00",
    x"29BF3418",
    x"29BF1C33",
    x"29BF0451",
    x"29BEEC72",
    x"29BED496",
    x"29BEBCBD",
    x"29BEA4E6",
    x"29BE8D13",
    x"29BE7543",
    x"29BE5D76",
    x"29BE45AC",
    x"29BE2DE5",
    x"29BE1620",
    x"29BDFE5F",
    x"29BDE6A1",
    x"29BDCEE5",
    x"29BDB72D",
    x"29BD9F78",
    x"29BD87C5",
    x"29BD7016",
    x"29BD5869",
    x"29BD40C0",
    x"29BD2919",
    x"29BD1175",
    x"29BCF9D5",
    x"29BCE237",
    x"29BCCA9C",
    x"29BCB304",
    x"29BC9B6F",
    x"29BC83DD",
    x"29BC6C4E",
    x"29BC54C2",
    x"29BC3D39",
    x"29BC25B3",
    x"29BC0E30",
    x"29BBF6AF",
    x"29BBDF32",
    x"29BBC7B8",
    x"29BBB040",
    x"29BB98CB",
    x"29BB815A",
    x"29BB69EB",
    x"29BB527F",
    x"29BB3B17",
    x"29BB23B1",
    x"29BB0C4E",
    x"29BAF4EE",
    x"29BADD90",
    x"29BAC636",
    x"29BAAEDF",
    x"29BA978A",
    x"29BA8039",
    x"29BA68EA",
    x"29BA519F",
    x"29BA3A56",
    x"29BA2310",
    x"29BA0BCD",
    x"29B9F48D",
    x"29B9DD50",
    x"29B9C616",
    x"29B9AEDF",
    x"29B997AA",
    x"29B98079",
    x"29B9694A",
    x"29B9521E",
    x"29B93AF5",
    x"29B923D0",
    x"29B90CAD",
    x"29B8F58C",
    x"29B8DE6F",
    x"29B8C755",
    x"29B8B03D",
    x"29B89929",
    x"29B88217",
    x"29B86B08",
    x"29B853FC",
    x"29B83CF3",
    x"29B825ED",
    x"29B80EEA",
    x"29B7F7E9",
    x"29B7E0EC",
    x"29B7C9F1",
    x"29B7B2F9",
    x"29B79C04",
    x"29B78512",
    x"29B76E23",
    x"29B75737",
    x"29B7404D",
    x"29B72967",
    x"29B71283",
    x"29B6FBA2",
    x"29B6E4C4",
    x"29B6CDE9",
    x"29B6B710",
    x"29B6A03B",
    x"29B68968",
    x"29B67299",
    x"29B65BCC",
    x"29B64502",
    x"29B62E3B",
    x"29B61776",
    x"29B600B5",
    x"29B5E9F6",
    x"29B5D33A",
    x"29B5BC81",
    x"29B5A5CB",
    x"29B58F18",
    x"29B57867",
    x"29B561BA",
    x"29B54B0F",
    x"29B53467",
    x"29B51DC2",
    x"29B5071F",
    x"29B4F080",
    x"29B4D9E3",
    x"29B4C349",
    x"29B4ACB2",
    x"29B4961E",
    x"29B47F8D",
    x"29B468FE",
    x"29B45273",
    x"29B43BEA",
    x"29B42564",
    x"29B40EE0",
    x"29B3F860",
    x"29B3E1E2",
    x"29B3CB68",
    x"29B3B4F0",
    x"29B39E7A",
    x"29B38808",
    x"29B37198",
    x"29B35B2B",
    x"29B344C2",
    x"29B32E5A",
    x"29B317F6",
    x"29B30194",
    x"29B2EB36",
    x"29B2D4DA",
    x"29B2BE80",
    x"29B2A82A",
    x"29B291D6",
    x"29B27B85",
    x"29B26537",
    x"29B24EEC",
    x"29B238A4",
    x"29B2225E",
    x"29B20C1B",
    x"29B1F5DB",
    x"29B1DF9E",
    x"29B1C963",
    x"29B1B32B",
    x"29B19CF6",
    x"29B186C4",
    x"29B17095",
    x"29B15A68",
    x"29B1443E",
    x"29B12E17",
    x"29B117F2",
    x"29B101D1",
    x"29B0EBB2",
    x"29B0D596",
    x"29B0BF7D",
    x"29B0A966",
    x"29B09352",
    x"29B07D41",
    x"29B06733",
    x"29B05127",
    x"29B03B1F",
    x"29B02519",
    x"29B00F15",
    x"29AFF915",
    x"29AFE317",
    x"29AFCD1C",
    x"29AFB724",
    x"29AFA12E",
    x"29AF8B3C",
    x"29AF754B",
    x"29AF5F5E",
    x"29AF4974",
    x"29AF338C",
    x"29AF1DA7",
    x"29AF07C4",
    x"29AEF1E5",
    x"29AEDC08",
    x"29AEC62E",
    x"29AEB056",
    x"29AE9A82",
    x"29AE84B0",
    x"29AE6EE1",
    x"29AE5914",
    x"29AE434A",
    x"29AE2D83",
    x"29AE17BF",
    x"29AE01FD",
    x"29ADEC3E",
    x"29ADD682",
    x"29ADC0C9",
    x"29ADAB12",
    x"29AD955E",
    x"29AD7FAD",
    x"29AD69FE",
    x"29AD5452",
    x"29AD3EA9",
    x"29AD2903",
    x"29AD135F",
    x"29ACFDBE",
    x"29ACE81F",
    x"29ACD284",
    x"29ACBCEB",
    x"29ACA754",
    x"29AC91C1",
    x"29AC7C30",
    x"29AC66A2",
    x"29AC5116",
    x"29AC3B8E",
    x"29AC2607",
    x"29AC1084",
    x"29ABFB03",
    x"29ABE585",
    x"29ABD00A",
    x"29ABBA91",
    x"29ABA51B",
    x"29AB8FA8",
    x"29AB7A37",
    x"29AB64C9",
    x"29AB4F5E",
    x"29AB39F6",
    x"29AB2490",
    x"29AB0F2C",
    x"29AAF9CC",
    x"29AAE46E",
    x"29AACF13",
    x"29AAB9BA",
    x"29AAA464",
    x"29AA8F11",
    x"29AA79C1",
    x"29AA6473",
    x"29AA4F27",
    x"29AA39DF",
    x"29AA2499",
    x"29AA0F56",
    x"29A9FA15",
    x"29A9E4D7",
    x"29A9CF9C",
    x"29A9BA63",
    x"29A9A52D",
    x"29A98FFA",
    x"29A97AC9",
    x"29A9659B",
    x"29A95070",
    x"29A93B47",
    x"29A92621",
    x"29A910FE",
    x"29A8FBDD",
    x"29A8E6BF",
    x"29A8D1A3",
    x"29A8BC8A",
    x"29A8A774",
    x"29A89260",
    x"29A87D4F",
    x"29A86841",
    x"29A85335",
    x"29A83E2C",
    x"29A82926",
    x"29A81422",
    x"29A7FF21",
    x"29A7EA22",
    x"29A7D526",
    x"29A7C02D",
    x"29A7AB36",
    x"29A79642",
    x"29A78151",
    x"29A76C62",
    x"29A75776",
    x"29A7428C",
    x"29A72DA5",
    x"29A718C1",
    x"29A703DF",
    x"29A6EF00",
    x"29A6DA23",
    x"29A6C549",
    x"29A6B072",
    x"29A69B9D",
    x"29A686CB",
    x"29A671FB",
    x"29A65D2E",
    x"29A64864",
    x"29A6339C",
    x"29A61ED7",
    x"29A60A14",
    x"29A5F555",
    x"29A5E097",
    x"29A5CBDC",
    x"29A5B724",
    x"29A5A26F",
    x"29A58DBC",
    x"29A5790B",
    x"29A5645D",
    x"29A54FB2",
    x"29A53B09",
    x"29A52663",
    x"29A511C0",
    x"29A4FD1F",
    x"29A4E881",
    x"29A4D3E5",
    x"29A4BF4C",
    x"29A4AAB5",
    x"29A49621",
    x"29A4818F",
    x"29A46D00",
    x"29A45874",
    x"29A443EA",
    x"29A42F63",
    x"29A41ADF",
    x"29A4065C",
    x"29A3F1DD",
    x"29A3DD60",
    x"29A3C8E6",
    x"29A3B46E",
    x"29A39FF8",
    x"29A38B86",
    x"29A37716",
    x"29A362A8",
    x"29A34E3D",
    x"29A339D4",
    x"29A3256E",
    x"29A3110B",
    x"29A2FCAA",
    x"29A2E84C",
    x"29A2D3F0",
    x"29A2BF97",
    x"29A2AB40",
    x"29A296EC",
    x"29A2829A",
    x"29A26E4B",
    x"29A259FF",
    x"29A245B5",
    x"29A2316D",
    x"29A21D29",
    x"29A208E6",
    x"29A1F4A6",
    x"29A1E069",
    x"29A1CC2E",
    x"29A1B7F6",
    x"29A1A3C0",
    x"29A18F8D",
    x"29A17B5C",
    x"29A1672E",
    x"29A15303",
    x"29A13ED9",
    x"29A12AB3",
    x"29A1168F",
    x"29A1026D",
    x"29A0EE4E",
    x"29A0DA32",
    x"29A0C618",
    x"29A0B200",
    x"29A09DEB",
    x"29A089D9",
    x"29A075C9",
    x"29A061BB",
    x"29A04DB0",
    x"29A039A8",
    x"29A025A2",
    x"29A0119E",
    x"299FFD9D",
    x"299FE99F",
    x"299FD5A3",
    x"299FC1AA",
    x"299FADB3",
    x"299F99BE",
    x"299F85CC",
    x"299F71DD",
    x"299F5DF0",
    x"299F4A05",
    x"299F361D",
    x"299F2238",
    x"299F0E55",
    x"299EFA74",
    x"299EE696",
    x"299ED2BA",
    x"299EBEE1",
    x"299EAB0B",
    x"299E9737",
    x"299E8365",
    x"299E6F96",
    x"299E5BC9",
    x"299E47FF",
    x"299E3437",
    x"299E2072",
    x"299E0CAF",
    x"299DF8EF",
    x"299DE531",
    x"299DD175",
    x"299DBDBC",
    x"299DAA06",
    x"299D9652",
    x"299D82A0",
    x"299D6EF1",
    x"299D5B45",
    x"299D479A",
    x"299D33F3",
    x"299D204D",
    x"299D0CAB",
    x"299CF90A",
    x"299CE56C",
    x"299CD1D1",
    x"299CBE38",
    x"299CAAA1",
    x"299C970D",
    x"299C837B",
    x"299C6FEC",
    x"299C5C60",
    x"299C48D5",
    x"299C354D",
    x"299C21C8",
    x"299C0E45",
    x"299BFAC4",
    x"299BE746",
    x"299BD3CA",
    x"299BC051",
    x"299BACDA",
    x"299B9966",
    x"299B85F4",
    x"299B7285",
    x"299B5F17",
    x"299B4BAD",
    x"299B3844",
    x"299B24DF",
    x"299B117B",
    x"299AFE1A",
    x"299AEABC",
    x"299AD760",
    x"299AC406",
    x"299AB0AF",
    x"299A9D5A",
    x"299A8A07",
    x"299A76B7",
    x"299A636A",
    x"299A501E",
    x"299A3CD6",
    x"299A298F",
    x"299A164B",
    x"299A030A",
    x"2999EFCA",
    x"2999DC8E",
    x"2999C953",
    x"2999B61B",
    x"2999A2E6",
    x"29998FB3",
    x"29997C82",
    x"29996953",
    x"29995627",
    x"299942FE",
    x"29992FD7",
    x"29991CB2",
    x"29990990",
    x"2998F670",
    x"2998E352",
    x"2998D037",
    x"2998BD1E",
    x"2998AA07",
    x"299896F3",
    x"299883E2",
    x"299870D2",
    x"29985DC6",
    x"29984ABB",
    x"299837B3",
    x"299824AD",
    x"299811AA",
    x"2997FEA9",
    x"2997EBAA",
    x"2997D8AE",
    x"2997C5B4",
    x"2997B2BC",
    x"29979FC7",
    x"29978CD4",
    x"299779E4",
    x"299766F6",
    x"2997540A",
    x"29974121",
    x"29972E3A",
    x"29971B55",
    x"29970873",
    x"2996F593",
    x"2996E2B6",
    x"2996CFDB",
    x"2996BD02",
    x"2996AA2B",
    x"29969757",
    x"29968485",
    x"299671B6",
    x"29965EE9",
    x"29964C1E",
    x"29963956",
    x"29962690",
    x"299613CC",
    x"2996010B",
    x"2995EE4C",
    x"2995DB8F",
    x"2995C8D5",
    x"2995B61D",
    x"2995A368",
    x"299590B4",
    x"29957E03",
    x"29956B55",
    x"299558A9",
    x"299545FF",
    x"29953357",
    x"299520B2",
    x"29950E0F",
    x"2994FB6E",
    x"2994E8D0",
    x"2994D634",
    x"2994C39B",
    x"2994B103",
    x"29949E6E",
    x"29948BDC",
    x"2994794B",
    x"299466BD",
    x"29945432",
    x"299441A8",
    x"29942F21",
    x"29941C9D",
    x"29940A1A",
    x"2993F79A",
    x"2993E51C",
    x"2993D2A1",
    x"2993C028",
    x"2993ADB1",
    x"29939B3C",
    x"299388CA",
    x"2993765A",
    x"299363EC",
    x"29935181",
    x"29933F18",
    x"29932CB1",
    x"29931A4D",
    x"299307EB",
    x"2992F58B",
    x"2992E32D",
    x"2992D0D2",
    x"2992BE79",
    x"2992AC22",
    x"299299CE",
    x"2992877C",
    x"2992752C",
    x"299262DF",
    x"29925093",
    x"29923E4A",
    x"29922C04",
    x"299219BF",
    x"2992077D",
    x"2991F53E",
    x"2991E300",
    x"2991D0C5",
    x"2991BE8C",
    x"2991AC55",
    x"29919A21",
    x"299187EF",
    x"299175BF",
    x"29916391",
    x"29915166",
    x"29913F3D",
    x"29912D16",
    x"29911AF2",
    x"299108CF",
    x"2990F6AF",
    x"2990E492",
    x"2990D276",
    x"2990C05D",
    x"2990AE46",
    x"29909C32",
    x"29908A1F",
    x"2990780F",
    x"29906601",
    x"299053F5",
    x"299041EC",
    x"29902FE5",
    x"29901DE0",
    x"29900BDE",
    x"298FF9DD",
    x"298FE7DF",
    x"298FD5E3",
    x"298FC3EA",
    x"298FB1F2",
    x"298F9FFD",
    x"298F8E0A",
    x"298F7C1A",
    x"298F6A2B",
    x"298F583F",
    x"298F4655",
    x"298F346D",
    x"298F2288",
    x"298F10A5",
    x"298EFEC4",
    x"298EECE5",
    x"298EDB09",
    x"298EC92E",
    x"298EB756",
    x"298EA581",
    x"298E93AD",
    x"298E81DC",
    x"298E700C",
    x"298E5E40",
    x"298E4C75",
    x"298E3AAC",
    x"298E28E6",
    x"298E1722",
    x"298E0560",
    x"298DF3A1",
    x"298DE1E4",
    x"298DD028",
    x"298DBE70",
    x"298DACB9",
    x"298D9B04",
    x"298D8952",
    x"298D77A2",
    x"298D65F4",
    x"298D5449",
    x"298D429F",
    x"298D30F8",
    x"298D1F53",
    x"298D0DB0",
    x"298CFC0F",
    x"298CEA71",
    x"298CD8D5",
    x"298CC73B",
    x"298CB5A3",
    x"298CA40D",
    x"298C927A",
    x"298C80E9",
    x"298C6F5A",
    x"298C5DCD",
    x"298C4C42",
    x"298C3ABA",
    x"298C2934",
    x"298C17B0",
    x"298C062E",
    x"298BF4AE",
    x"298BE331",
    x"298BD1B5",
    x"298BC03C",
    x"298BAEC5",
    x"298B9D50",
    x"298B8BDE",
    x"298B7A6D",
    x"298B68FF",
    x"298B5793",
    x"298B4629",
    x"298B34C2",
    x"298B235C",
    x"298B11F9",
    x"298B0098",
    x"298AEF39",
    x"298ADDDC",
    x"298ACC81",
    x"298ABB29",
    x"298AA9D2",
    x"298A987E",
    x"298A872C",
    x"298A75DC",
    x"298A648F",
    x"298A5343",
    x"298A41FA",
    x"298A30B3",
    x"298A1F6E",
    x"298A0E2B",
    x"2989FCEA",
    x"2989EBAC",
    x"2989DA6F",
    x"2989C935",
    x"2989B7FD",
    x"2989A6C7",
    x"29899593",
    x"29898462",
    x"29897332",
    x"29896205",
    x"298950DA",
    x"29893FB1",
    x"29892E8A",
    x"29891D65",
    x"29890C43",
    x"2988FB22",
    x"2988EA04",
    x"2988D8E8",
    x"2988C7CE",
    x"2988B6B6",
    x"2988A5A0",
    x"2988948C",
    x"2988837B",
    x"2988726B",
    x"2988615E",
    x"29885053",
    x"29883F4A",
    x"29882E43",
    x"29881D3E",
    x"29880C3C",
    x"2987FB3B",
    x"2987EA3D",
    x"2987D941",
    x"2987C847",
    x"2987B74F",
    x"2987A659",
    x"29879565",
    x"29878474",
    x"29877384",
    x"29876297",
    x"298751AB",
    x"298740C2",
    x"29872FDB",
    x"29871EF6",
    x"29870E13",
    x"2986FD33",
    x"2986EC54",
    x"2986DB78",
    x"2986CA9D",
    x"2986B9C5",
    x"2986A8EF",
    x"2986981B",
    x"29868749",
    x"29867679",
    x"298665AB",
    x"298654E0",
    x"29864416",
    x"2986334F",
    x"29862289",
    x"298611C6",
    x"29860105",
    x"2985F046",
    x"2985DF89",
    x"2985CECE",
    x"2985BE15",
    x"2985AD5E",
    x"29859CAA",
    x"29858BF7",
    x"29857B47",
    x"29856A98",
    x"298559EC",
    x"29854942",
    x"2985389A",
    x"298527F4",
    x"29851750",
    x"298506AE",
    x"2984F60E",
    x"2984E570",
    x"2984D4D5",
    x"2984C43B",
    x"2984B3A4",
    x"2984A30E",
    x"2984927B",
    x"298481EA",
    x"2984715A",
    x"298460CD",
    x"29845042",
    x"29843FB9",
    x"29842F32",
    x"29841EAD",
    x"29840E2B",
    x"2983FDAA",
    x"2983ED2B",
    x"2983DCAF",
    x"2983CC34",
    x"2983BBBB",
    x"2983AB45",
    x"29839AD1",
    x"29838A5E",
    x"298379EE",
    x"29836980",
    x"29835914",
    x"298348AA",
    x"29833842",
    x"298327DC",
    x"29831778",
    x"29830716",
    x"2982F6B6",
    x"2982E658",
    x"2982D5FC",
    x"2982C5A2",
    x"2982B54B",
    x"2982A4F5",
    x"298294A2",
    x"29828450",
    x"29827400",
    x"298263B3",
    x"29825368",
    x"2982431E",
    x"298232D7",
    x"29822291",
    x"2982124E",
    x"2982020D",
    x"2981F1CE",
    x"2981E190",
    x"2981D155",
    x"2981C11C",
    x"2981B0E5",
    x"2981A0B0",
    x"2981907D",
    x"2981804C",
    x"2981701D",
    x"29815FF0",
    x"29814FC5",
    x"29813F9C",
    x"29812F75",
    x"29811F50",
    x"29810F2D",
    x"2980FF0C",
    x"2980EEED",
    x"2980DED0",
    x"2980CEB6",
    x"2980BE9D",
    x"2980AE86",
    x"29809E71",
    x"29808E5E",
    x"29807E4D",
    x"29806E3F",
    x"29805E32",
    x"29804E27",
    x"29803E1E",
    x"29802E18",
    x"29801E13",
    x"29800E10",
    x"297FFC1F",
    x"297FDC21",
    x"297FBC28",
    x"297F9C32",
    x"297F7C41",
    x"297F5C53",
    x"297F3C69",
    x"297F1C84",
    x"297EFCA2",
    x"297EDCC5",
    x"297EBCEB",
    x"297E9D16",
    x"297E7D44",
    x"297E5D76",
    x"297E3DAC",
    x"297E1DE7",
    x"297DFE25",
    x"297DDE67",
    x"297DBEAD",
    x"297D9EF8",
    x"297D7F46",
    x"297D5F98",
    x"297D3FEE",
    x"297D2048",
    x"297D00A6",
    x"297CE108",
    x"297CC16D",
    x"297CA1D7",
    x"297C8245",
    x"297C62B7",
    x"297C432C",
    x"297C23A6",
    x"297C0423",
    x"297BE4A5",
    x"297BC52A",
    x"297BA5B4",
    x"297B8641",
    x"297B66D2",
    x"297B4767",
    x"297B2800",
    x"297B089D",
    x"297AE93E",
    x"297AC9E3",
    x"297AAA8C",
    x"297A8B38",
    x"297A6BE9",
    x"297A4C9D",
    x"297A2D56",
    x"297A0E12",
    x"2979EED2",
    x"2979CF96",
    x"2979B05E",
    x"2979912A",
    x"297971FA",
    x"297952CE",
    x"297933A5",
    x"29791481",
    x"2978F560",
    x"2978D643",
    x"2978B72A",
    x"29789816",
    x"29787904",
    x"297859F7",
    x"29783AEE",
    x"29781BE9",
    x"2977FCE7",
    x"2977DDE9",
    x"2977BEEF",
    x"29779FFA",
    x"29778107",
    x"29776219",
    x"2977432F",
    x"29772449",
    x"29770566",
    x"2976E687",
    x"2976C7AC",
    x"2976A8D5",
    x"29768A02",
    x"29766B33",
    x"29764C67",
    x"29762DA0",
    x"29760EDC",
    x"2975F01C",
    x"2975D160",
    x"2975B2A8",
    x"297593F3",
    x"29757543",
    x"29755696",
    x"297537ED",
    x"29751948",
    x"2974FAA7",
    x"2974DC09",
    x"2974BD70",
    x"29749EDA",
    x"29748048",
    x"297461BA",
    x"2974432F",
    x"297424A9",
    x"29740626",
    x"2973E7A7",
    x"2973C92C",
    x"2973AAB5",
    x"29738C42",
    x"29736DD2",
    x"29734F66",
    x"297330FE",
    x"2973129A",
    x"2972F43A",
    x"2972D5DD",
    x"2972B784",
    x"2972992F",
    x"29727ADE",
    x"29725C90",
    x"29723E47",
    x"29722001",
    x"297201BF",
    x"2971E380",
    x"2971C546",
    x"2971A70F",
    x"297188DC",
    x"29716AAD",
    x"29714C81",
    x"29712E5A",
    x"29711036",
    x"2970F216",
    x"2970D3F9",
    x"2970B5E1",
    x"297097CC",
    x"297079BB",
    x"29705BAD",
    x"29703DA4",
    x"29701F9E",
    x"2970019C",
    x"296FE39E",
    x"296FC5A3",
    x"296FA7AC",
    x"296F89B9",
    x"296F6BCA",
    x"296F4DDE",
    x"296F2FF6",
    x"296F1212",
    x"296EF432",
    x"296ED655",
    x"296EB87C",
    x"296E9AA7",
    x"296E7CD5",
    x"296E5F08",
    x"296E413E",
    x"296E2377",
    x"296E05B5",
    x"296DE7F6",
    x"296DCA3B",
    x"296DAC83",
    x"296D8ED0",
    x"296D7120",
    x"296D5373",
    x"296D35CB",
    x"296D1826",
    x"296CFA85",
    x"296CDCE7",
    x"296CBF4E",
    x"296CA1B8",
    x"296C8425",
    x"296C6696",
    x"296C490C",
    x"296C2B84",
    x"296C0E01",
    x"296BF081",
    x"296BD305",
    x"296BB58C",
    x"296B9817",
    x"296B7AA6",
    x"296B5D38",
    x"296B3FCF",
    x"296B2268",
    x"296B0506",
    x"296AE7A7",
    x"296ACA4C",
    x"296AACF5",
    x"296A8FA1",
    x"296A7251",
    x"296A5504",
    x"296A37BC",
    x"296A1A76",
    x"2969FD35",
    x"2969DFF7",
    x"2969C2BD",
    x"2969A586",
    x"29698854",
    x"29696B24",
    x"29694DF9",
    x"296930D1",
    x"296913AD",
    x"2968F68C",
    x"2968D96F",
    x"2968BC56",
    x"29689F40",
    x"2968822E",
    x"2968651F",
    x"29684814",
    x"29682B0D",
    x"29680E0A",
    x"2967F10A",
    x"2967D40D",
    x"2967B715",
    x"29679A20",
    x"29677D2E",
    x"29676040",
    x"29674356",
    x"29672670",
    x"2967098D",
    x"2966ECAD",
    x"2966CFD1",
    x"2966B2F9",
    x"29669625",
    x"29667954",
    x"29665C86",
    x"29663FBC",
    x"296622F6",
    x"29660634",
    x"2965E975",
    x"2965CCB9",
    x"2965B002",
    x"2965934D",
    x"2965769D",
    x"296559F0",
    x"29653D46",
    x"296520A0",
    x"296503FE",
    x"2964E75F",
    x"2964CAC4",
    x"2964AE2D",
    x"29649199",
    x"29647508",
    x"2964587B",
    x"29643BF2",
    x"29641F6C",
    x"296402EA",
    x"2963E66C",
    x"2963C9F1",
    x"2963AD79",
    x"29639105",
    x"29637495",
    x"29635828",
    x"29633BBF",
    x"29631F59",
    x"296302F7",
    x"2962E699",
    x"2962CA3D",
    x"2962ADE6",
    x"29629192",
    x"29627542",
    x"296258F5",
    x"29623CAB",
    x"29622066",
    x"29620423",
    x"2961E7E5",
    x"2961CBA9",
    x"2961AF72",
    x"2961933D",
    x"2961770D",
    x"29615AE0",
    x"29613EB6",
    x"29612290",
    x"2961066D",
    x"2960EA4E",
    x"2960CE33",
    x"2960B21B",
    x"29609606",
    x"296079F5",
    x"29605DE8",
    x"296041DE",
    x"296025D7",
    x"296009D4",
    x"295FEDD5",
    x"295FD1D9",
    x"295FB5E0",
    x"295F99EB",
    x"295F7DFA",
    x"295F620C",
    x"295F4621",
    x"295F2A3A",
    x"295F0E57",
    x"295EF277",
    x"295ED69A",
    x"295EBAC1",
    x"295E9EEC",
    x"295E8319",
    x"295E674B",
    x"295E4B80",
    x"295E2FB8",
    x"295E13F4",
    x"295DF833",
    x"295DDC76",
    x"295DC0BC",
    x"295DA505",
    x"295D8953",
    x"295D6DA3",
    x"295D51F7",
    x"295D364F",
    x"295D1AAA",
    x"295CFF08",
    x"295CE36A",
    x"295CC7CF",
    x"295CAC38",
    x"295C90A4",
    x"295C7514",
    x"295C5987",
    x"295C3DFD",
    x"295C2277",
    x"295C06F5",
    x"295BEB76",
    x"295BCFFA",
    x"295BB482",
    x"295B990D",
    x"295B7D9B",
    x"295B622D",
    x"295B46C3",
    x"295B2B5C",
    x"295B0FF8",
    x"295AF498",
    x"295AD93B",
    x"295ABDE1",
    x"295AA28B",
    x"295A8739",
    x"295A6BE9",
    x"295A509E",
    x"295A3555",
    x"295A1A10",
    x"2959FECF",
    x"2959E391",
    x"2959C856",
    x"2959AD1F",
    x"295991EB",
    x"295976BA",
    x"29595B8D",
    x"29594063",
    x"2959253D",
    x"29590A1A",
    x"2958EEFA",
    x"2958D3DE",
    x"2958B8C5",
    x"29589DB0",
    x"2958829E",
    x"2958678F",
    x"29584C84",
    x"2958317C",
    x"29581678",
    x"2957FB77",
    x"2957E079",
    x"2957C57E",
    x"2957AA87",
    x"29578F94",
    x"295774A4",
    x"295759B7",
    x"29573ECD",
    x"295723E7",
    x"29570904",
    x"2956EE25",
    x"2956D349",
    x"2956B870",
    x"29569D9B",
    x"295682C8",
    x"295667FA",
    x"29564D2E",
    x"29563267",
    x"295617A2",
    x"2955FCE1",
    x"2955E223",
    x"2955C768",
    x"2955ACB1",
    x"295591FD",
    x"2955774C",
    x"29555C9F",
    x"295541F5",
    x"2955274F",
    x"29550CAB",
    x"2954F20B",
    x"2954D76F",
    x"2954BCD6",
    x"2954A240",
    x"295487AD",
    x"29546D1E",
    x"29545292",
    x"29543809",
    x"29541D84",
    x"29540302",
    x"2953E883",
    x"2953CE08",
    x"2953B38F",
    x"2953991B",
    x"29537EA9",
    x"2953643B",
    x"295349D0",
    x"29532F69",
    x"29531504",
    x"2952FAA3",
    x"2952E046",
    x"2952C5EB",
    x"2952AB94",
    x"29529140",
    x"295276F0",
    x"29525CA3",
    x"29524259",
    x"29522812",
    x"29520DCF",
    x"2951F38F",
    x"2951D952",
    x"2951BF18",
    x"2951A4E2",
    x"29518AAF",
    x"2951707F",
    x"29515653",
    x"29513C2A",
    x"29512204",
    x"295107E1",
    x"2950EDC2",
    x"2950D3A6",
    x"2950B98D",
    x"29509F77",
    x"29508565",
    x"29506B56",
    x"2950514A",
    x"29503742",
    x"29501D3C",
    x"2950033A",
    x"294FE93C",
    x"294FCF40",
    x"294FB548",
    x"294F9B53",
    x"294F8161",
    x"294F6772",
    x"294F4D87",
    x"294F339F",
    x"294F19BA",
    x"294EFFD9",
    x"294EE5FA",
    x"294ECC1F",
    x"294EB247",
    x"294E9873",
    x"294E7EA1",
    x"294E64D3",
    x"294E4B08",
    x"294E3140",
    x"294E177C",
    x"294DFDBA",
    x"294DE3FC",
    x"294DCA41",
    x"294DB08A",
    x"294D96D5",
    x"294D7D24",
    x"294D6376",
    x"294D49CB",
    x"294D3023",
    x"294D167F",
    x"294CFCDE",
    x"294CE340",
    x"294CC9A5",
    x"294CB00D",
    x"294C9679",
    x"294C7CE8",
    x"294C635A",
    x"294C49CF",
    x"294C3047",
    x"294C16C3",
    x"294BFD42",
    x"294BE3C3",
    x"294BCA49",
    x"294BB0D1",
    x"294B975C",
    x"294B7DEB",
    x"294B647D",
    x"294B4B12",
    x"294B31AA",
    x"294B1846",
    x"294AFEE4",
    x"294AE586",
    x"294ACC2B",
    x"294AB2D3",
    x"294A997E",
    x"294A802C",
    x"294A66DE",
    x"294A4D93",
    x"294A344B",
    x"294A1B06",
    x"294A01C4",
    x"2949E885",
    x"2949CF4A",
    x"2949B611",
    x"29499CDC",
    x"294983AA",
    x"29496A7B",
    x"29495150",
    x"29493827",
    x"29491F01",
    x"294905DF",
    x"2948ECC0",
    x"2948D3A4",
    x"2948BA8B",
    x"2948A175",
    x"29488863",
    x"29486F53",
    x"29485647",
    x"29483D3E",
    x"29482438",
    x"29480B35",
    x"2947F235",
    x"2947D938",
    x"2947C03E",
    x"2947A748",
    x"29478E55",
    x"29477564",
    x"29475C77",
    x"2947438D",
    x"29472AA6",
    x"294711C3",
    x"2946F8E2",
    x"2946E004",
    x"2946C72A",
    x"2946AE53",
    x"2946957E",
    x"29467CAD",
    x"294663DF",
    x"29464B14",
    x"2946324C",
    x"29461988",
    x"294600C6",
    x"2945E808",
    x"2945CF4C",
    x"2945B694",
    x"29459DDE",
    x"2945852C",
    x"29456C7D",
    x"294553D1",
    x"29453B28",
    x"29452282",
    x"294509E0",
    x"2944F140",
    x"2944D8A3",
    x"2944C00A",
    x"2944A773",
    x"29448EE0",
    x"29447650",
    x"29445DC2",
    x"29444538",
    x"29442CB1",
    x"2944142D",
    x"2943FBAC",
    x"2943E32E",
    x"2943CAB3",
    x"2943B23B",
    x"294399C7",
    x"29438155",
    x"294368E6",
    x"2943507B",
    x"29433812",
    x"29431FAD",
    x"2943074A",
    x"2942EEEB",
    x"2942D68E",
    x"2942BE35",
    x"2942A5DF",
    x"29428D8C",
    x"2942753C",
    x"29425CEE",
    x"294244A4",
    x"29422C5D",
    x"29421419",
    x"2941FBD8",
    x"2941E39A",
    x"2941CB5F",
    x"2941B327",
    x"29419AF2",
    x"294182C1",
    x"29416A92",
    x"29415266",
    x"29413A3D",
    x"29412217",
    x"294109F5",
    x"2940F1D5",
    x"2940D9B8",
    x"2940C19F",
    x"2940A988",
    x"29409174",
    x"29407963",
    x"29406156",
    x"2940494B",
    x"29403143",
    x"2940193F",
    x"2940013D",
    x"293FE93E",
    x"293FD143",
    x"293FB94A",
    x"293FA155",
    x"293F8962",
    x"293F7172",
    x"293F5985",
    x"293F419C",
    x"293F29B5",
    x"293F11D1",
    x"293EF9F1",
    x"293EE213",
    x"293ECA38",
    x"293EB260",
    x"293E9A8C",
    x"293E82BA",
    x"293E6AEB",
    x"293E531F",
    x"293E3B56",
    x"293E2390",
    x"293E0BCD",
    x"293DF40D",
    x"293DDC50",
    x"293DC496",
    x"293DACDF",
    x"293D952B",
    x"293D7D7A",
    x"293D65CC",
    x"293D4E20",
    x"293D3678",
    x"293D1ED3",
    x"293D0730",
    x"293CEF91",
    x"293CD7F4",
    x"293CC05B",
    x"293CA8C4",
    x"293C9131",
    x"293C79A0",
    x"293C6212",
    x"293C4A87",
    x"293C3300",
    x"293C1B7B",
    x"293C03F9",
    x"293BEC7A",
    x"293BD4FE",
    x"293BBD84",
    x"293BA60E",
    x"293B8E9B",
    x"293B772B",
    x"293B5FBD",
    x"293B4853",
    x"293B30EB",
    x"293B1986",
    x"293B0225",
    x"293AEAC6",
    x"293AD36A",
    x"293ABC11",
    x"293AA4BB",
    x"293A8D68",
    x"293A7618",
    x"293A5ECA",
    x"293A4780",
    x"293A3038",
    x"293A18F4",
    x"293A01B2",
    x"2939EA73",
    x"2939D338",
    x"2939BBFF",
    x"2939A4C9",
    x"29398D95",
    x"29397665",
    x"29395F38",
    x"2939480D",
    x"293930E6",
    x"293919C1",
    x"2939029F",
    x"2938EB81",
    x"2938D465",
    x"2938BD4B",
    x"2938A635",
    x"29388F22",
    x"29387811",
    x"29386104",
    x"293849F9",
    x"293832F1",
    x"29381BEC",
    x"293804EA",
    x"2937EDEB",
    x"2937D6EF",
    x"2937BFF5",
    x"2937A8FF",
    x"2937920B",
    x"29377B1A",
    x"2937642C",
    x"29374D41",
    x"29373659",
    x"29371F74",
    x"29370891",
    x"2936F1B2",
    x"2936DAD5",
    x"2936C3FB",
    x"2936AD24",
    x"29369650",
    x"29367F7E",
    x"293668B0",
    x"293651E4",
    x"29363B1B",
    x"29362455",
    x"29360D92",
    x"2935F6D2",
    x"2935E015",
    x"2935C95A",
    x"2935B2A2",
    x"29359BED",
    x"2935853B",
    x"29356E8C",
    x"293557E0",
    x"29354136",
    x"29352A8F",
    x"293513EB",
    x"2934FD4A",
    x"2934E6AC",
    x"2934D011",
    x"2934B978",
    x"2934A2E2",
    x"29348C4F",
    x"293475BF",
    x"29345F32",
    x"293448A7",
    x"29343220",
    x"29341B9B",
    x"29340519",
    x"2933EE9A",
    x"2933D81D",
    x"2933C1A4",
    x"2933AB2D",
    x"293394B9",
    x"29337E48",
    x"293367D9",
    x"2933516E",
    x"29333B05",
    x"2933249F",
    x"29330E3C",
    x"2932F7DB",
    x"2932E17E",
    x"2932CB23",
    x"2932B4CB",
    x"29329E76",
    x"29328823",
    x"293271D4",
    x"29325B87",
    x"2932453D",
    x"29322EF6",
    x"293218B1",
    x"2932026F",
    x"2931EC30",
    x"2931D5F4",
    x"2931BFBB",
    x"2931A984",
    x"29319351",
    x"29317D20",
    x"293166F1",
    x"293150C6",
    x"29313A9D",
    x"29312477",
    x"29310E54",
    x"2930F834",
    x"2930E216",
    x"2930CBFB",
    x"2930B5E3",
    x"29309FCE",
    x"293089BB",
    x"293073AB",
    x"29305D9E",
    x"29304794",
    x"2930318C",
    x"29301B87",
    x"29300585",
    x"292FEF86",
    x"292FD989",
    x"292FC390",
    x"292FAD98",
    x"292F97A4",
    x"292F81B3",
    x"292F6BC4",
    x"292F55D8",
    x"292F3FEE",
    x"292F2A08",
    x"292F1424",
    x"292EFE43",
    x"292EE864",
    x"292ED289",
    x"292EBCB0",
    x"292EA6D9",
    x"292E9106",
    x"292E7B35",
    x"292E6567",
    x"292E4F9C",
    x"292E39D3",
    x"292E240D",
    x"292E0E4A",
    x"292DF88A",
    x"292DE2CC",
    x"292DCD11",
    x"292DB759",
    x"292DA1A3",
    x"292D8BF0",
    x"292D7640",
    x"292D6093",
    x"292D4AE8",
    x"292D3540",
    x"292D1F9B",
    x"292D09F8",
    x"292CF458",
    x"292CDEBB",
    x"292CC921",
    x"292CB389",
    x"292C9DF4",
    x"292C8861",
    x"292C72D2",
    x"292C5D45",
    x"292C47BA",
    x"292C3233",
    x"292C1CAE",
    x"292C072B",
    x"292BF1AC",
    x"292BDC2F",
    x"292BC6B5",
    x"292BB13D",
    x"292B9BC9",
    x"292B8656",
    x"292B70E7",
    x"292B5B7A",
    x"292B4610",
    x"292B30A9",
    x"292B1B44",
    x"292B05E2",
    x"292AF082",
    x"292ADB26",
    x"292AC5CC",
    x"292AB074",
    x"292A9B20",
    x"292A85CE",
    x"292A707E",
    x"292A5B31",
    x"292A45E7",
    x"292A30A0",
    x"292A1B5B",
    x"292A0619",
    x"2929F0DA",
    x"2929DB9D",
    x"2929C663",
    x"2929B12B",
    x"29299BF6",
    x"292986C4",
    x"29297195",
    x"29295C68",
    x"2929473E",
    x"29293216",
    x"29291CF1",
    x"292907CF",
    x"2928F2AF",
    x"2928DD92",
    x"2928C878",
    x"2928B360",
    x"29289E4B",
    x"29288938",
    x"29287429",
    x"29285F1B",
    x"29284A11",
    x"29283509",
    x"29282004",
    x"29280B01",
    x"2927F601",
    x"2927E103",
    x"2927CC09",
    x"2927B710",
    x"2927A21B",
    x"29278D28",
    x"29277838",
    x"2927634A",
    x"29274E5F",
    x"29273976",
    x"29272490",
    x"29270FAD",
    x"2926FACC",
    x"2926E5EE",
    x"2926D113",
    x"2926BC3A",
    x"2926A764",
    x"29269290",
    x"29267DBF",
    x"292668F1",
    x"29265425",
    x"29263F5C",
    x"29262A95",
    x"292615D1",
    x"29260110",
    x"2925EC51",
    x"2925D795",
    x"2925C2DB",
    x"2925AE24",
    x"2925996F",
    x"292584BE",
    x"2925700E",
    x"29255B62",
    x"292546B7",
    x"29253210",
    x"29251D6B",
    x"292508C9",
    x"2924F429",
    x"2924DF8B",
    x"2924CAF1",
    x"2924B659",
    x"2924A1C3",
    x"29248D30",
    x"292478A0",
    x"29246412",
    x"29244F87",
    x"29243AFE",
    x"29242678",
    x"292411F5",
    x"2923FD74",
    x"2923E8F5",
    x"2923D479",
    x"2923C000",
    x"2923AB89",
    x"29239715",
    x"292382A4",
    x"29236E35",
    x"292359C8",
    x"2923455E",
    x"292330F7",
    x"29231C92",
    x"29230830",
    x"2922F3D0",
    x"2922DF73",
    x"2922CB18",
    x"2922B6C0",
    x"2922A26A",
    x"29228E17",
    x"292279C7",
    x"29226579",
    x"2922512D",
    x"29223CE5",
    x"2922289E",
    x"2922145A",
    x"29220019",
    x"2921EBDA",
    x"2921D79E",
    x"2921C364",
    x"2921AF2D",
    x"29219AF9",
    x"292186C7",
    x"29217297",
    x"29215E6A",
    x"29214A3F",
    x"29213617",
    x"292121F2",
    x"29210DCF",
    x"2920F9AE",
    x"2920E590",
    x"2920D175",
    x"2920BD5C",
    x"2920A946",
    x"29209532",
    x"29208120",
    x"29206D11",
    x"29205905",
    x"292044FB",
    x"292030F4",
    x"29201CEF",
    x"292008ED",
    x"291FF4ED",
    x"291FE0EF",
    x"291FCCF5",
    x"291FB8FC",
    x"291FA506",
    x"291F9113",
    x"291F7D22",
    x"291F6934",
    x"291F5548",
    x"291F415E",
    x"291F2D77",
    x"291F1993",
    x"291F05B1",
    x"291EF1D2",
    x"291EDDF5",
    x"291ECA1A",
    x"291EB642",
    x"291EA26C",
    x"291E8E99",
    x"291E7AC9",
    x"291E66FB",
    x"291E532F",
    x"291E3F66",
    x"291E2B9F",
    x"291E17DB",
    x"291E0419",
    x"291DF05A",
    x"291DDC9D",
    x"291DC8E3",
    x"291DB52B",
    x"291DA176",
    x"291D8DC3",
    x"291D7A12",
    x"291D6664",
    x"291D52B8",
    x"291D3F0F",
    x"291D2B69",
    x"291D17C5",
    x"291D0423",
    x"291CF083",
    x"291CDCE7",
    x"291CC94C",
    x"291CB5B4",
    x"291CA21F",
    x"291C8E8C",
    x"291C7AFB",
    x"291C676D",
    x"291C53E1",
    x"291C4058",
    x"291C2CD1",
    x"291C194D",
    x"291C05CB",
    x"291BF24B",
    x"291BDECE",
    x"291BCB54",
    x"291BB7DC",
    x"291BA466",
    x"291B90F2",
    x"291B7D82",
    x"291B6A13",
    x"291B56A7",
    x"291B433D",
    x"291B2FD6",
    x"291B1C71",
    x"291B090F",
    x"291AF5AF",
    x"291AE252",
    x"291ACEF7",
    x"291ABB9E",
    x"291AA848",
    x"291A94F4",
    x"291A81A2",
    x"291A6E53",
    x"291A5B07",
    x"291A47BD",
    x"291A3475",
    x"291A2130",
    x"291A0DED",
    x"2919FAAC",
    x"2919E76E",
    x"2919D432",
    x"2919C0F9",
    x"2919ADC2",
    x"29199A8D",
    x"2919875B",
    x"2919742C",
    x"291960FE",
    x"29194DD3",
    x"29193AAB",
    x"29192785",
    x"29191461",
    x"29190140",
    x"2918EE21",
    x"2918DB04",
    x"2918C7EA",
    x"2918B4D2",
    x"2918A1BD",
    x"29188EAA",
    x"29187B99",
    x"2918688B",
    x"2918557F",
    x"29184275",
    x"29182F6E",
    x"29181C6A",
    x"29180967",
    x"2917F667",
    x"2917E36A",
    x"2917D06E",
    x"2917BD75",
    x"2917AA7F",
    x"2917978B",
    x"29178499",
    x"291771AA",
    x"29175EBD",
    x"29174BD2",
    x"291738EA",
    x"29172604",
    x"29171320",
    x"2917003F",
    x"2916ED60",
    x"2916DA84",
    x"2916C7AA",
    x"2916B4D2",
    x"2916A1FC",
    x"29168F29",
    x"29167C59",
    x"2916698A",
    x"291656BE",
    x"291643F4",
    x"2916312D",
    x"29161E68",
    x"29160BA6",
    x"2915F8E5",
    x"2915E627",
    x"2915D36C",
    x"2915C0B2",
    x"2915ADFC",
    x"29159B47",
    x"29158895",
    x"291575E5",
    x"29156337",
    x"2915508C",
    x"29153DE3",
    x"29152B3D",
    x"29151898",
    x"291505F6",
    x"2914F357",
    x"2914E0BA",
    x"2914CE1F",
    x"2914BB86",
    x"2914A8F0",
    x"2914965C",
    x"291483CA",
    x"2914713B",
    x"29145EAE",
    x"29144C23",
    x"2914399B",
    x"29142715",
    x"29141491",
    x"29140210",
    x"2913EF91",
    x"2913DD14",
    x"2913CA99",
    x"2913B821",
    x"2913A5AB",
    x"29139338",
    x"291380C6",
    x"29136E57",
    x"29135BEB",
    x"29134980",
    x"29133718",
    x"291324B3",
    x"2913124F",
    x"2912FFEE",
    x"2912ED8F",
    x"2912DB33",
    x"2912C8D8",
    x"2912B681",
    x"2912A42B",
    x"291291D7",
    x"29127F86",
    x"29126D38",
    x"29125AEB",
    x"291248A1",
    x"29123659",
    x"29122413",
    x"291211D0",
    x"2911FF8F",
    x"2911ED50",
    x"2911DB14",
    x"2911C8D9",
    x"2911B6A1",
    x"2911A46C",
    x"29119238",
    x"29118007",
    x"29116DD8",
    x"29115BAC",
    x"29114981",
    x"29113759",
    x"29112533",
    x"29111310",
    x"291100EF",
    x"2910EED0",
    x"2910DCB3",
    x"2910CA99",
    x"2910B880",
    x"2910A66A",
    x"29109457",
    x"29108245",
    x"29107036",
    x"29105E29",
    x"29104C1F",
    x"29103A16",
    x"29102810",
    x"2910160C",
    x"2910040B",
    x"290FF20B",
    x"290FE00E",
    x"290FCE13",
    x"290FBC1B",
    x"290FAA24",
    x"290F9830",
    x"290F863E",
    x"290F744E",
    x"290F6261",
    x"290F5076",
    x"290F3E8D",
    x"290F2CA6",
    x"290F1AC2",
    x"290F08E0",
    x"290EF700",
    x"290EE522",
    x"290ED346",
    x"290EC16D",
    x"290EAF96",
    x"290E9DC1",
    x"290E8BEE",
    x"290E7A1E",
    x"290E6850",
    x"290E5684",
    x"290E44BA",
    x"290E32F3",
    x"290E212E",
    x"290E0F6B",
    x"290DFDAA",
    x"290DEBEB",
    x"290DDA2F",
    x"290DC875",
    x"290DB6BD",
    x"290DA507",
    x"290D9353",
    x"290D81A2",
    x"290D6FF3",
    x"290D5E46",
    x"290D4C9B",
    x"290D3AF3",
    x"290D294D",
    x"290D17A9",
    x"290D0607",
    x"290CF467",
    x"290CE2CA",
    x"290CD12E",
    x"290CBF95",
    x"290CADFE",
    x"290C9C6A",
    x"290C8AD7",
    x"290C7947",
    x"290C67B9",
    x"290C562D",
    x"290C44A4",
    x"290C331C",
    x"290C2197",
    x"290C1014",
    x"290BFE93",
    x"290BED14",
    x"290BDB97",
    x"290BCA1D",
    x"290BB8A5",
    x"290BA72F",
    x"290B95BB",
    x"290B8449",
    x"290B72DA",
    x"290B616D",
    x"290B5002",
    x"290B3E99",
    x"290B2D32",
    x"290B1BCD",
    x"290B0A6B",
    x"290AF90B",
    x"290AE7AD",
    x"290AD651",
    x"290AC4F7",
    x"290AB3A0",
    x"290AA24A",
    x"290A90F7",
    x"290A7FA6",
    x"290A6E57",
    x"290A5D0B",
    x"290A4BC0",
    x"290A3A78",
    x"290A2931",
    x"290A17ED",
    x"290A06AB",
    x"2909F56C",
    x"2909E42E",
    x"2909D2F3",
    x"2909C1B9",
    x"2909B082",
    x"29099F4D",
    x"29098E1A",
    x"29097CEA",
    x"29096BBB",
    x"29095A8F",
    x"29094964",
    x"2909383C",
    x"29092716",
    x"290915F3",
    x"290904D1",
    x"2908F3B1",
    x"2908E294",
    x"2908D179",
    x"2908C060",
    x"2908AF49",
    x"29089E34",
    x"29088D21",
    x"29087C10",
    x"29086B02",
    x"290859F6",
    x"290848EC",
    x"290837E4",
    x"290826DE",
    x"290815DA",
    x"290804D8",
    x"2907F3D9",
    x"2907E2DB",
    x"2907D1E0",
    x"2907C0E7",
    x"2907AFF0",
    x"29079EFB",
    x"29078E08",
    x"29077D17",
    x"29076C29",
    x"29075B3C",
    x"29074A52",
    x"2907396A",
    x"29072883",
    x"2907179F",
    x"290706BE",
    x"2906F5DE",
    x"2906E500",
    x"2906D425",
    x"2906C34B",
    x"2906B274",
    x"2906A19E",
    x"290690CB",
    x"29067FFA",
    x"29066F2B",
    x"29065E5E",
    x"29064D94",
    x"29063CCB",
    x"29062C05",
    x"29061B40",
    x"29060A7E",
    x"2905F9BD",
    x"2905E8FF",
    x"2905D843",
    x"2905C789",
    x"2905B6D1",
    x"2905A61B",
    x"29059568",
    x"290584B6",
    x"29057407",
    x"29056359",
    x"290552AE",
    x"29054204",
    x"2905315D",
    x"290520B8",
    x"29051015",
    x"2904FF74",
    x"2904EED5",
    x"2904DE38",
    x"2904CD9E",
    x"2904BD05",
    x"2904AC6E",
    x"29049BDA",
    x"29048B47",
    x"29047AB7",
    x"29046A29",
    x"2904599D",
    x"29044912",
    x"2904388A",
    x"29042804",
    x"29041780",
    x"290406FE",
    x"2903F67E",
    x"2903E601",
    x"2903D585",
    x"2903C50B",
    x"2903B494",
    x"2903A41E",
    x"290393AB",
    x"29038339",
    x"290372CA",
    x"2903625D",
    x"290351F1",
    x"29034188",
    x"29033121",
    x"290320BC",
    x"29031059",
    x"2902FFF8",
    x"2902EF99",
    x"2902DF3C",
    x"2902CEE1",
    x"2902BE88",
    x"2902AE31",
    x"29029DDD",
    x"29028D8A",
    x"29027D39",
    x"29026CEB",
    x"29025C9E",
    x"29024C53",
    x"29023C0B",
    x"29022BC4",
    x"29021B80",
    x"29020B3D",
    x"2901FAFD",
    x"2901EABF",
    x"2901DA82",
    x"2901CA48",
    x"2901BA10",
    x"2901A9DA",
    x"290199A5",
    x"29018973",
    x"29017943",
    x"29016915",
    x"290158E9",
    x"290148BF",
    x"29013897",
    x"29012870",
    x"2901184C",
    x"2901082A",
    x"2900F80A",
    x"2900E7EC",
    x"2900D7D0",
    x"2900C7B6",
    x"2900B79E",
    x"2900A789",
    x"29009775",
    x"29008763",
    x"29007753",
    x"29006745",
    x"29005739",
    x"2900472F",
    x"29003727",
    x"29002721",
    x"2900171D",
    x"2900071B",
    x"28FFEE37",
    x"28FFCE3B",
    x"28FFAE44",
    x"28FF8E50",
    x"28FF6E60",
    x"28FF4E74",
    x"28FF2E8C",
    x"28FF0EA9",
    x"28FEEEC9",
    x"28FECEED",
    x"28FEAF15",
    x"28FE8F41",
    x"28FE6F71",
    x"28FE4FA5",
    x"28FE2FDD",
    x"28FE1019",
    x"28FDF059",
    x"28FDD09D",
    x"28FDB0E5",
    x"28FD9131",
    x"28FD7181",
    x"28FD51D5",
    x"28FD322C",
    x"28FD1288",
    x"28FCF2E8",
    x"28FCD34B",
    x"28FCB3B3",
    x"28FC941E",
    x"28FC748E",
    x"28FC5501",
    x"28FC3579",
    x"28FC15F4",
    x"28FBF673",
    x"28FBD6F6",
    x"28FBB77D",
    x"28FB9808",
    x"28FB7897",
    x"28FB592A",
    x"28FB39C1",
    x"28FB1A5C",
    x"28FAFAFB",
    x"28FADB9D",
    x"28FABC44",
    x"28FA9CEE",
    x"28FA7D9C",
    x"28FA5E4F",
    x"28FA3F05",
    x"28FA1FBF",
    x"28FA007D",
    x"28F9E13F",
    x"28F9C205",
    x"28F9A2CE",
    x"28F9839C",
    x"28F9646D",
    x"28F94543",
    x"28F9261C",
    x"28F906F9",
    x"28F8E7DA",
    x"28F8C8BF",
    x"28F8A9A8",
    x"28F88A95",
    x"28F86B85",
    x"28F84C7A",
    x"28F82D72",
    x"28F80E6F",
    x"28F7EF6F",
    x"28F7D073",
    x"28F7B17B",
    x"28F79286",
    x"28F77396",
    x"28F754A9",
    x"28F735C1",
    x"28F716DC",
    x"28F6F7FB",
    x"28F6D91E",
    x"28F6BA45",
    x"28F69B6F",
    x"28F67C9E",
    x"28F65DD0",
    x"28F63F06",
    x"28F62041",
    x"28F6017E",
    x"28F5E2C0",
    x"28F5C406",
    x"28F5A54F",
    x"28F5869C",
    x"28F567EE",
    x"28F54942",
    x"28F52A9B",
    x"28F50BF8",
    x"28F4ED58",
    x"28F4CEBC",
    x"28F4B025",
    x"28F49190",
    x"28F47300",
    x"28F45474",
    x"28F435EB",
    x"28F41766",
    x"28F3F8E5",
    x"28F3DA68",
    x"28F3BBEF",
    x"28F39D79",
    x"28F37F07",
    x"28F36099",
    x"28F3422F",
    x"28F323C9",
    x"28F30566",
    x"28F2E707",
    x"28F2C8AC",
    x"28F2AA55",
    x"28F28C02",
    x"28F26DB2",
    x"28F24F66",
    x"28F2311E",
    x"28F212DA",
    x"28F1F49A",
    x"28F1D65D",
    x"28F1B824",
    x"28F199EF",
    x"28F17BBE",
    x"28F15D90",
    x"28F13F66",
    x"28F12140",
    x"28F1031E",
    x"28F0E4FF",
    x"28F0C6E5",
    x"28F0A8CE",
    x"28F08ABA",
    x"28F06CAB",
    x"28F04E9F",
    x"28F03097",
    x"28F01293",
    x"28EFF493",
    x"28EFD696",
    x"28EFB89D",
    x"28EF9AA8",
    x"28EF7CB6",
    x"28EF5EC9",
    x"28EF40DF",
    x"28EF22F8",
    x"28EF0516",
    x"28EEE737",
    x"28EEC95C",
    x"28EEAB85",
    x"28EE8DB1",
    x"28EE6FE1",
    x"28EE5215",
    x"28EE344D",
    x"28EE1688",
    x"28EDF8C7",
    x"28EDDB0A",
    x"28EDBD50",
    x"28ED9F9B",
    x"28ED81E8",
    x"28ED643A",
    x"28ED468F",
    x"28ED28E8",
    x"28ED0B45",
    x"28ECEDA6",
    x"28ECD00A",
    x"28ECB272",
    x"28EC94DD",
    x"28EC774C",
    x"28EC59BF",
    x"28EC3C36",
    x"28EC1EB0",
    x"28EC012E",
    x"28EBE3B0",
    x"28EBC635",
    x"28EBA8BE",
    x"28EB8B4B",
    x"28EB6DDC",
    x"28EB5070",
    x"28EB3308",
    x"28EB15A3",
    x"28EAF842",
    x"28EADAE5",
    x"28EABD8B",
    x"28EAA036",
    x"28EA82E3",
    x"28EA6595",
    x"28EA484A",
    x"28EA2B03",
    x"28EA0DBF",
    x"28E9F07F",
    x"28E9D343",
    x"28E9B60A",
    x"28E998D6",
    x"28E97BA4",
    x"28E95E77",
    x"28E9414D",
    x"28E92426",
    x"28E90704",
    x"28E8E9E5",
    x"28E8CCC9",
    x"28E8AFB1",
    x"28E8929D",
    x"28E8758D",
    x"28E85880",
    x"28E83B77",
    x"28E81E71",
    x"28E8016F",
    x"28E7E471",
    x"28E7C776",
    x"28E7AA7F",
    x"28E78D8B",
    x"28E7709B",
    x"28E753AF",
    x"28E736C6",
    x"28E719E1",
    x"28E6FD00",
    x"28E6E022",
    x"28E6C348",
    x"28E6A671",
    x"28E6899E",
    x"28E66CCF",
    x"28E65003",
    x"28E6333B",
    x"28E61676",
    x"28E5F9B5",
    x"28E5DCF8",
    x"28E5C03E",
    x"28E5A388",
    x"28E586D5",
    x"28E56A26",
    x"28E54D7B",
    x"28E530D3",
    x"28E5142E",
    x"28E4F78E",
    x"28E4DAF1",
    x"28E4BE57",
    x"28E4A1C1",
    x"28E4852F",
    x"28E468A0",
    x"28E44C14",
    x"28E42F8D",
    x"28E41308",
    x"28E3F688",
    x"28E3DA0B",
    x"28E3BD91",
    x"28E3A11B",
    x"28E384A9",
    x"28E3683A",
    x"28E34BCF",
    x"28E32F67",
    x"28E31303",
    x"28E2F6A3",
    x"28E2DA46",
    x"28E2BDEC",
    x"28E2A196",
    x"28E28544",
    x"28E268F5",
    x"28E24CA9",
    x"28E23062",
    x"28E2141D",
    x"28E1F7DD",
    x"28E1DB9F",
    x"28E1BF66",
    x"28E1A32F",
    x"28E186FD",
    x"28E16ACE",
    x"28E14EA2",
    x"28E1327A",
    x"28E11655",
    x"28E0FA34",
    x"28E0DE17",
    x"28E0C1FD",
    x"28E0A5E6",
    x"28E089D3",
    x"28E06DC4",
    x"28E051B8",
    x"28E035B0",
    x"28E019AB",
    x"28DFFDA9",
    x"28DFE1AB",
    x"28DFC5B1",
    x"28DFA9BA",
    x"28DF8DC6",
    x"28DF71D6",
    x"28DF55EA",
    x"28DF3A01",
    x"28DF1E1B",
    x"28DF0239",
    x"28DEE65B",
    x"28DECA80",
    x"28DEAEA8",
    x"28DE92D4",
    x"28DE7703",
    x"28DE5B36",
    x"28DE3F6D",
    x"28DE23A6",
    x"28DE07E4",
    x"28DDEC24",
    x"28DDD069",
    x"28DDB4B0",
    x"28DD98FC",
    x"28DD7D4A",
    x"28DD619C",
    x"28DD45F2",
    x"28DD2A4B",
    x"28DD0EA7",
    x"28DCF307",
    x"28DCD76A",
    x"28DCBBD1",
    x"28DCA03B",
    x"28DC84A9",
    x"28DC691A",
    x"28DC4D8F",
    x"28DC3207",
    x"28DC1682",
    x"28DBFB01",
    x"28DBDF84",
    x"28DBC409",
    x"28DBA893",
    x"28DB8D1F",
    x"28DB71AF",
    x"28DB5643",
    x"28DB3ADA",
    x"28DB1F74",
    x"28DB0412",
    x"28DAE8B3",
    x"28DACD58",
    x"28DAB200",
    x"28DA96AB",
    x"28DA7B5A",
    x"28DA600C",
    x"28DA44C2",
    x"28DA297B",
    x"28DA0E38",
    x"28D9F2F8",
    x"28D9D7BB",
    x"28D9BC82",
    x"28D9A14C",
    x"28D98619",
    x"28D96AEA",
    x"28D94FBF",
    x"28D93496",
    x"28D91971",
    x"28D8FE50",
    x"28D8E332",
    x"28D8C817",
    x"28D8AD00",
    x"28D891EC",
    x"28D876DB",
    x"28D85BCE",
    x"28D840C4",
    x"28D825BE",
    x"28D80ABB",
    x"28D7EFBB",
    x"28D7D4BF",
    x"28D7B9C6",
    x"28D79ED1",
    x"28D783DE",
    x"28D768F0",
    x"28D74E04",
    x"28D7331C",
    x"28D71837",
    x"28D6FD56",
    x"28D6E278",
    x"28D6C79D",
    x"28D6ACC6",
    x"28D691F2",
    x"28D67722",
    x"28D65C55",
    x"28D6418B",
    x"28D626C4",
    x"28D60C01",
    x"28D5F141",
    x"28D5D685",
    x"28D5BBCB",
    x"28D5A116",
    x"28D58663",
    x"28D56BB4",
    x"28D55108",
    x"28D53660",
    x"28D51BBB",
    x"28D50119",
    x"28D4E67A",
    x"28D4CBDF",
    x"28D4B147",
    x"28D496B3",
    x"28D47C22",
    x"28D46194",
    x"28D44709",
    x"28D42C82",
    x"28D411FE",
    x"28D3F77E",
    x"28D3DD00",
    x"28D3C286",
    x"28D3A810",
    x"28D38D9C",
    x"28D3732C",
    x"28D358C0",
    x"28D33E56",
    x"28D323F0",
    x"28D3098D",
    x"28D2EF2E",
    x"28D2D4D1",
    x"28D2BA78",
    x"28D2A023",
    x"28D285D0",
    x"28D26B81",
    x"28D25136",
    x"28D236ED",
    x"28D21CA8",
    x"28D20266",
    x"28D1E827",
    x"28D1CDEC",
    x"28D1B3B4",
    x"28D1997F",
    x"28D17F4D",
    x"28D1651F",
    x"28D14AF4",
    x"28D130CC",
    x"28D116A8",
    x"28D0FC87",
    x"28D0E269",
    x"28D0C84E",
    x"28D0AE37",
    x"28D09422",
    x"28D07A12",
    x"28D06004",
    x"28D045FA",
    x"28D02BF2",
    x"28D011EF",
    x"28CFF7EE",
    x"28CFDDF1",
    x"28CFC3F7",
    x"28CFAA00",
    x"28CF900C",
    x"28CF761C",
    x"28CF5C2E",
    x"28CF4245",
    x"28CF285E",
    x"28CF0E7A",
    x"28CEF49A",
    x"28CEDABD",
    x"28CEC0E4",
    x"28CEA70D",
    x"28CE8D3A",
    x"28CE736A",
    x"28CE599D",
    x"28CE3FD3",
    x"28CE260D",
    x"28CE0C4A",
    x"28CDF28A",
    x"28CDD8CD",
    x"28CDBF14",
    x"28CDA55D",
    x"28CD8BAA",
    x"28CD71FB",
    x"28CD584E",
    x"28CD3EA4",
    x"28CD24FE",
    x"28CD0B5B",
    x"28CCF1BB",
    x"28CCD81F",
    x"28CCBE85",
    x"28CCA4EF",
    x"28CC8B5C",
    x"28CC71CC",
    x"28CC5840",
    x"28CC3EB6",
    x"28CC2530",
    x"28CC0BAD",
    x"28CBF22D",
    x"28CBD8B0",
    x"28CBBF37",
    x"28CBA5C1",
    x"28CB8C4E",
    x"28CB72DE",
    x"28CB5971",
    x"28CB4007",
    x"28CB26A1",
    x"28CB0D3E",
    x"28CAF3DD",
    x"28CADA81",
    x"28CAC127",
    x"28CAA7D0",
    x"28CA8E7D",
    x"28CA752D",
    x"28CA5BE0",
    x"28CA4296",
    x"28CA294F",
    x"28CA100B",
    x"28C9F6CB",
    x"28C9DD8E",
    x"28C9C454",
    x"28C9AB1D",
    x"28C991E9",
    x"28C978B8",
    x"28C95F8B",
    x"28C94660",
    x"28C92D39",
    x"28C91415",
    x"28C8FAF4",
    x"28C8E1D6",
    x"28C8C8BC",
    x"28C8AFA4",
    x"28C89690",
    x"28C87D7E",
    x"28C86470",
    x"28C84B65",
    x"28C8325D",
    x"28C81959",
    x"28C80057",
    x"28C7E759",
    x"28C7CE5D",
    x"28C7B565",
    x"28C79C70",
    x"28C7837E",
    x"28C76A8F",
    x"28C751A3",
    x"28C738BB",
    x"28C71FD5",
    x"28C706F3",
    x"28C6EE13",
    x"28C6D537",
    x"28C6BC5E",
    x"28C6A388",
    x"28C68AB5",
    x"28C671E5",
    x"28C65919",
    x"28C6404F",
    x"28C62789",
    x"28C60EC5",
    x"28C5F605",
    x"28C5DD48",
    x"28C5C48E",
    x"28C5ABD7",
    x"28C59323",
    x"28C57A72",
    x"28C561C4",
    x"28C54919",
    x"28C53072",
    x"28C517CD",
    x"28C4FF2C",
    x"28C4E68D",
    x"28C4CDF2",
    x"28C4B55A",
    x"28C49CC5",
    x"28C48433",
    x"28C46BA4",
    x"28C45318",
    x"28C43A8F",
    x"28C42209",
    x"28C40986",
    x"28C3F107",
    x"28C3D88A",
    x"28C3C011",
    x"28C3A79A",
    x"28C38F27",
    x"28C376B6",
    x"28C35E49",
    x"28C345DF",
    x"28C32D78",
    x"28C31513",
    x"28C2FCB2",
    x"28C2E454",
    x"28C2CBF9",
    x"28C2B3A1",
    x"28C29B4C",
    x"28C282FA",
    x"28C26AAC",
    x"28C25260",
    x"28C23A17",
    x"28C221D1",
    x"28C2098F",
    x"28C1F14F",
    x"28C1D912",
    x"28C1C0D9",
    x"28C1A8A2",
    x"28C1906E",
    x"28C1783E",
    x"28C16010",
    x"28C147E6",
    x"28C12FBE",
    x"28C1179A",
    x"28C0FF78",
    x"28C0E75A",
    x"28C0CF3F",
    x"28C0B726",
    x"28C09F11",
    x"28C086FE",
    x"28C06EEF",
    x"28C056E3",
    x"28C03ED9",
    x"28C026D3",
    x"28C00ED0",
    x"28BFF6CF",
    x"28BFDED2",
    x"28BFC6D8",
    x"28BFAEE0",
    x"28BF96EC",
    x"28BF7EFB",
    x"28BF670C",
    x"28BF4F21",
    x"28BF3738",
    x"28BF1F53",
    x"28BF0771",
    x"28BEEF91",
    x"28BED7B5",
    x"28BEBFDB",
    x"28BEA805",
    x"28BE9031",
    x"28BE7861",
    x"28BE6093",
    x"28BE48C9",
    x"28BE3101",
    x"28BE193C",
    x"28BE017B",
    x"28BDE9BC",
    x"28BDD200",
    x"28BDBA47",
    x"28BDA292",
    x"28BD8ADF",
    x"28BD732F",
    x"28BD5B82",
    x"28BD43D8",
    x"28BD2C31",
    x"28BD148D",
    x"28BCFCEC",
    x"28BCE54E",
    x"28BCCDB3",
    x"28BCB61A",
    x"28BC9E85",
    x"28BC86F3",
    x"28BC6F63",
    x"28BC57D7",
    x"28BC404D",
    x"28BC28C7",
    x"28BC1143",
    x"28BBF9C2",
    x"28BBE245",
    x"28BBCACA",
    x"28BBB352",
    x"28BB9BDD",
    x"28BB846B",
    x"28BB6CFC",
    x"28BB5590",
    x"28BB3E27",
    x"28BB26C0",
    x"28BB0F5D",
    x"28BAF7FC",
    x"28BAE09F",
    x"28BAC944",
    x"28BAB1ED",
    x"28BA9A98",
    x"28BA8346",
    x"28BA6BF7",
    x"28BA54AB",
    x"28BA3D62",
    x"28BA261C",
    x"28BA0ED8",
    x"28B9F798",
    x"28B9E05A",
    x"28B9C920",
    x"28B9B1E8",
    x"28B99AB3",
    x"28B98381",
    x"28B96C52",
    x"28B95526",
    x"28B93DFD",
    x"28B926D7",
    x"28B90FB3",
    x"28B8F893",
    x"28B8E175",
    x"28B8CA5A",
    x"28B8B343",
    x"28B89C2E",
    x"28B8851C",
    x"28B86E0C",
    x"28B85700",
    x"28B83FF7",
    x"28B828F0",
    x"28B811EC",
    x"28B7FAEC",
    x"28B7E3EE",
    x"28B7CCF3",
    x"28B7B5FA",
    x"28B79F05",
    x"28B78813",
    x"28B77123",
    x"28B75A36",
    x"28B7434D",
    x"28B72C66",
    x"28B71581",
    x"28B6FEA0",
    x"28B6E7C2",
    x"28B6D0E6",
    x"28B6BA0E",
    x"28B6A338",
    x"28B68C65",
    x"28B67595",
    x"28B65EC7",
    x"28B647FD",
    x"28B63135",
    x"28B61A71",
    x"28B603AF",
    x"28B5ECF0",
    x"28B5D634",
    x"28B5BF7A",
    x"28B5A8C4",
    x"28B59210",
    x"28B57B5F",
    x"28B564B1",
    x"28B54E06",
    x"28B5375E",
    x"28B520B8",
    x"28B50A15",
    x"28B4F376",
    x"28B4DCD9",
    x"28B4C63E",
    x"28B4AFA7",
    x"28B49912",
    x"28B48281",
    x"28B46BF2",
    x"28B45566",
    x"28B43EDD",
    x"28B42856",
    x"28B411D2",
    x"28B3FB52",
    x"28B3E4D4",
    x"28B3CE58",
    x"28B3B7E0",
    x"28B3A16A",
    x"28B38AF8",
    x"28B37488",
    x"28B35E1B",
    x"28B347B0",
    x"28B33149",
    x"28B31AE4",
    x"28B30482",
    x"28B2EE23",
    x"28B2D7C6",
    x"28B2C16D",
    x"28B2AB16",
    x"28B294C2",
    x"28B27E71",
    x"28B26822",
    x"28B251D7",
    x"28B23B8E",
    x"28B22548",
    x"28B20F05",
    x"28B1F8C4",
    x"28B1E286",
    x"28B1CC4B",
    x"28B1B613",
    x"28B19FDE",
    x"28B189AB",
    x"28B1737C",
    x"28B15D4F",
    x"28B14724",
    x"28B130FD",
    x"28B11AD8",
    x"28B104B6",
    x"28B0EE97",
    x"28B0D87A",
    x"28B0C261",
    x"28B0AC4A",
    x"28B09636",
    x"28B08024",
    x"28B06A16",
    x"28B0540A",
    x"28B03E01",
    x"28B027FA",
    x"28B011F7",
    x"28AFFBF6",
    x"28AFE5F8",
    x"28AFCFFC",
    x"28AFBA04",
    x"28AFA40E",
    x"28AF8E1B",
    x"28AF782A",
    x"28AF623D",
    x"28AF4C52",
    x"28AF3669",
    x"28AF2084",
    x"28AF0AA1",
    x"28AEF4C1",
    x"28AEDEE4",
    x"28AEC90A",
    x"28AEB332",
    x"28AE9D5D",
    x"28AE878B",
    x"28AE71BB",
    x"28AE5BEE",
    x"28AE4624",
    x"28AE305D",
    x"28AE1A98",
    x"28AE04D6",
    x"28ADEF17",
    x"28ADD95A",
    x"28ADC3A0",
    x"28ADADE9",
    x"28AD9835",
    x"28AD8283",
    x"28AD6CD4",
    x"28AD5728",
    x"28AD417E",
    x"28AD2BD8",
    x"28AD1633",
    x"28AD0092",
    x"28ACEAF3",
    x"28ACD557",
    x"28ACBFBE",
    x"28ACAA27",
    x"28AC9493",
    x"28AC7F02",
    x"28AC6974",
    x"28AC53E8",
    x"28AC3E5F",
    x"28AC28D8",
    x"28AC1355",
    x"28ABFDD3",
    x"28ABE855",
    x"28ABD2D9",
    x"28ABBD60",
    x"28ABA7EA",
    x"28AB9276",
    x"28AB7D05",
    x"28AB6797",
    x"28AB522B",
    x"28AB3CC3",
    x"28AB275C",
    x"28AB11F9",
    x"28AAFC98",
    x"28AAE73A",
    x"28AAD1DE",
    x"28AABC85",
    x"28AAA72F",
    x"28AA91DB",
    x"28AA7C8A",
    x"28AA673C",
    x"28AA51F1",
    x"28AA3CA8",
    x"28AA2761",
    x"28AA121E",
    x"28A9FCDD",
    x"28A9E79F",
    x"28A9D263",
    x"28A9BD2A",
    x"28A9A7F4",
    x"28A992C0",
    x"28A97D8F",
    x"28A96861",
    x"28A95335",
    x"28A93E0C",
    x"28A928E5",
    x"28A913C2",
    x"28A8FEA0",
    x"28A8E982",
    x"28A8D466",
    x"28A8BF4D",
    x"28A8AA36",
    x"28A89522",
    x"28A88011",
    x"28A86B02",
    x"28A855F6",
    x"28A840ED",
    x"28A82BE6",
    x"28A816E2",
    x"28A801E0",
    x"28A7ECE1",
    x"28A7D7E5",
    x"28A7C2EB",
    x"28A7ADF4",
    x"28A79900",
    x"28A7840E",
    x"28A76F1F",
    x"28A75A32",
    x"28A74548",
    x"28A73061",
    x"28A71B7C",
    x"28A7069A",
    x"28A6F1BB",
    x"28A6DCDE",
    x"28A6C803",
    x"28A6B32C",
    x"28A69E57",
    x"28A68984",
    x"28A674B4",
    x"28A65FE7",
    x"28A64B1C",
    x"28A63654",
    x"28A6218F",
    x"28A60CCC",
    x"28A5F80B",
    x"28A5E34E",
    x"28A5CE93",
    x"28A5B9DA",
    x"28A5A524",
    x"28A59071",
    x"28A57BC0",
    x"28A56712",
    x"28A55266",
    x"28A53DBD",
    x"28A52917",
    x"28A51473",
    x"28A4FFD2",
    x"28A4EB33",
    x"28A4D697",
    x"28A4C1FD",
    x"28A4AD66",
    x"28A498D2",
    x"28A48440",
    x"28A46FB1",
    x"28A45B24",
    x"28A4469A",
    x"28A43213",
    x"28A41D8E",
    x"28A4090B",
    x"28A3F48B",
    x"28A3E00E",
    x"28A3CB93",
    x"28A3B71B",
    x"28A3A2A6",
    x"28A38E33",
    x"28A379C2",
    x"28A36554",
    x"28A350E9",
    x"28A33C80",
    x"28A3281A",
    x"28A313B6",
    x"28A2FF55",
    x"28A2EAF6",
    x"28A2D69A",
    x"28A2C240",
    x"28A2ADE9",
    x"28A29995",
    x"28A28543",
    x"28A270F4",
    x"28A25CA7",
    x"28A2485C",
    x"28A23415",
    x"28A21FCF",
    x"28A20B8D",
    x"28A1F74D",
    x"28A1E30F",
    x"28A1CED4",
    x"28A1BA9B",
    x"28A1A665",
    x"28A19232",
    x"28A17E01",
    x"28A169D2",
    x"28A155A6",
    x"28A1417D",
    x"28A12D56",
    x"28A11931",
    x"28A1050F",
    x"28A0F0F0",
    x"28A0DCD3",
    x"28A0C8B9",
    x"28A0B4A1",
    x"28A0A08C",
    x"28A08C79",
    x"28A07869",
    x"28A0645B",
    x"28A0504F",
    x"28A03C47",
    x"28A02840",
    x"28A0143D",
    x"28A0003B",
    x"289FEC3D",
    x"289FD840",
    x"289FC447",
    x"289FB04F",
    x"289F9C5A",
    x"289F8868",
    x"289F7478",
    x"289F608B",
    x"289F4CA0",
    x"289F38B8",
    x"289F24D2",
    x"289F10EF",
    x"289EFD0E",
    x"289EE92F",
    x"289ED553",
    x"289EC17A",
    x"289EADA3",
    x"289E99CF",
    x"289E85FD",
    x"289E722D",
    x"289E5E60",
    x"289E4A96",
    x"289E36CD",
    x"289E2308",
    x"289E0F45",
    x"289DFB84",
    x"289DE7C6",
    x"289DD40A",
    x"289DC051",
    x"289DAC9A",
    x"289D98E6",
    x"289D8534",
    x"289D7184",
    x"289D5DD7",
    x"289D4A2D",
    x"289D3685",
    x"289D22DF",
    x"289D0F3C",
    x"289CFB9B",
    x"289CE7FD",
    x"289CD461",
    x"289CC0C8",
    x"289CAD31",
    x"289C999D",
    x"289C860B",
    x"289C727B",
    x"289C5EEE",
    x"289C4B64",
    x"289C37DB",
    x"289C2456",
    x"289C10D2",
    x"289BFD51",
    x"289BE9D3",
    x"289BD657",
    x"289BC2DD",
    x"289BAF66",
    x"289B9BF2",
    x"289B887F",
    x"289B750F",
    x"289B61A2",
    x"289B4E37",
    x"289B3ACE",
    x"289B2768",
    x"289B1405",
    x"289B00A3",
    x"289AED44",
    x"289AD9E8",
    x"289AC68E",
    x"289AB336",
    x"289A9FE1",
    x"289A8C8E",
    x"289A793E",
    x"289A65F0",
    x"289A52A5",
    x"289A3F5B",
    x"289A2C15",
    x"289A18D0",
    x"289A058F",
    x"2899F24F",
    x"2899DF12",
    x"2899CBD7",
    x"2899B89F",
    x"2899A569",
    x"28999236",
    x"28997F05",
    x"28996BD6",
    x"289958AA",
    x"28994580",
    x"28993258",
    x"28991F33",
    x"28990C10",
    x"2898F8F0",
    x"2898E5D2",
    x"2898D2B7",
    x"2898BF9D",
    x"2898AC87",
    x"28989972",
    x"28988660",
    x"28987351",
    x"28986044",
    x"28984D39",
    x"28983A30",
    x"2898272A",
    x"28981426",
    x"28980125",
    x"2897EE26",
    x"2897DB2A",
    x"2897C82F",
    x"2897B538",
    x"2897A242",
    x"28978F4F",
    x"28977C5E",
    x"28976970",
    x"28975684",
    x"2897439A",
    x"289730B3",
    x"28971DCE",
    x"28970AEC",
    x"2896F80B",
    x"2896E52E",
    x"2896D252",
    x"2896BF79",
    x"2896ACA2",
    x"289699CE",
    x"289686FC",
    x"2896742C",
    x"2896615F",
    x"28964E94",
    x"28963BCB",
    x"28962905",
    x"28961641",
    x"2896037F",
    x"2895F0C0",
    x"2895DE03",
    x"2895CB48",
    x"2895B890",
    x"2895A5DA",
    x"28959327",
    x"28958075",
    x"28956DC7",
    x"28955B1A",
    x"28954870",
    x"289535C8",
    x"28952322",
    x"2895107F",
    x"2894FDDE",
    x"2894EB40",
    x"2894D8A3",
    x"2894C60A",
    x"2894B372",
    x"2894A0DD",
    x"28948E4A",
    x"28947BB9",
    x"2894692B",
    x"2894569F",
    x"28944415",
    x"2894318E",
    x"28941F09",
    x"28940C86",
    x"2893FA06",
    x"2893E787",
    x"2893D50C",
    x"2893C292",
    x"2893B01B",
    x"28939DA6",
    x"28938B34",
    x"289378C3",
    x"28936655",
    x"289353EA",
    x"28934180",
    x"28932F19",
    x"28931CB5",
    x"28930A52",
    x"2892F7F2",
    x"2892E594",
    x"2892D339",
    x"2892C0DF",
    x"2892AE89",
    x"28929C34",
    x"289289E1",
    x"28927791",
    x"28926544",
    x"289252F8",
    x"289240AF",
    x"28922E68",
    x"28921C23",
    x"289209E1",
    x"2891F7A1",
    x"2891E563",
    x"2891D327",
    x"2891C0EE",
    x"2891AEB7",
    x"28919C82",
    x"28918A50",
    x"28917820",
    x"289165F2",
    x"289153C6",
    x"2891419D",
    x"28912F76",
    x"28911D51",
    x"28910B2F",
    x"2890F90E",
    x"2890E6F0",
    x"2890D4D5",
    x"2890C2BB",
    x"2890B0A4",
    x"28909E8F",
    x"28908C7C",
    x"28907A6C",
    x"2890685E",
    x"28905652",
    x"28904448",
    x"28903241",
    x"2890203C",
    x"28900E39",
    x"288FFC38",
    x"288FEA3A",
    x"288FD83D",
    x"288FC644",
    x"288FB44C",
    x"288FA257",
    x"288F9063",
    x"288F7E72",
    x"288F6C84",
    x"288F5A97",
    x"288F48AD",
    x"288F36C5",
    x"288F24DF",
    x"288F12FC",
    x"288F011B",
    x"288EEF3C",
    x"288EDD5F",
    x"288ECB84",
    x"288EB9AC",
    x"288EA7D6",
    x"288E9602",
    x"288E8430",
    x"288E7261",
    x"288E6094",
    x"288E4EC9",
    x"288E3D00",
    x"288E2B3A",
    x"288E1975",
    x"288E07B3",
    x"288DF5F3",
    x"288DE436",
    x"288DD27A",
    x"288DC0C1",
    x"288DAF0A",
    x"288D9D55",
    x"288D8BA3",
    x"288D79F2",
    x"288D6844",
    x"288D5698",
    x"288D44EF",
    x"288D3347",
    x"288D21A2",
    x"288D0FFF",
    x"288CFE5E",
    x"288CECBF",
    x"288CDB23",
    x"288CC988",
    x"288CB7F0",
    x"288CA65A",
    x"288C94C7",
    x"288C8335",
    x"288C71A6",
    x"288C6019",
    x"288C4E8E",
    x"288C3D05",
    x"288C2B7F",
    x"288C19FA",
    x"288C0878",
    x"288BF6F8",
    x"288BE57A",
    x"288BD3FF",
    x"288BC285",
    x"288BB10E",
    x"288B9F99",
    x"288B8E26",
    x"288B7CB6",
    x"288B6B47",
    x"288B59DB",
    x"288B4871",
    x"288B3709",
    x"288B25A3",
    x"288B143F",
    x"288B02DE",
    x"288AF17E",
    x"288AE021",
    x"288ACEC6",
    x"288ABD6E",
    x"288AAC17",
    x"288A9AC3",
    x"288A8970",
    x"288A7820",
    x"288A66D2",
    x"288A5587",
    x"288A443D",
    x"288A32F6",
    x"288A21B0",
    x"288A106D",
    x"2889FF2C",
    x"2889EDED",
    x"2889DCB1",
    x"2889CB76",
    x"2889BA3E",
    x"2889A908",
    x"288997D4",
    x"288986A2",
    x"28897572",
    x"28896444",
    x"28895319",
    x"288941EF",
    x"288930C8",
    x"28891FA3",
    x"28890E80",
    x"2888FD60",
    x"2888EC41",
    x"2888DB25",
    x"2888CA0A",
    x"2888B8F2",
    x"2888A7DC",
    x"288896C8",
    x"288885B6",
    x"288874A7",
    x"28886399",
    x"2888528E",
    x"28884185",
    x"2888307D",
    x"28881F78",
    x"28880E76",
    x"2887FD75",
    x"2887EC76",
    x"2887DB7A",
    x"2887CA7F",
    x"2887B987",
    x"2887A891",
    x"2887979D",
    x"288786AB",
    x"288775BB",
    x"288764CE",
    x"288753E2",
    x"288742F9",
    x"28873211",
    x"2887212C",
    x"28871049",
    x"2886FF68",
    x"2886EE89",
    x"2886DDAC",
    x"2886CCD2",
    x"2886BBF9",
    x"2886AB23",
    x"28869A4E",
    x"2886897C",
    x"288678AC",
    x"288667DE",
    x"28865712",
    x"28864648",
    x"28863580",
    x"288624BB",
    x"288613F7",
    x"28860336",
    x"2885F277",
    x"2885E1B9",
    x"2885D0FE",
    x"2885C045",
    x"2885AF8E",
    x"28859ED9",
    x"28858E26",
    x"28857D76",
    x"28856CC7",
    x"28855C1A",
    x"28854B70",
    x"28853AC8",
    x"28852A21",
    x"2885197D",
    x"288508DB",
    x"2884F83B",
    x"2884E79D",
    x"2884D701",
    x"2884C667",
    x"2884B5CF",
    x"2884A53A",
    x"288494A6",
    x"28848414",
    x"28847385",
    x"288462F8",
    x"2884526C",
    x"288441E3",
    x"2884315C",
    x"288420D7",
    x"28841054",
    x"2883FFD3",
    x"2883EF54",
    x"2883DED7",
    x"2883CE5C",
    x"2883BDE3",
    x"2883AD6C",
    x"28839CF8",
    x"28838C85",
    x"28837C15",
    x"28836BA6",
    x"28835B3A",
    x"28834ACF",
    x"28833A67",
    x"28832A01",
    x"2883199C",
    x"2883093A",
    x"2882F8DA",
    x"2882E87C",
    x"2882D820",
    x"2882C7C6",
    x"2882B76E",
    x"2882A718",
    x"288296C4",
    x"28828673",
    x"28827623",
    x"288265D5",
    x"28825589",
    x"28824540",
    x"288234F8",
    x"288224B2",
    x"2882146F",
    x"2882042D",
    x"2881F3EE",
    x"2881E3B0",
    x"2881D375",
    x"2881C33B",
    x"2881B304",
    x"2881A2CF",
    x"2881929B",
    x"2881826A",
    x"2881723B",
    x"2881620D",
    x"288151E2",
    x"288141B9",
    x"28813192",
    x"2881216D",
    x"28811149",
    x"28810128",
    x"2880F109",
    x"2880E0EC",
    x"2880D0D1",
    x"2880C0B8",
    x"2880B0A1",
    x"2880A08C",
    x"28809079",
    x"28808068",
    x"28807058",
    x"2880604B",
    x"28805040",
    x"28804037",
    x"28803030",
    x"2880202B",
    x"28801028",
    x"28800027",
    x"287FE050",
    x"287FC056",
    x"287FA060",
    x"287F806E",
    x"287F6080",
    x"287F4096",
    x"287F20B0",
    x"287F00CE",
    x"287EE0F0",
    x"287EC116",
    x"287EA140",
    x"287E816E",
    x"287E619F",
    x"287E41D5",
    x"287E220F",
    x"287E024D",
    x"287DE28E",
    x"287DC2D4",
    x"287DA31E",
    x"287D836B",
    x"287D63BD",
    x"287D4412",
    x"287D246C",
    x"287D04C9",
    x"287CE52B",
    x"287CC590",
    x"287CA5F9",
    x"287C8666",
    x"287C66D8",
    x"287C474D",
    x"287C27C6",
    x"287C0843",
    x"287BE8C4",
    x"287BC948",
    x"287BA9D1",
    x"287B8A5E",
    x"287B6AEF",
    x"287B4B83",
    x"287B2C1C",
    x"287B0CB8",
    x"287AED59",
    x"287ACDFD",
    x"287AAEA5",
    x"287A8F51",
    x"287A7001",
    x"287A50B5",
    x"287A316D",
    x"287A1229",
    x"2879F2E9",
    x"2879D3AC",
    x"2879B474",
    x"2879953F",
    x"2879760E",
    x"287956E2",
    x"287937B9",
    x"28791894",
    x"2878F973",
    x"2878DA55",
    x"2878BB3C",
    x"28789C26",
    x"28787D15",
    x"28785E07",
    x"28783EFD",
    x"28781FF7",
    x"287800F5",
    x"2877E1F7",
    x"2877C2FD",
    x"2877A406",
    x"28778514",
    x"28776625",
    x"2877473A",
    x"28772853",
    x"28770970",
    x"2876EA91",
    x"2876CBB6",
    x"2876ACDE",
    x"28768E0A",
    x"28766F3B",
    x"2876506F",
    x"287631A6",
    x"287612E2",
    x"2875F422",
    x"2875D565",
    x"2875B6AC",
    x"287597F7",
    x"28757946",
    x"28755A99",
    x"28753BF0",
    x"28751D4A",
    x"2874FEA8",
    x"2874E00B",
    x"2874C170",
    x"2874A2DA",
    x"28748448",
    x"287465B9",
    x"2874472E",
    x"287428A7",
    x"28740A24",
    x"2873EBA5",
    x"2873CD29",
    x"2873AEB1",
    x"2873903E",
    x"287371CD",
    x"28735361",
    x"287334F9",
    x"28731694",
    x"2872F833",
    x"2872D9D6",
    x"2872BB7C",
    x"28729D27",
    x"28727ED5",
    x"28726087",
    x"2872423D",
    x"287223F7",
    x"287205B4",
    x"2871E775",
    x"2871C93A",
    x"2871AB03",
    x"28718CCF",
    x"28716EA0",
    x"28715074",
    x"2871324C",
    x"28711427",
    x"2870F607",
    x"2870D7EA",
    x"2870B9D1",
    x"28709BBB",
    x"28707DAA",
    x"28705F9C",
    x"28704192",
    x"2870238B",
    x"28700589",
    x"286FE78A",
    x"286FC98F",
    x"286FAB98",
    x"286F8DA4",
    x"286F6FB4",
    x"286F51C8",
    x"286F33E0",
    x"286F15FB",
    x"286EF81A",
    x"286EDA3D",
    x"286EBC64",
    x"286E9E8E",
    x"286E80BC",
    x"286E62EE",
    x"286E4523",
    x"286E275D",
    x"286E099A",
    x"286DEBDA",
    x"286DCE1F",
    x"286DB067",
    x"286D92B2",
    x"286D7502",
    x"286D5755",
    x"286D39AC",
    x"286D1C07",
    x"286CFE65",
    x"286CE0C7",
    x"286CC32D",
    x"286CA596",
    x"286C8804",
    x"286C6A74",
    x"286C4CE9",
    x"286C2F61",
    x"286C11DD",
    x"286BF45D",
    x"286BD6E0",
    x"286BB967",
    x"286B9BF2",
    x"286B7E80",
    x"286B6112",
    x"286B43A8",
    x"286B2641",
    x"286B08DE",
    x"286AEB7F",
    x"286ACE23",
    x"286AB0CB",
    x"286A9377",
    x"286A7626",
    x"286A58DA",
    x"286A3B90",
    x"286A1E4B",
    x"286A0109",
    x"2869E3CA",
    x"2869C690",
    x"2869A959",
    x"28698C25",
    x"28696EF6",
    x"286951CA",
    x"286934A1",
    x"2869177D",
    x"2868FA5B",
    x"2868DD3E",
    x"2868C024",
    x"2868A30E",
    x"286885FB",
    x"286868EC",
    x"28684BE1",
    x"28682ED9",
    x"286811D5",
    x"2867F4D5",
    x"2867D7D8",
    x"2867BADF",
    x"28679DE9",
    x"286780F8",
    x"28676409",
    x"2867471F",
    x"28672A37",
    x"28670D54",
    x"2866F074",
    x"2866D398",
    x"2866B6BF",
    x"286699EA",
    x"28667D19",
    x"2866604B",
    x"28664381",
    x"286626BA",
    x"286609F7",
    x"2865ED38",
    x"2865D07C",
    x"2865B3C3",
    x"2865970F",
    x"28657A5E",
    x"28655DB0",
    x"28654106",
    x"28652460",
    x"286507BD",
    x"2864EB1E",
    x"2864CE82",
    x"2864B1EA",
    x"28649556",
    x"286478C5",
    x"28645C38",
    x"00000000"
  );

begin

  p_mem_read : process (clk) begin
    if rising_edge(clk) then
      data_out <= mem(to_integer(unsigned(address)));
    end if;
  end process;

end architecture;
