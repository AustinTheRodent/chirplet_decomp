
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sine_rom is
  port
  (
    clk       : in  std_logic;
    address   : in  std_logic_vector(15 downto 0);
    data_out  : out std_logic_vector(31 downto 0)
  );
end entity;

architecture rtl of sine_rom is

  constant C_DATA_WIDTH  : integer := 32;
  constant C_ADDR_WIDTH  : integer := 16;

  constant RAM_DEPTH :integer := 2**C_ADDR_WIDTH;

  type RAM is array (integer range <>) of std_logic_vector (C_DATA_WIDTH-1 downto 0);
  signal mem : RAM (0 to RAM_DEPTH-1) :=
  (
    x"00000000",
    x"38C90FDB",
    x"39490FDB",
    x"3996CBE4",
    x"39C90FDA",
    x"39FB53D1",
    x"3A16CBE3",
    x"3A2FEDDE",
    x"3A490FD9",
    x"3A6231D4",
    x"3A7B53CF",
    x"3A8A3AE5",
    x"3A96CBE2",
    x"3AA35CDF",
    x"3AAFEDDC",
    x"3ABC7ED9",
    x"3AC90FD5",
    x"3AD5A0D2",
    x"3AE231CF",
    x"3AEEC2CB",
    x"3AFB53C7",
    x"3B03F262",
    x"3B0A3AE0",
    x"3B10835D",
    x"3B16CBDB",
    x"3B1D1459",
    x"3B235CD7",
    x"3B29A554",
    x"3B2FEDD1",
    x"3B36364F",
    x"3B3C7ECC",
    x"3B42C749",
    x"3B490FC6",
    x"3B4F5843",
    x"3B55A0C0",
    x"3B5BE93C",
    x"3B6231B9",
    x"3B687A35",
    x"3B6EC2B1",
    x"3B750B2D",
    x"3B7B53A9",
    x"3B80CE12",
    x"3B83F250",
    x"3B87168E",
    x"3B8A3ACB",
    x"3B8D5F09",
    x"3B908346",
    x"3B93A784",
    x"3B96CBC1",
    x"3B99EFFE",
    x"3B9D143B",
    x"3BA03878",
    x"3BA35CB5",
    x"3BA680F2",
    x"3BA9A52F",
    x"3BACC96B",
    x"3BAFEDA8",
    x"3BB311E4",
    x"3BB63621",
    x"3BB95A5D",
    x"3BBC7E99",
    x"3BBFA2D5",
    x"3BC2C711",
    x"3BC5EB4C",
    x"3BC90F88",
    x"3BCC33C3",
    x"3BCF57FF",
    x"3BD27C3A",
    x"3BD5A075",
    x"3BD8C4B0",
    x"3BDBE8EB",
    x"3BDF0D26",
    x"3BE23160",
    x"3BE5559B",
    x"3BE879D5",
    x"3BEB9E0F",
    x"3BEEC249",
    x"3BF1E683",
    x"3BF50ABD",
    x"3BF82EF6",
    x"3BFB5330",
    x"3BFE7769",
    x"3C00CDD1",
    x"3C025FEE",
    x"3C03F20A",
    x"3C058426",
    x"3C071643",
    x"3C08A85F",
    x"3C0A3A7B",
    x"3C0BCC97",
    x"3C0D5EB3",
    x"3C0EF0CF",
    x"3C1082EA",
    x"3C121506",
    x"3C13A722",
    x"3C15393D",
    x"3C16CB58",
    x"3C185D74",
    x"3C19EF8F",
    x"3C1B81AA",
    x"3C1D13C5",
    x"3C1EA5E0",
    x"3C2037FB",
    x"3C21CA16",
    x"3C235C30",
    x"3C24EE4B",
    x"3C268065",
    x"3C281280",
    x"3C29A49A",
    x"3C2B36B4",
    x"3C2CC8CE",
    x"3C2E5AE8",
    x"3C2FED02",
    x"3C317F1B",
    x"3C331135",
    x"3C34A34F",
    x"3C363568",
    x"3C37C781",
    x"3C39599A",
    x"3C3AEBB4",
    x"3C3C7DCC",
    x"3C3E0FE5",
    x"3C3FA1FE",
    x"3C413417",
    x"3C42C62F",
    x"3C445847",
    x"3C45EA60",
    x"3C477C78",
    x"3C490E90",
    x"3C4AA0A8",
    x"3C4C32C0",
    x"3C4DC4D7",
    x"3C4F56EF",
    x"3C50E906",
    x"3C527B1D",
    x"3C540D35",
    x"3C559F4C",
    x"3C573162",
    x"3C58C379",
    x"3C5A5590",
    x"3C5BE7A6",
    x"3C5D79BD",
    x"3C5F0BD3",
    x"3C609DE9",
    x"3C622FFF",
    x"3C63C215",
    x"3C65542B",
    x"3C66E640",
    x"3C687856",
    x"3C6A0A6B",
    x"3C6B9C80",
    x"3C6D2E95",
    x"3C6EC0AA",
    x"3C7052BF",
    x"3C71E4D3",
    x"3C7376E7",
    x"3C7508FC",
    x"3C769B10",
    x"3C782D24",
    x"3C79BF38",
    x"3C7B514B",
    x"3C7CE35F",
    x"3C7E7572",
    x"3C8003C3",
    x"3C80CCCC",
    x"3C8195D6",
    x"3C825EDF",
    x"3C8327E8",
    x"3C83F0F2",
    x"3C84B9FB",
    x"3C858304",
    x"3C864C0D",
    x"3C871516",
    x"3C87DE1E",
    x"3C88A727",
    x"3C897030",
    x"3C8A3938",
    x"3C8B0241",
    x"3C8BCB49",
    x"3C8C9452",
    x"3C8D5D5A",
    x"3C8E2662",
    x"3C8EEF6A",
    x"3C8FB872",
    x"3C90817A",
    x"3C914A82",
    x"3C921389",
    x"3C92DC91",
    x"3C93A599",
    x"3C946EA0",
    x"3C9537A7",
    x"3C9600AF",
    x"3C96C9B6",
    x"3C9792BD",
    x"3C985BC4",
    x"3C9924CB",
    x"3C99EDD2",
    x"3C9AB6D8",
    x"3C9B7FDF",
    x"3C9C48E6",
    x"3C9D11EC",
    x"3C9DDAF2",
    x"3C9EA3F9",
    x"3C9F6CFF",
    x"3CA03605",
    x"3CA0FF0B",
    x"3CA1C811",
    x"3CA29116",
    x"3CA35A1C",
    x"3CA42322",
    x"3CA4EC27",
    x"3CA5B52C",
    x"3CA67E32",
    x"3CA74737",
    x"3CA8103C",
    x"3CA8D941",
    x"3CA9A246",
    x"3CAA6B4B",
    x"3CAB344F",
    x"3CABFD54",
    x"3CACC658",
    x"3CAD8F5D",
    x"3CAE5861",
    x"3CAF2165",
    x"3CAFEA69",
    x"3CB0B36D",
    x"3CB17C71",
    x"3CB24575",
    x"3CB30E78",
    x"3CB3D77C",
    x"3CB4A07F",
    x"3CB56982",
    x"3CB63286",
    x"3CB6FB89",
    x"3CB7C48C",
    x"3CB88D8E",
    x"3CB95691",
    x"3CBA1F94",
    x"3CBAE896",
    x"3CBBB199",
    x"3CBC7A9B",
    x"3CBD439D",
    x"3CBE0C9F",
    x"3CBED5A1",
    x"3CBF9EA3",
    x"3CC067A5",
    x"3CC130A6",
    x"3CC1F9A8",
    x"3CC2C2A9",
    x"3CC38BAA",
    x"3CC454AB",
    x"3CC51DAC",
    x"3CC5E6AD",
    x"3CC6AFAE",
    x"3CC778AF",
    x"3CC841AF",
    x"3CC90AB0",
    x"3CC9D3B0",
    x"3CCA9CB0",
    x"3CCB65B0",
    x"3CCC2EB0",
    x"3CCCF7B0",
    x"3CCDC0B0",
    x"3CCE89AF",
    x"3CCF52AF",
    x"3CD01BAE",
    x"3CD0E4AD",
    x"3CD1ADAC",
    x"3CD276AB",
    x"3CD33FAA",
    x"3CD408A9",
    x"3CD4D1A7",
    x"3CD59AA6",
    x"3CD663A4",
    x"3CD72CA2",
    x"3CD7F5A0",
    x"3CD8BE9E",
    x"3CD9879C",
    x"3CDA5099",
    x"3CDB1997",
    x"3CDBE294",
    x"3CDCAB91",
    x"3CDD748F",
    x"3CDE3D8C",
    x"3CDF0688",
    x"3CDFCF85",
    x"3CE09882",
    x"3CE1617E",
    x"3CE22A7A",
    x"3CE2F377",
    x"3CE3BC73",
    x"3CE4856E",
    x"3CE54E6A",
    x"3CE61766",
    x"3CE6E061",
    x"3CE7A95D",
    x"3CE87258",
    x"3CE93B53",
    x"3CEA044E",
    x"3CEACD49",
    x"3CEB9643",
    x"3CEC5F3E",
    x"3CED2838",
    x"3CEDF132",
    x"3CEEBA2C",
    x"3CEF8326",
    x"3CF04C20",
    x"3CF1151A",
    x"3CF1DE13",
    x"3CF2A70D",
    x"3CF37006",
    x"3CF438FF",
    x"3CF501F8",
    x"3CF5CAF0",
    x"3CF693E9",
    x"3CF75CE2",
    x"3CF825DA",
    x"3CF8EED2",
    x"3CF9B7CA",
    x"3CFA80C2",
    x"3CFB49BA",
    x"3CFC12B1",
    x"3CFCDBA9",
    x"3CFDA4A0",
    x"3CFE6D97",
    x"3CFF368E",
    x"3CFFFF85",
    x"3D00643E",
    x"3D00C8B9",
    x"3D012D34",
    x"3D0191AF",
    x"3D01F62A",
    x"3D025AA5",
    x"3D02BF20",
    x"3D03239B",
    x"3D038815",
    x"3D03EC90",
    x"3D04510B",
    x"3D04B585",
    x"3D0519FF",
    x"3D057E7A",
    x"3D05E2F4",
    x"3D06476E",
    x"3D06ABE8",
    x"3D071062",
    x"3D0774DC",
    x"3D07D956",
    x"3D083DCF",
    x"3D08A249",
    x"3D0906C3",
    x"3D096B3C",
    x"3D09CFB6",
    x"3D0A342F",
    x"3D0A98A8",
    x"3D0AFD21",
    x"3D0B619A",
    x"3D0BC613",
    x"3D0C2A8C",
    x"3D0C8F05",
    x"3D0CF37E",
    x"3D0D57F6",
    x"3D0DBC6F",
    x"3D0E20E7",
    x"3D0E8560",
    x"3D0EE9D8",
    x"3D0F4E50",
    x"3D0FB2C8",
    x"3D101740",
    x"3D107BB8",
    x"3D10E030",
    x"3D1144A8",
    x"3D11A920",
    x"3D120D97",
    x"3D12720F",
    x"3D12D686",
    x"3D133AFE",
    x"3D139F75",
    x"3D1403EC",
    x"3D146863",
    x"3D14CCDA",
    x"3D153151",
    x"3D1595C8",
    x"3D15FA3F",
    x"3D165EB5",
    x"3D16C32C",
    x"3D1727A2",
    x"3D178C18",
    x"3D17F08F",
    x"3D185505",
    x"3D18B97B",
    x"3D191DF1",
    x"3D198267",
    x"3D19E6DD",
    x"3D1A4B52",
    x"3D1AAFC8",
    x"3D1B143D",
    x"3D1B78B3",
    x"3D1BDD28",
    x"3D1C419D",
    x"3D1CA613",
    x"3D1D0A88",
    x"3D1D6EFD",
    x"3D1DD372",
    x"3D1E37E6",
    x"3D1E9C5B",
    x"3D1F00D0",
    x"3D1F6544",
    x"3D1FC9B8",
    x"3D202E2D",
    x"3D2092A1",
    x"3D20F715",
    x"3D215B89",
    x"3D21BFFD",
    x"3D222471",
    x"3D2288E4",
    x"3D22ED58",
    x"3D2351CB",
    x"3D23B63F",
    x"3D241AB2",
    x"3D247F25",
    x"3D24E399",
    x"3D25480C",
    x"3D25AC7E",
    x"3D2610F1",
    x"3D267564",
    x"3D26D9D7",
    x"3D273E49",
    x"3D27A2BC",
    x"3D28072E",
    x"3D286BA0",
    x"3D28D012",
    x"3D293484",
    x"3D2998F6",
    x"3D29FD68",
    x"3D2A61DA",
    x"3D2AC64B",
    x"3D2B2ABD",
    x"3D2B8F2E",
    x"3D2BF39F",
    x"3D2C5811",
    x"3D2CBC82",
    x"3D2D20F3",
    x"3D2D8564",
    x"3D2DE9D4",
    x"3D2E4E45",
    x"3D2EB2B6",
    x"3D2F1726",
    x"3D2F7B96",
    x"3D2FE007",
    x"3D304477",
    x"3D30A8E7",
    x"3D310D57",
    x"3D3171C6",
    x"3D31D636",
    x"3D323AA6",
    x"3D329F15",
    x"3D330385",
    x"3D3367F4",
    x"3D33CC63",
    x"3D3430D2",
    x"3D349541",
    x"3D34F9B0",
    x"3D355E1F",
    x"3D35C28D",
    x"3D3626FC",
    x"3D368B6A",
    x"3D36EFD9",
    x"3D375447",
    x"3D37B8B5",
    x"3D381D23",
    x"3D388191",
    x"3D38E5FE",
    x"3D394A6C",
    x"3D39AEDA",
    x"3D3A1347",
    x"3D3A77B4",
    x"3D3ADC22",
    x"3D3B408F",
    x"3D3BA4FC",
    x"3D3C0968",
    x"3D3C6DD5",
    x"3D3CD242",
    x"3D3D36AE",
    x"3D3D9B1B",
    x"3D3DFF87",
    x"3D3E63F3",
    x"3D3EC85F",
    x"3D3F2CCB",
    x"3D3F9137",
    x"3D3FF5A3",
    x"3D405A0E",
    x"3D40BE7A",
    x"3D4122E5",
    x"3D418750",
    x"3D41EBBB",
    x"3D425026",
    x"3D42B491",
    x"3D4318FC",
    x"3D437D67",
    x"3D43E1D1",
    x"3D44463C",
    x"3D44AAA6",
    x"3D450F10",
    x"3D45737A",
    x"3D45D7E4",
    x"3D463C4E",
    x"3D46A0B8",
    x"3D470521",
    x"3D47698B",
    x"3D47CDF4",
    x"3D48325D",
    x"3D4896C7",
    x"3D48FB30",
    x"3D495F98",
    x"3D49C401",
    x"3D4A286A",
    x"3D4A8CD2",
    x"3D4AF13B",
    x"3D4B55A3",
    x"3D4BBA0B",
    x"3D4C1E73",
    x"3D4C82DB",
    x"3D4CE743",
    x"3D4D4BAA",
    x"3D4DB012",
    x"3D4E1479",
    x"3D4E78E1",
    x"3D4EDD48",
    x"3D4F41AF",
    x"3D4FA616",
    x"3D500A7C",
    x"3D506EE3",
    x"3D50D34A",
    x"3D5137B0",
    x"3D519C16",
    x"3D52007C",
    x"3D5264E2",
    x"3D52C948",
    x"3D532DAE",
    x"3D539214",
    x"3D53F679",
    x"3D545ADF",
    x"3D54BF44",
    x"3D5523A9",
    x"3D55880E",
    x"3D55EC73",
    x"3D5650D8",
    x"3D56B53C",
    x"3D5719A1",
    x"3D577E05",
    x"3D57E269",
    x"3D5846CD",
    x"3D58AB31",
    x"3D590F95",
    x"3D5973F9",
    x"3D59D85C",
    x"3D5A3CC0",
    x"3D5AA123",
    x"3D5B0586",
    x"3D5B69E9",
    x"3D5BCE4C",
    x"3D5C32AF",
    x"3D5C9712",
    x"3D5CFB74",
    x"3D5D5FD7",
    x"3D5DC439",
    x"3D5E289B",
    x"3D5E8CFD",
    x"3D5EF15F",
    x"3D5F55C0",
    x"3D5FBA22",
    x"3D601E83",
    x"3D6082E5",
    x"3D60E746",
    x"3D614BA7",
    x"3D61B008",
    x"3D621469",
    x"3D6278C9",
    x"3D62DD2A",
    x"3D63418A",
    x"3D63A5EA",
    x"3D640A4A",
    x"3D646EAA",
    x"3D64D30A",
    x"3D65376A",
    x"3D659BC9",
    x"3D660029",
    x"3D666488",
    x"3D66C8E7",
    x"3D672D46",
    x"3D6791A5",
    x"3D67F604",
    x"3D685A62",
    x"3D68BEC1",
    x"3D69231F",
    x"3D69877D",
    x"3D69EBDB",
    x"3D6A5039",
    x"3D6AB496",
    x"3D6B18F4",
    x"3D6B7D51",
    x"3D6BE1AF",
    x"3D6C460C",
    x"3D6CAA69",
    x"3D6D0EC6",
    x"3D6D7323",
    x"3D6DD77F",
    x"3D6E3BDC",
    x"3D6EA038",
    x"3D6F0494",
    x"3D6F68F0",
    x"3D6FCD4C",
    x"3D7031A8",
    x"3D709603",
    x"3D70FA5E",
    x"3D715EBA",
    x"3D71C315",
    x"3D722770",
    x"3D728BCB",
    x"3D72F025",
    x"3D735480",
    x"3D73B8DA",
    x"3D741D35",
    x"3D74818F",
    x"3D74E5E9",
    x"3D754A42",
    x"3D75AE9C",
    x"3D7612F6",
    x"3D76774F",
    x"3D76DBA8",
    x"3D774001",
    x"3D77A45A",
    x"3D7808B3",
    x"3D786D0C",
    x"3D78D164",
    x"3D7935BC",
    x"3D799A15",
    x"3D79FE6D",
    x"3D7A62C5",
    x"3D7AC71C",
    x"3D7B2B74",
    x"3D7B8FCB",
    x"3D7BF422",
    x"3D7C587A",
    x"3D7CBCD1",
    x"3D7D2127",
    x"3D7D857E",
    x"3D7DE9D5",
    x"3D7E4E2B",
    x"3D7EB281",
    x"3D7F16D7",
    x"3D7F7B2D",
    x"3D7FDF83",
    x"3D8021EC",
    x"3D805417",
    x"3D808642",
    x"3D80B86C",
    x"3D80EA97",
    x"3D811CC1",
    x"3D814EEB",
    x"3D818116",
    x"3D81B340",
    x"3D81E56A",
    x"3D821794",
    x"3D8249BE",
    x"3D827BE8",
    x"3D82AE11",
    x"3D82E03B",
    x"3D831265",
    x"3D83448E",
    x"3D8376B8",
    x"3D83A8E1",
    x"3D83DB0A",
    x"3D840D34",
    x"3D843F5D",
    x"3D847186",
    x"3D84A3AF",
    x"3D84D5D8",
    x"3D850801",
    x"3D853A29",
    x"3D856C52",
    x"3D859E7B",
    x"3D85D0A3",
    x"3D8602CC",
    x"3D8634F4",
    x"3D86671C",
    x"3D869944",
    x"3D86CB6C",
    x"3D86FD94",
    x"3D872FBC",
    x"3D8761E4",
    x"3D87940C",
    x"3D87C634",
    x"3D87F85B",
    x"3D882A83",
    x"3D885CAA",
    x"3D888ED2",
    x"3D88C0F9",
    x"3D88F320",
    x"3D892547",
    x"3D89576E",
    x"3D898995",
    x"3D89BBBC",
    x"3D89EDE3",
    x"3D8A200A",
    x"3D8A5230",
    x"3D8A8457",
    x"3D8AB67D",
    x"3D8AE8A4",
    x"3D8B1ACA",
    x"3D8B4CF0",
    x"3D8B7F16",
    x"3D8BB13C",
    x"3D8BE362",
    x"3D8C1588",
    x"3D8C47AE",
    x"3D8C79D4",
    x"3D8CABF9",
    x"3D8CDE1F",
    x"3D8D1044",
    x"3D8D426A",
    x"3D8D748F",
    x"3D8DA6B4",
    x"3D8DD8D9",
    x"3D8E0AFE",
    x"3D8E3D23",
    x"3D8E6F48",
    x"3D8EA16D",
    x"3D8ED391",
    x"3D8F05B6",
    x"3D8F37DA",
    x"3D8F69FF",
    x"3D8F9C23",
    x"3D8FCE47",
    x"3D90006C",
    x"3D903290",
    x"3D9064B4",
    x"3D9096D8",
    x"3D90C8FB",
    x"3D90FB1F",
    x"3D912D43",
    x"3D915F66",
    x"3D91918A",
    x"3D91C3AD",
    x"3D91F5D0",
    x"3D9227F4",
    x"3D925A17",
    x"3D928C3A",
    x"3D92BE5D",
    x"3D92F07F",
    x"3D9322A2",
    x"3D9354C5",
    x"3D9386E7",
    x"3D93B90A",
    x"3D93EB2C",
    x"3D941D4F",
    x"3D944F71",
    x"3D948193",
    x"3D94B3B5",
    x"3D94E5D7",
    x"3D9517F9",
    x"3D954A1B",
    x"3D957C3C",
    x"3D95AE5E",
    x"3D95E07F",
    x"3D9612A1",
    x"3D9644C2",
    x"3D9676E3",
    x"3D96A905",
    x"3D96DB26",
    x"3D970D47",
    x"3D973F67",
    x"3D977188",
    x"3D97A3A9",
    x"3D97D5CA",
    x"3D9807EA",
    x"3D983A0A",
    x"3D986C2B",
    x"3D989E4B",
    x"3D98D06B",
    x"3D99028B",
    x"3D9934AB",
    x"3D9966CB",
    x"3D9998EB",
    x"3D99CB0A",
    x"3D99FD2A",
    x"3D9A2F4A",
    x"3D9A6169",
    x"3D9A9388",
    x"3D9AC5A7",
    x"3D9AF7C7",
    x"3D9B29E6",
    x"3D9B5C05",
    x"3D9B8E23",
    x"3D9BC042",
    x"3D9BF261",
    x"3D9C247F",
    x"3D9C569E",
    x"3D9C88BC",
    x"3D9CBADA",
    x"3D9CECF9",
    x"3D9D1F17",
    x"3D9D5135",
    x"3D9D8353",
    x"3D9DB570",
    x"3D9DE78E",
    x"3D9E19AC",
    x"3D9E4BC9",
    x"3D9E7DE7",
    x"3D9EB004",
    x"3D9EE221",
    x"3D9F143E",
    x"3D9F465B",
    x"3D9F7878",
    x"3D9FAA95",
    x"3D9FDCB2",
    x"3DA00ECF",
    x"3DA040EB",
    x"3DA07308",
    x"3DA0A524",
    x"3DA0D740",
    x"3DA1095C",
    x"3DA13B78",
    x"3DA16D94",
    x"3DA19FB0",
    x"3DA1D1CC",
    x"3DA203E8",
    x"3DA23603",
    x"3DA2681F",
    x"3DA29A3A",
    x"3DA2CC55",
    x"3DA2FE71",
    x"3DA3308C",
    x"3DA362A7",
    x"3DA394C2",
    x"3DA3C6DC",
    x"3DA3F8F7",
    x"3DA42B12",
    x"3DA45D2C",
    x"3DA48F47",
    x"3DA4C161",
    x"3DA4F37B",
    x"3DA52595",
    x"3DA557AF",
    x"3DA589C9",
    x"3DA5BBE3",
    x"3DA5EDFD",
    x"3DA62016",
    x"3DA65230",
    x"3DA68449",
    x"3DA6B663",
    x"3DA6E87C",
    x"3DA71A95",
    x"3DA74CAE",
    x"3DA77EC7",
    x"3DA7B0E0",
    x"3DA7E2F8",
    x"3DA81511",
    x"3DA84729",
    x"3DA87942",
    x"3DA8AB5A",
    x"3DA8DD72",
    x"3DA90F8A",
    x"3DA941A2",
    x"3DA973BA",
    x"3DA9A5D2",
    x"3DA9D7EA",
    x"3DAA0A01",
    x"3DAA3C19",
    x"3DAA6E30",
    x"3DAAA048",
    x"3DAAD25F",
    x"3DAB0476",
    x"3DAB368D",
    x"3DAB68A4",
    x"3DAB9ABA",
    x"3DABCCD1",
    x"3DABFEE8",
    x"3DAC30FE",
    x"3DAC6314",
    x"3DAC952B",
    x"3DACC741",
    x"3DACF957",
    x"3DAD2B6D",
    x"3DAD5D83",
    x"3DAD8F98",
    x"3DADC1AE",
    x"3DADF3C3",
    x"3DAE25D9",
    x"3DAE57EE",
    x"3DAE8A03",
    x"3DAEBC18",
    x"3DAEEE2D",
    x"3DAF2042",
    x"3DAF5257",
    x"3DAF846C",
    x"3DAFB680",
    x"3DAFE895",
    x"3DB01AA9",
    x"3DB04CBD",
    x"3DB07ED2",
    x"3DB0B0E6",
    x"3DB0E2FA",
    x"3DB1150D",
    x"3DB14721",
    x"3DB17935",
    x"3DB1AB48",
    x"3DB1DD5C",
    x"3DB20F6F",
    x"3DB24182",
    x"3DB27395",
    x"3DB2A5A8",
    x"3DB2D7BB",
    x"3DB309CE",
    x"3DB33BE0",
    x"3DB36DF3",
    x"3DB3A005",
    x"3DB3D218",
    x"3DB4042A",
    x"3DB4363C",
    x"3DB4684E",
    x"3DB49A60",
    x"3DB4CC72",
    x"3DB4FE83",
    x"3DB53095",
    x"3DB562A6",
    x"3DB594B8",
    x"3DB5C6C9",
    x"3DB5F8DA",
    x"3DB62AEB",
    x"3DB65CFC",
    x"3DB68F0D",
    x"3DB6C11D",
    x"3DB6F32E",
    x"3DB7253E",
    x"3DB7574F",
    x"3DB7895F",
    x"3DB7BB6F",
    x"3DB7ED7F",
    x"3DB81F8F",
    x"3DB8519F",
    x"3DB883AF",
    x"3DB8B5BE",
    x"3DB8E7CE",
    x"3DB919DD",
    x"3DB94BEC",
    x"3DB97DFB",
    x"3DB9B00A",
    x"3DB9E219",
    x"3DBA1428",
    x"3DBA4637",
    x"3DBA7845",
    x"3DBAAA54",
    x"3DBADC62",
    x"3DBB0E70",
    x"3DBB407E",
    x"3DBB728C",
    x"3DBBA49A",
    x"3DBBD6A8",
    x"3DBC08B6",
    x"3DBC3AC3",
    x"3DBC6CD1",
    x"3DBC9EDE",
    x"3DBCD0EB",
    x"3DBD02F8",
    x"3DBD3505",
    x"3DBD6712",
    x"3DBD991F",
    x"3DBDCB2C",
    x"3DBDFD38",
    x"3DBE2F45",
    x"3DBE6151",
    x"3DBE935D",
    x"3DBEC569",
    x"3DBEF775",
    x"3DBF2981",
    x"3DBF5B8D",
    x"3DBF8D98",
    x"3DBFBFA4",
    x"3DBFF1AF",
    x"3DC023BA",
    x"3DC055C6",
    x"3DC087D1",
    x"3DC0B9DC",
    x"3DC0EBE6",
    x"3DC11DF1",
    x"3DC14FFC",
    x"3DC18206",
    x"3DC1B410",
    x"3DC1E61B",
    x"3DC21825",
    x"3DC24A2F",
    x"3DC27C39",
    x"3DC2AE42",
    x"3DC2E04C",
    x"3DC31255",
    x"3DC3445F",
    x"3DC37668",
    x"3DC3A871",
    x"3DC3DA7A",
    x"3DC40C83",
    x"3DC43E8C",
    x"3DC47095",
    x"3DC4A29D",
    x"3DC4D4A6",
    x"3DC506AE",
    x"3DC538B6",
    x"3DC56ABE",
    x"3DC59CC6",
    x"3DC5CECE",
    x"3DC600D6",
    x"3DC632DE",
    x"3DC664E5",
    x"3DC696ED",
    x"3DC6C8F4",
    x"3DC6FAFB",
    x"3DC72D02",
    x"3DC75F09",
    x"3DC79110",
    x"3DC7C316",
    x"3DC7F51D",
    x"3DC82723",
    x"3DC8592A",
    x"3DC88B30",
    x"3DC8BD36",
    x"3DC8EF3C",
    x"3DC92142",
    x"3DC95347",
    x"3DC9854D",
    x"3DC9B752",
    x"3DC9E958",
    x"3DCA1B5D",
    x"3DCA4D62",
    x"3DCA7F67",
    x"3DCAB16C",
    x"3DCAE371",
    x"3DCB1575",
    x"3DCB477A",
    x"3DCB797E",
    x"3DCBAB82",
    x"3DCBDD86",
    x"3DCC0F8A",
    x"3DCC418E",
    x"3DCC7392",
    x"3DCCA596",
    x"3DCCD799",
    x"3DCD099C",
    x"3DCD3BA0",
    x"3DCD6DA3",
    x"3DCD9FA6",
    x"3DCDD1A9",
    x"3DCE03AB",
    x"3DCE35AE",
    x"3DCE67B1",
    x"3DCE99B3",
    x"3DCECBB5",
    x"3DCEFDB7",
    x"3DCF2FB9",
    x"3DCF61BB",
    x"3DCF93BD",
    x"3DCFC5BF",
    x"3DCFF7C0",
    x"3DD029C2",
    x"3DD05BC3",
    x"3DD08DC4",
    x"3DD0BFC5",
    x"3DD0F1C6",
    x"3DD123C7",
    x"3DD155C7",
    x"3DD187C8",
    x"3DD1B9C8",
    x"3DD1EBC8",
    x"3DD21DC8",
    x"3DD24FC8",
    x"3DD281C8",
    x"3DD2B3C8",
    x"3DD2E5C8",
    x"3DD317C7",
    x"3DD349C7",
    x"3DD37BC6",
    x"3DD3ADC5",
    x"3DD3DFC4",
    x"3DD411C3",
    x"3DD443C1",
    x"3DD475C0",
    x"3DD4A7BE",
    x"3DD4D9BD",
    x"3DD50BBB",
    x"3DD53DB9",
    x"3DD56FB7",
    x"3DD5A1B5",
    x"3DD5D3B3",
    x"3DD605B0",
    x"3DD637AE",
    x"3DD669AB",
    x"3DD69BA8",
    x"3DD6CDA5",
    x"3DD6FFA2",
    x"3DD7319F",
    x"3DD7639C",
    x"3DD79598",
    x"3DD7C795",
    x"3DD7F991",
    x"3DD82B8D",
    x"3DD85D89",
    x"3DD88F85",
    x"3DD8C181",
    x"3DD8F37C",
    x"3DD92578",
    x"3DD95773",
    x"3DD9896E",
    x"3DD9BB69",
    x"3DD9ED64",
    x"3DDA1F5F",
    x"3DDA515A",
    x"3DDA8354",
    x"3DDAB54F",
    x"3DDAE749",
    x"3DDB1943",
    x"3DDB4B3D",
    x"3DDB7D37",
    x"3DDBAF31",
    x"3DDBE12B",
    x"3DDC1324",
    x"3DDC451E",
    x"3DDC7717",
    x"3DDCA910",
    x"3DDCDB09",
    x"3DDD0D02",
    x"3DDD3EFB",
    x"3DDD70F3",
    x"3DDDA2EC",
    x"3DDDD4E4",
    x"3DDE06DC",
    x"3DDE38D4",
    x"3DDE6ACC",
    x"3DDE9CC4",
    x"3DDECEBC",
    x"3DDF00B3",
    x"3DDF32AB",
    x"3DDF64A2",
    x"3DDF9699",
    x"3DDFC890",
    x"3DDFFA87",
    x"3DE02C7D",
    x"3DE05E74",
    x"3DE0906A",
    x"3DE0C261",
    x"3DE0F457",
    x"3DE1264D",
    x"3DE15843",
    x"3DE18A39",
    x"3DE1BC2E",
    x"3DE1EE24",
    x"3DE22019",
    x"3DE2520E",
    x"3DE28403",
    x"3DE2B5F8",
    x"3DE2E7ED",
    x"3DE319E2",
    x"3DE34BD6",
    x"3DE37DCB",
    x"3DE3AFBF",
    x"3DE3E1B3",
    x"3DE413A7",
    x"3DE4459B",
    x"3DE4778F",
    x"3DE4A982",
    x"3DE4DB76",
    x"3DE50D69",
    x"3DE53F5C",
    x"3DE5714F",
    x"3DE5A342",
    x"3DE5D535",
    x"3DE60727",
    x"3DE6391A",
    x"3DE66B0C",
    x"3DE69CFE",
    x"3DE6CEF0",
    x"3DE700E2",
    x"3DE732D4",
    x"3DE764C6",
    x"3DE796B7",
    x"3DE7C8A9",
    x"3DE7FA9A",
    x"3DE82C8B",
    x"3DE85E7C",
    x"3DE8906D",
    x"3DE8C25D",
    x"3DE8F44E",
    x"3DE9263E",
    x"3DE9582E",
    x"3DE98A1F",
    x"3DE9BC0E",
    x"3DE9EDFE",
    x"3DEA1FEE",
    x"3DEA51DE",
    x"3DEA83CD",
    x"3DEAB5BC",
    x"3DEAE7AB",
    x"3DEB199A",
    x"3DEB4B89",
    x"3DEB7D78",
    x"3DEBAF66",
    x"3DEBE155",
    x"3DEC1343",
    x"3DEC4531",
    x"3DEC771F",
    x"3DECA90D",
    x"3DECDAFB",
    x"3DED0CE8",
    x"3DED3ED5",
    x"3DED70C3",
    x"3DEDA2B0",
    x"3DEDD49D",
    x"3DEE068A",
    x"3DEE3876",
    x"3DEE6A63",
    x"3DEE9C4F",
    x"3DEECE3C",
    x"3DEF0028",
    x"3DEF3214",
    x"3DEF63FF",
    x"3DEF95EB",
    x"3DEFC7D7",
    x"3DEFF9C2",
    x"3DF02BAD",
    x"3DF05D98",
    x"3DF08F83",
    x"3DF0C16E",
    x"3DF0F359",
    x"3DF12543",
    x"3DF1572E",
    x"3DF18918",
    x"3DF1BB02",
    x"3DF1ECEC",
    x"3DF21ED6",
    x"3DF250BF",
    x"3DF282A9",
    x"3DF2B492",
    x"3DF2E67C",
    x"3DF31865",
    x"3DF34A4E",
    x"3DF37C36",
    x"3DF3AE1F",
    x"3DF3E007",
    x"3DF411F0",
    x"3DF443D8",
    x"3DF475C0",
    x"3DF4A7A8",
    x"3DF4D990",
    x"3DF50B77",
    x"3DF53D5F",
    x"3DF56F46",
    x"3DF5A12D",
    x"3DF5D314",
    x"3DF604FB",
    x"3DF636E2",
    x"3DF668C8",
    x"3DF69AAF",
    x"3DF6CC95",
    x"3DF6FE7B",
    x"3DF73061",
    x"3DF76247",
    x"3DF7942C",
    x"3DF7C612",
    x"3DF7F7F7",
    x"3DF829DD",
    x"3DF85BC2",
    x"3DF88DA7",
    x"3DF8BF8B",
    x"3DF8F170",
    x"3DF92354",
    x"3DF95539",
    x"3DF9871D",
    x"3DF9B901",
    x"3DF9EAE5",
    x"3DFA1CC8",
    x"3DFA4EAC",
    x"3DFA808F",
    x"3DFAB273",
    x"3DFAE456",
    x"3DFB1639",
    x"3DFB481C",
    x"3DFB79FE",
    x"3DFBABE1",
    x"3DFBDDC3",
    x"3DFC0FA5",
    x"3DFC4187",
    x"3DFC7369",
    x"3DFCA54B",
    x"3DFCD72D",
    x"3DFD090E",
    x"3DFD3AEF",
    x"3DFD6CD1",
    x"3DFD9EB2",
    x"3DFDD092",
    x"3DFE0273",
    x"3DFE3454",
    x"3DFE6634",
    x"3DFE9814",
    x"3DFEC9F4",
    x"3DFEFBD4",
    x"3DFF2DB4",
    x"3DFF5F94",
    x"3DFF9173",
    x"3DFFC352",
    x"3DFFF531",
    x"3E001388",
    x"3E002C78",
    x"3E004567",
    x"3E005E56",
    x"3E007745",
    x"3E009035",
    x"3E00A924",
    x"3E00C213",
    x"3E00DB01",
    x"3E00F3F0",
    x"3E010CDF",
    x"3E0125CE",
    x"3E013EBC",
    x"3E0157AB",
    x"3E017099",
    x"3E018987",
    x"3E01A276",
    x"3E01BB64",
    x"3E01D452",
    x"3E01ED40",
    x"3E02062E",
    x"3E021F1C",
    x"3E02380A",
    x"3E0250F7",
    x"3E0269E5",
    x"3E0282D2",
    x"3E029BC0",
    x"3E02B4AD",
    x"3E02CD9B",
    x"3E02E688",
    x"3E02FF75",
    x"3E031862",
    x"3E03314F",
    x"3E034A3C",
    x"3E036329",
    x"3E037C16",
    x"3E039502",
    x"3E03ADEF",
    x"3E03C6DB",
    x"3E03DFC8",
    x"3E03F8B4",
    x"3E0411A0",
    x"3E042A8D",
    x"3E044379",
    x"3E045C65",
    x"3E047551",
    x"3E048E3D",
    x"3E04A729",
    x"3E04C014",
    x"3E04D900",
    x"3E04F1EB",
    x"3E050AD7",
    x"3E0523C2",
    x"3E053CAE",
    x"3E055599",
    x"3E056E84",
    x"3E05876F",
    x"3E05A05A",
    x"3E05B945",
    x"3E05D230",
    x"3E05EB1B",
    x"3E060405",
    x"3E061CF0",
    x"3E0635DB",
    x"3E064EC5",
    x"3E0667AF",
    x"3E06809A",
    x"3E069984",
    x"3E06B26E",
    x"3E06CB58",
    x"3E06E442",
    x"3E06FD2C",
    x"3E071616",
    x"3E072EFF",
    x"3E0747E9",
    x"3E0760D2",
    x"3E0779BC",
    x"3E0792A5",
    x"3E07AB8F",
    x"3E07C478",
    x"3E07DD61",
    x"3E07F64A",
    x"3E080F33",
    x"3E08281C",
    x"3E084105",
    x"3E0859ED",
    x"3E0872D6",
    x"3E088BBF",
    x"3E08A4A7",
    x"3E08BD90",
    x"3E08D678",
    x"3E08EF60",
    x"3E090848",
    x"3E092130",
    x"3E093A18",
    x"3E095300",
    x"3E096BE8",
    x"3E0984D0",
    x"3E099DB7",
    x"3E09B69F",
    x"3E09CF86",
    x"3E09E86E",
    x"3E0A0155",
    x"3E0A1A3C",
    x"3E0A3324",
    x"3E0A4C0B",
    x"3E0A64F2",
    x"3E0A7DD9",
    x"3E0A96BF",
    x"3E0AAFA6",
    x"3E0AC88D",
    x"3E0AE173",
    x"3E0AFA5A",
    x"3E0B1340",
    x"3E0B2C27",
    x"3E0B450D",
    x"3E0B5DF3",
    x"3E0B76D9",
    x"3E0B8FBF",
    x"3E0BA8A5",
    x"3E0BC18B",
    x"3E0BDA71",
    x"3E0BF356",
    x"3E0C0C3C",
    x"3E0C2521",
    x"3E0C3E07",
    x"3E0C56EC",
    x"3E0C6FD1",
    x"3E0C88B6",
    x"3E0CA19B",
    x"3E0CBA80",
    x"3E0CD365",
    x"3E0CEC4A",
    x"3E0D052F",
    x"3E0D1E13",
    x"3E0D36F8",
    x"3E0D4FDC",
    x"3E0D68C1",
    x"3E0D81A5",
    x"3E0D9A89",
    x"3E0DB36D",
    x"3E0DCC51",
    x"3E0DE535",
    x"3E0DFE19",
    x"3E0E16FD",
    x"3E0E2FE1",
    x"3E0E48C4",
    x"3E0E61A8",
    x"3E0E7A8B",
    x"3E0E936F",
    x"3E0EAC52",
    x"3E0EC535",
    x"3E0EDE18",
    x"3E0EF6FB",
    x"3E0F0FDE",
    x"3E0F28C1",
    x"3E0F41A4",
    x"3E0F5A86",
    x"3E0F7369",
    x"3E0F8C4B",
    x"3E0FA52E",
    x"3E0FBE10",
    x"3E0FD6F2",
    x"3E0FEFD5",
    x"3E1008B7",
    x"3E102199",
    x"3E103A7B",
    x"3E10535C",
    x"3E106C3E",
    x"3E108520",
    x"3E109E01",
    x"3E10B6E3",
    x"3E10CFC4",
    x"3E10E8A5",
    x"3E110186",
    x"3E111A68",
    x"3E113349",
    x"3E114C2A",
    x"3E11650A",
    x"3E117DEB",
    x"3E1196CC",
    x"3E11AFAC",
    x"3E11C88D",
    x"3E11E16D",
    x"3E11FA4E",
    x"3E12132E",
    x"3E122C0E",
    x"3E1244EE",
    x"3E125DCE",
    x"3E1276AE",
    x"3E128F8E",
    x"3E12A86D",
    x"3E12C14D",
    x"3E12DA2C",
    x"3E12F30C",
    x"3E130BEB",
    x"3E1324CA",
    x"3E133DAA",
    x"3E135689",
    x"3E136F68",
    x"3E138847",
    x"3E13A125",
    x"3E13BA04",
    x"3E13D2E3",
    x"3E13EBC1",
    x"3E1404A0",
    x"3E141D7E",
    x"3E14365C",
    x"3E144F3B",
    x"3E146819",
    x"3E1480F7",
    x"3E1499D5",
    x"3E14B2B2",
    x"3E14CB90",
    x"3E14E46E",
    x"3E14FD4B",
    x"3E151629",
    x"3E152F06",
    x"3E1547E4",
    x"3E1560C1",
    x"3E15799E",
    x"3E15927B",
    x"3E15AB58",
    x"3E15C435",
    x"3E15DD11",
    x"3E15F5EE",
    x"3E160ECB",
    x"3E1627A7",
    x"3E164083",
    x"3E165960",
    x"3E16723C",
    x"3E168B18",
    x"3E16A3F4",
    x"3E16BCD0",
    x"3E16D5AC",
    x"3E16EE88",
    x"3E170763",
    x"3E17203F",
    x"3E17391A",
    x"3E1751F6",
    x"3E176AD1",
    x"3E1783AC",
    x"3E179C87",
    x"3E17B562",
    x"3E17CE3D",
    x"3E17E718",
    x"3E17FFF3",
    x"3E1818CE",
    x"3E1831A8",
    x"3E184A83",
    x"3E18635D",
    x"3E187C37",
    x"3E189511",
    x"3E18ADEC",
    x"3E18C6C6",
    x"3E18DFA0",
    x"3E18F879",
    x"3E191153",
    x"3E192A2D",
    x"3E194306",
    x"3E195BE0",
    x"3E1974B9",
    x"3E198D92",
    x"3E19A66C",
    x"3E19BF45",
    x"3E19D81E",
    x"3E19F0F7",
    x"3E1A09CF",
    x"3E1A22A8",
    x"3E1A3B81",
    x"3E1A5459",
    x"3E1A6D32",
    x"3E1A860A",
    x"3E1A9EE2",
    x"3E1AB7BB",
    x"3E1AD093",
    x"3E1AE96B",
    x"3E1B0242",
    x"3E1B1B1A",
    x"3E1B33F2",
    x"3E1B4CCA",
    x"3E1B65A1",
    x"3E1B7E79",
    x"3E1B9750",
    x"3E1BB027",
    x"3E1BC8FE",
    x"3E1BE1D5",
    x"3E1BFAAC",
    x"3E1C1383",
    x"3E1C2C5A",
    x"3E1C4530",
    x"3E1C5E07",
    x"3E1C76DE",
    x"3E1C8FB4",
    x"3E1CA88A",
    x"3E1CC160",
    x"3E1CDA36",
    x"3E1CF30D",
    x"3E1D0BE2",
    x"3E1D24B8",
    x"3E1D3D8E",
    x"3E1D5664",
    x"3E1D6F39",
    x"3E1D880F",
    x"3E1DA0E4",
    x"3E1DB9B9",
    x"3E1DD28E",
    x"3E1DEB63",
    x"3E1E0438",
    x"3E1E1D0D",
    x"3E1E35E2",
    x"3E1E4EB7",
    x"3E1E678B",
    x"3E1E8060",
    x"3E1E9934",
    x"3E1EB208",
    x"3E1ECADD",
    x"3E1EE3B1",
    x"3E1EFC85",
    x"3E1F1559",
    x"3E1F2E2C",
    x"3E1F4700",
    x"3E1F5FD4",
    x"3E1F78A7",
    x"3E1F917B",
    x"3E1FAA4E",
    x"3E1FC321",
    x"3E1FDBF4",
    x"3E1FF4C8",
    x"3E200D9A",
    x"3E20266D",
    x"3E203F40",
    x"3E205813",
    x"3E2070E5",
    x"3E2089B8",
    x"3E20A28A",
    x"3E20BB5C",
    x"3E20D42F",
    x"3E20ED01",
    x"3E2105D3",
    x"3E211EA5",
    x"3E213776",
    x"3E215048",
    x"3E21691A",
    x"3E2181EB",
    x"3E219ABD",
    x"3E21B38E",
    x"3E21CC5F",
    x"3E21E530",
    x"3E21FE01",
    x"3E2216D2",
    x"3E222FA3",
    x"3E224874",
    x"3E226144",
    x"3E227A15",
    x"3E2292E5",
    x"3E22ABB6",
    x"3E22C486",
    x"3E22DD56",
    x"3E22F626",
    x"3E230EF6",
    x"3E2327C6",
    x"3E234095",
    x"3E235965",
    x"3E237235",
    x"3E238B04",
    x"3E23A3D3",
    x"3E23BCA3",
    x"3E23D572",
    x"3E23EE41",
    x"3E240710",
    x"3E241FDF",
    x"3E2438AD",
    x"3E24517C",
    x"3E246A4B",
    x"3E248319",
    x"3E249BE7",
    x"3E24B4B6",
    x"3E24CD84",
    x"3E24E652",
    x"3E24FF20",
    x"3E2517EE",
    x"3E2530BC",
    x"3E254989",
    x"3E256257",
    x"3E257B24",
    x"3E2593F2",
    x"3E25ACBF",
    x"3E25C58C",
    x"3E25DE59",
    x"3E25F726",
    x"3E260FF3",
    x"3E2628C0",
    x"3E26418C",
    x"3E265A59",
    x"3E267325",
    x"3E268BF2",
    x"3E26A4BE",
    x"3E26BD8A",
    x"3E26D656",
    x"3E26EF22",
    x"3E2707EE",
    x"3E2720BA",
    x"3E273985",
    x"3E275251",
    x"3E276B1C",
    x"3E2783E8",
    x"3E279CB3",
    x"3E27B57E",
    x"3E27CE49",
    x"3E27E714",
    x"3E27FFDF",
    x"3E2818AA",
    x"3E283174",
    x"3E284A3F",
    x"3E286309",
    x"3E287BD4",
    x"3E28949E",
    x"3E28AD68",
    x"3E28C632",
    x"3E28DEFC",
    x"3E28F7C6",
    x"3E291090",
    x"3E292959",
    x"3E294223",
    x"3E295AEC",
    x"3E2973B6",
    x"3E298C7F",
    x"3E29A548",
    x"3E29BE11",
    x"3E29D6DA",
    x"3E29EFA3",
    x"3E2A086B",
    x"3E2A2134",
    x"3E2A39FD",
    x"3E2A52C5",
    x"3E2A6B8D",
    x"3E2A8456",
    x"3E2A9D1E",
    x"3E2AB5E6",
    x"3E2ACEAE",
    x"3E2AE775",
    x"3E2B003D",
    x"3E2B1905",
    x"3E2B31CC",
    x"3E2B4A93",
    x"3E2B635B",
    x"3E2B7C22",
    x"3E2B94E9",
    x"3E2BADB0",
    x"3E2BC677",
    x"3E2BDF3E",
    x"3E2BF804",
    x"3E2C10CB",
    x"3E2C2991",
    x"3E2C4258",
    x"3E2C5B1E",
    x"3E2C73E4",
    x"3E2C8CAA",
    x"3E2CA570",
    x"3E2CBE36",
    x"3E2CD6FB",
    x"3E2CEFC1",
    x"3E2D0887",
    x"3E2D214C",
    x"3E2D3A11",
    x"3E2D52D6",
    x"3E2D6B9C",
    x"3E2D8461",
    x"3E2D9D25",
    x"3E2DB5EA",
    x"3E2DCEAF",
    x"3E2DE773",
    x"3E2E0038",
    x"3E2E18FC",
    x"3E2E31C1",
    x"3E2E4A85",
    x"3E2E6349",
    x"3E2E7C0D",
    x"3E2E94D1",
    x"3E2EAD94",
    x"3E2EC658",
    x"3E2EDF1B",
    x"3E2EF7DF",
    x"3E2F10A2",
    x"3E2F2965",
    x"3E2F4228",
    x"3E2F5AEB",
    x"3E2F73AE",
    x"3E2F8C71",
    x"3E2FA534",
    x"3E2FBDF6",
    x"3E2FD6B9",
    x"3E2FEF7B",
    x"3E30083D",
    x"3E302100",
    x"3E3039C2",
    x"3E305284",
    x"3E306B45",
    x"3E308407",
    x"3E309CC9",
    x"3E30B58A",
    x"3E30CE4C",
    x"3E30E70D",
    x"3E30FFCE",
    x"3E31188F",
    x"3E313150",
    x"3E314A11",
    x"3E3162D2",
    x"3E317B92",
    x"3E319453",
    x"3E31AD13",
    x"3E31C5D4",
    x"3E31DE94",
    x"3E31F754",
    x"3E321014",
    x"3E3228D4",
    x"3E324194",
    x"3E325A54",
    x"3E327313",
    x"3E328BD3",
    x"3E32A492",
    x"3E32BD51",
    x"3E32D610",
    x"3E32EECF",
    x"3E33078E",
    x"3E33204D",
    x"3E33390C",
    x"3E3351CB",
    x"3E336A89",
    x"3E338348",
    x"3E339C06",
    x"3E33B4C4",
    x"3E33CD82",
    x"3E33E640",
    x"3E33FEFE",
    x"3E3417BC",
    x"3E343079",
    x"3E344937",
    x"3E3461F4",
    x"3E347AB2",
    x"3E34936F",
    x"3E34AC2C",
    x"3E34C4E9",
    x"3E34DDA6",
    x"3E34F662",
    x"3E350F1F",
    x"3E3527DC",
    x"3E354098",
    x"3E355954",
    x"3E357211",
    x"3E358ACD",
    x"3E35A389",
    x"3E35BC45",
    x"3E35D501",
    x"3E35EDBC",
    x"3E360678",
    x"3E361F33",
    x"3E3637EF",
    x"3E3650AA",
    x"3E366965",
    x"3E368220",
    x"3E369ADB",
    x"3E36B396",
    x"3E36CC50",
    x"3E36E50B",
    x"3E36FDC5",
    x"3E371680",
    x"3E372F3A",
    x"3E3747F4",
    x"3E3760AE",
    x"3E377968",
    x"3E379222",
    x"3E37AADC",
    x"3E37C395",
    x"3E37DC4F",
    x"3E37F508",
    x"3E380DC1",
    x"3E38267A",
    x"3E383F33",
    x"3E3857EC",
    x"3E3870A5",
    x"3E38895E",
    x"3E38A217",
    x"3E38BACF",
    x"3E38D387",
    x"3E38EC40",
    x"3E3904F8",
    x"3E391DB0",
    x"3E393668",
    x"3E394F20",
    x"3E3967D7",
    x"3E39808F",
    x"3E399946",
    x"3E39B1FE",
    x"3E39CAB5",
    x"3E39E36C",
    x"3E39FC23",
    x"3E3A14DA",
    x"3E3A2D91",
    x"3E3A4647",
    x"3E3A5EFE",
    x"3E3A77B4",
    x"3E3A906B",
    x"3E3AA921",
    x"3E3AC1D7",
    x"3E3ADA8D",
    x"3E3AF343",
    x"3E3B0BF9",
    x"3E3B24AF",
    x"3E3B3D64",
    x"3E3B561A",
    x"3E3B6ECF",
    x"3E3B8784",
    x"3E3BA039",
    x"3E3BB8EE",
    x"3E3BD1A3",
    x"3E3BEA58",
    x"3E3C030D",
    x"3E3C1BC1",
    x"3E3C3476",
    x"3E3C4D2A",
    x"3E3C65DE",
    x"3E3C7E92",
    x"3E3C9746",
    x"3E3CAFFA",
    x"3E3CC8AE",
    x"3E3CE161",
    x"3E3CFA15",
    x"3E3D12C8",
    x"3E3D2B7C",
    x"3E3D442F",
    x"3E3D5CE2",
    x"3E3D7595",
    x"3E3D8E48",
    x"3E3DA6FA",
    x"3E3DBFAD",
    x"3E3DD860",
    x"3E3DF112",
    x"3E3E09C4",
    x"3E3E2276",
    x"3E3E3B28",
    x"3E3E53DA",
    x"3E3E6C8C",
    x"3E3E853E",
    x"3E3E9DEF",
    x"3E3EB6A1",
    x"3E3ECF52",
    x"3E3EE804",
    x"3E3F00B5",
    x"3E3F1966",
    x"3E3F3217",
    x"3E3F4AC7",
    x"3E3F6378",
    x"3E3F7C29",
    x"3E3F94D9",
    x"3E3FAD89",
    x"3E3FC639",
    x"3E3FDEEA",
    x"3E3FF79A",
    x"3E401049",
    x"3E4028F9",
    x"3E4041A9",
    x"3E405A58",
    x"3E407308",
    x"3E408BB7",
    x"3E40A466",
    x"3E40BD15",
    x"3E40D5C4",
    x"3E40EE73",
    x"3E410722",
    x"3E411FD0",
    x"3E41387F",
    x"3E41512D",
    x"3E4169DB",
    x"3E418289",
    x"3E419B37",
    x"3E41B3E5",
    x"3E41CC93",
    x"3E41E541",
    x"3E41FDEE",
    x"3E42169B",
    x"3E422F49",
    x"3E4247F6",
    x"3E4260A3",
    x"3E427950",
    x"3E4291FD",
    x"3E42AAAA",
    x"3E42C356",
    x"3E42DC03",
    x"3E42F4AF",
    x"3E430D5B",
    x"3E432607",
    x"3E433EB3",
    x"3E43575F",
    x"3E43700B",
    x"3E4388B7",
    x"3E43A162",
    x"3E43BA0E",
    x"3E43D2B9",
    x"3E43EB64",
    x"3E44040F",
    x"3E441CBA",
    x"3E443565",
    x"3E444E10",
    x"3E4466BA",
    x"3E447F65",
    x"3E44980F",
    x"3E44B0B9",
    x"3E44C963",
    x"3E44E20D",
    x"3E44FAB7",
    x"3E451361",
    x"3E452C0B",
    x"3E4544B4",
    x"3E455D5E",
    x"3E457607",
    x"3E458EB0",
    x"3E45A759",
    x"3E45C002",
    x"3E45D8AB",
    x"3E45F153",
    x"3E4609FC",
    x"3E4622A5",
    x"3E463B4D",
    x"3E4653F5",
    x"3E466C9D",
    x"3E468545",
    x"3E469DED",
    x"3E46B695",
    x"3E46CF3C",
    x"3E46E7E4",
    x"3E47008B",
    x"3E471932",
    x"3E4731DA",
    x"3E474A81",
    x"3E476328",
    x"3E477BCE",
    x"3E479475",
    x"3E47AD1B",
    x"3E47C5C2",
    x"3E47DE68",
    x"3E47F70E",
    x"3E480FB4",
    x"3E48285A",
    x"3E484100",
    x"3E4859A6",
    x"3E48724B",
    x"3E488AF1",
    x"3E48A396",
    x"3E48BC3B",
    x"3E48D4E0",
    x"3E48ED85",
    x"3E49062A",
    x"3E491ECF",
    x"3E493774",
    x"3E495018",
    x"3E4968BC",
    x"3E498161",
    x"3E499A05",
    x"3E49B2A9",
    x"3E49CB4D",
    x"3E49E3F0",
    x"3E49FC94",
    x"3E4A1538",
    x"3E4A2DDB",
    x"3E4A467E",
    x"3E4A5F21",
    x"3E4A77C4",
    x"3E4A9067",
    x"3E4AA90A",
    x"3E4AC1AD",
    x"3E4ADA4F",
    x"3E4AF2F2",
    x"3E4B0B94",
    x"3E4B2436",
    x"3E4B3CD8",
    x"3E4B557A",
    x"3E4B6E1C",
    x"3E4B86BE",
    x"3E4B9F5F",
    x"3E4BB801",
    x"3E4BD0A2",
    x"3E4BE943",
    x"3E4C01E4",
    x"3E4C1A85",
    x"3E4C3326",
    x"3E4C4BC7",
    x"3E4C6467",
    x"3E4C7D08",
    x"3E4C95A8",
    x"3E4CAE48",
    x"3E4CC6E8",
    x"3E4CDF88",
    x"3E4CF828",
    x"3E4D10C8",
    x"3E4D2967",
    x"3E4D4207",
    x"3E4D5AA6",
    x"3E4D7345",
    x"3E4D8BE4",
    x"3E4DA483",
    x"3E4DBD22",
    x"3E4DD5C1",
    x"3E4DEE60",
    x"3E4E06FE",
    x"3E4E1F9C",
    x"3E4E383B",
    x"3E4E50D9",
    x"3E4E6977",
    x"3E4E8215",
    x"3E4E9AB2",
    x"3E4EB350",
    x"3E4ECBED",
    x"3E4EE48B",
    x"3E4EFD28",
    x"3E4F15C5",
    x"3E4F2E62",
    x"3E4F46FF",
    x"3E4F5F9C",
    x"3E4F7838",
    x"3E4F90D5",
    x"3E4FA971",
    x"3E4FC20D",
    x"3E4FDAA9",
    x"3E4FF345",
    x"3E500BE1",
    x"3E50247D",
    x"3E503D19",
    x"3E5055B4",
    x"3E506E4F",
    x"3E5086EB",
    x"3E509F86",
    x"3E50B821",
    x"3E50D0BC",
    x"3E50E956",
    x"3E5101F1",
    x"3E511A8B",
    x"3E513326",
    x"3E514BC0",
    x"3E51645A",
    x"3E517CF4",
    x"3E51958E",
    x"3E51AE28",
    x"3E51C6C1",
    x"3E51DF5B",
    x"3E51F7F4",
    x"3E52108D",
    x"3E522926",
    x"3E5241BF",
    x"3E525A58",
    x"3E5272F1",
    x"3E528B89",
    x"3E52A422",
    x"3E52BCBA",
    x"3E52D552",
    x"3E52EDEA",
    x"3E530682",
    x"3E531F1A",
    x"3E5337B2",
    x"3E535049",
    x"3E5368E1",
    x"3E538178",
    x"3E539A0F",
    x"3E53B2A6",
    x"3E53CB3D",
    x"3E53E3D4",
    x"3E53FC6B",
    x"3E541501",
    x"3E542D98",
    x"3E54462E",
    x"3E545EC4",
    x"3E54775A",
    x"3E548FF0",
    x"3E54A886",
    x"3E54C11B",
    x"3E54D9B1",
    x"3E54F246",
    x"3E550ADC",
    x"3E552371",
    x"3E553C06",
    x"3E55549B",
    x"3E556D2F",
    x"3E5585C4",
    x"3E559E58",
    x"3E55B6ED",
    x"3E55CF81",
    x"3E55E815",
    x"3E5600A9",
    x"3E56193D",
    x"3E5631D1",
    x"3E564A64",
    x"3E5662F8",
    x"3E567B8B",
    x"3E56941E",
    x"3E56ACB1",
    x"3E56C544",
    x"3E56DDD7",
    x"3E56F66A",
    x"3E570EFC",
    x"3E57278F",
    x"3E574021",
    x"3E5758B3",
    x"3E577145",
    x"3E5789D7",
    x"3E57A269",
    x"3E57BAFB",
    x"3E57D38C",
    x"3E57EC1D",
    x"3E5804AF",
    x"3E581D40",
    x"3E5835D1",
    x"3E584E62",
    x"3E5866F2",
    x"3E587F83",
    x"3E589813",
    x"3E58B0A4",
    x"3E58C934",
    x"3E58E1C4",
    x"3E58FA54",
    x"3E5912E4",
    x"3E592B74",
    x"3E594403",
    x"3E595C93",
    x"3E597522",
    x"3E598DB1",
    x"3E59A640",
    x"3E59BECF",
    x"3E59D75E",
    x"3E59EFEC",
    x"3E5A087B",
    x"3E5A2109",
    x"3E5A3997",
    x"3E5A5226",
    x"3E5A6AB4",
    x"3E5A8341",
    x"3E5A9BCF",
    x"3E5AB45D",
    x"3E5ACCEA",
    x"3E5AE578",
    x"3E5AFE05",
    x"3E5B1692",
    x"3E5B2F1F",
    x"3E5B47AC",
    x"3E5B6038",
    x"3E5B78C5",
    x"3E5B9151",
    x"3E5BA9DD",
    x"3E5BC26A",
    x"3E5BDAF6",
    x"3E5BF381",
    x"3E5C0C0D",
    x"3E5C2499",
    x"3E5C3D24",
    x"3E5C55B0",
    x"3E5C6E3B",
    x"3E5C86C6",
    x"3E5C9F51",
    x"3E5CB7DC",
    x"3E5CD066",
    x"3E5CE8F1",
    x"3E5D017B",
    x"3E5D1A05",
    x"3E5D3290",
    x"3E5D4B1A",
    x"3E5D63A4",
    x"3E5D7C2D",
    x"3E5D94B7",
    x"3E5DAD40",
    x"3E5DC5CA",
    x"3E5DDE53",
    x"3E5DF6DC",
    x"3E5E0F65",
    x"3E5E27EE",
    x"3E5E4076",
    x"3E5E58FF",
    x"3E5E7187",
    x"3E5E8A10",
    x"3E5EA298",
    x"3E5EBB20",
    x"3E5ED3A8",
    x"3E5EEC2F",
    x"3E5F04B7",
    x"3E5F1D3E",
    x"3E5F35C6",
    x"3E5F4E4D",
    x"3E5F66D4",
    x"3E5F7F5B",
    x"3E5F97E2",
    x"3E5FB068",
    x"3E5FC8EF",
    x"3E5FE175",
    x"3E5FF9FC",
    x"3E601282",
    x"3E602B08",
    x"3E60438E",
    x"3E605C13",
    x"3E607499",
    x"3E608D1E",
    x"3E60A5A4",
    x"3E60BE29",
    x"3E60D6AE",
    x"3E60EF33",
    x"3E6107B8",
    x"3E61203C",
    x"3E6138C1",
    x"3E615145",
    x"3E6169C9",
    x"3E61824D",
    x"3E619AD1",
    x"3E61B355",
    x"3E61CBD9",
    x"3E61E45C",
    x"3E61FCE0",
    x"3E621563",
    x"3E622DE6",
    x"3E624669",
    x"3E625EEC",
    x"3E62776F",
    x"3E628FF1",
    x"3E62A874",
    x"3E62C0F6",
    x"3E62D978",
    x"3E62F1FA",
    x"3E630A7C",
    x"3E6322FE",
    x"3E633B80",
    x"3E635401",
    x"3E636C83",
    x"3E638504",
    x"3E639D85",
    x"3E63B606",
    x"3E63CE87",
    x"3E63E707",
    x"3E63FF88",
    x"3E641808",
    x"3E643089",
    x"3E644909",
    x"3E646189",
    x"3E647A09",
    x"3E649288",
    x"3E64AB08",
    x"3E64C387",
    x"3E64DC07",
    x"3E64F486",
    x"3E650D05",
    x"3E652584",
    x"3E653E02",
    x"3E655681",
    x"3E656F00",
    x"3E65877E",
    x"3E659FFC",
    x"3E65B87A",
    x"3E65D0F8",
    x"3E65E976",
    x"3E6601F3",
    x"3E661A71",
    x"3E6632EE",
    x"3E664B6C",
    x"3E6663E9",
    x"3E667C66",
    x"3E6694E2",
    x"3E66AD5F",
    x"3E66C5DC",
    x"3E66DE58",
    x"3E66F6D4",
    x"3E670F50",
    x"3E6727CC",
    x"3E674048",
    x"3E6758C4",
    x"3E67713F",
    x"3E6789BB",
    x"3E67A236",
    x"3E67BAB1",
    x"3E67D32C",
    x"3E67EBA7",
    x"3E680422",
    x"3E681C9C",
    x"3E683517",
    x"3E684D91",
    x"3E68660B",
    x"3E687E85",
    x"3E6896FF",
    x"3E68AF79",
    x"3E68C7F3",
    x"3E68E06C",
    x"3E68F8E5",
    x"3E69115F",
    x"3E6929D8",
    x"3E694251",
    x"3E695AC9",
    x"3E697342",
    x"3E698BBA",
    x"3E69A433",
    x"3E69BCAB",
    x"3E69D523",
    x"3E69ED9B",
    x"3E6A0613",
    x"3E6A1E8A",
    x"3E6A3702",
    x"3E6A4F79",
    x"3E6A67F0",
    x"3E6A8067",
    x"3E6A98DE",
    x"3E6AB155",
    x"3E6AC9CC",
    x"3E6AE242",
    x"3E6AFAB9",
    x"3E6B132F",
    x"3E6B2BA5",
    x"3E6B441B",
    x"3E6B5C91",
    x"3E6B7506",
    x"3E6B8D7C",
    x"3E6BA5F1",
    x"3E6BBE66",
    x"3E6BD6DC",
    x"3E6BEF51",
    x"3E6C07C5",
    x"3E6C203A",
    x"3E6C38AF",
    x"3E6C5123",
    x"3E6C6997",
    x"3E6C820B",
    x"3E6C9A7F",
    x"3E6CB2F3",
    x"3E6CCB67",
    x"3E6CE3DA",
    x"3E6CFC4E",
    x"3E6D14C1",
    x"3E6D2D34",
    x"3E6D45A7",
    x"3E6D5E1A",
    x"3E6D768C",
    x"3E6D8EFF",
    x"3E6DA771",
    x"3E6DBFE3",
    x"3E6DD856",
    x"3E6DF0C7",
    x"3E6E0939",
    x"3E6E21AB",
    x"3E6E3A1C",
    x"3E6E528E",
    x"3E6E6AFF",
    x"3E6E8370",
    x"3E6E9BE1",
    x"3E6EB452",
    x"3E6ECCC3",
    x"3E6EE533",
    x"3E6EFDA3",
    x"3E6F1614",
    x"3E6F2E84",
    x"3E6F46F4",
    x"3E6F5F63",
    x"3E6F77D3",
    x"3E6F9043",
    x"3E6FA8B2",
    x"3E6FC121",
    x"3E6FD990",
    x"3E6FF1FF",
    x"3E700A6E",
    x"3E7022DD",
    x"3E703B4B",
    x"3E7053B9",
    x"3E706C28",
    x"3E708496",
    x"3E709D04",
    x"3E70B571",
    x"3E70CDDF",
    x"3E70E64C",
    x"3E70FEBA",
    x"3E711727",
    x"3E712F94",
    x"3E714801",
    x"3E71606E",
    x"3E7178DA",
    x"3E719147",
    x"3E71A9B3",
    x"3E71C21F",
    x"3E71DA8B",
    x"3E71F2F7",
    x"3E720B63",
    x"3E7223CE",
    x"3E723C3A",
    x"3E7254A5",
    x"3E726D10",
    x"3E72857B",
    x"3E729DE6",
    x"3E72B651",
    x"3E72CEBC",
    x"3E72E726",
    x"3E72FF90",
    x"3E7317FA",
    x"3E733064",
    x"3E7348CE",
    x"3E736138",
    x"3E7379A1",
    x"3E73920B",
    x"3E73AA74",
    x"3E73C2DD",
    x"3E73DB46",
    x"3E73F3AF",
    x"3E740C18",
    x"3E742480",
    x"3E743CE8",
    x"3E745551",
    x"3E746DB9",
    x"3E748621",
    x"3E749E88",
    x"3E74B6F0",
    x"3E74CF57",
    x"3E74E7BF",
    x"3E750026",
    x"3E75188D",
    x"3E7530F4",
    x"3E75495B",
    x"3E7561C1",
    x"3E757A28",
    x"3E75928E",
    x"3E75AAF4",
    x"3E75C35A",
    x"3E75DBC0",
    x"3E75F426",
    x"3E760C8B",
    x"3E7624F1",
    x"3E763D56",
    x"3E7655BB",
    x"3E766E20",
    x"3E768685",
    x"3E769EEA",
    x"3E76B74E",
    x"3E76CFB2",
    x"3E76E817",
    x"3E77007B",
    x"3E7718DF",
    x"3E773142",
    x"3E7749A6",
    x"3E77620A",
    x"3E777A6D",
    x"3E7792D0",
    x"3E77AB33",
    x"3E77C396",
    x"3E77DBF9",
    x"3E77F45B",
    x"3E780CBE",
    x"3E782520",
    x"3E783D82",
    x"3E7855E4",
    x"3E786E46",
    x"3E7886A8",
    x"3E789F09",
    x"3E78B76B",
    x"3E78CFCC",
    x"3E78E82D",
    x"3E79008E",
    x"3E7918EF",
    x"3E79314F",
    x"3E7949B0",
    x"3E796210",
    x"3E797A70",
    x"3E7992D0",
    x"3E79AB30",
    x"3E79C390",
    x"3E79DBF0",
    x"3E79F44F",
    x"3E7A0CAE",
    x"3E7A250D",
    x"3E7A3D6C",
    x"3E7A55CB",
    x"3E7A6E2A",
    x"3E7A8688",
    x"3E7A9EE7",
    x"3E7AB745",
    x"3E7ACFA3",
    x"3E7AE801",
    x"3E7B005F",
    x"3E7B18BC",
    x"3E7B311A",
    x"3E7B4977",
    x"3E7B61D4",
    x"3E7B7A31",
    x"3E7B928E",
    x"3E7BAAEB",
    x"3E7BC348",
    x"3E7BDBA4",
    x"3E7BF400",
    x"3E7C0C5C",
    x"3E7C24B8",
    x"3E7C3D14",
    x"3E7C5570",
    x"3E7C6DCB",
    x"3E7C8627",
    x"3E7C9E82",
    x"3E7CB6DD",
    x"3E7CCF38",
    x"3E7CE793",
    x"3E7CFFED",
    x"3E7D1848",
    x"3E7D30A2",
    x"3E7D48FC",
    x"3E7D6156",
    x"3E7D79B0",
    x"3E7D9209",
    x"3E7DAA63",
    x"3E7DC2BC",
    x"3E7DDB16",
    x"3E7DF36F",
    x"3E7E0BC8",
    x"3E7E2420",
    x"3E7E3C79",
    x"3E7E54D1",
    x"3E7E6D2A",
    x"3E7E8582",
    x"3E7E9DDA",
    x"3E7EB632",
    x"3E7ECE89",
    x"3E7EE6E1",
    x"3E7EFF38",
    x"3E7F178F",
    x"3E7F2FE7",
    x"3E7F483D",
    x"3E7F6094",
    x"3E7F78EB",
    x"3E7F9141",
    x"3E7FA998",
    x"3E7FC1EE",
    x"3E7FDA44",
    x"3E7FF29A",
    x"3E800578",
    x"3E8011A2",
    x"3E801DCD",
    x"3E8029F8",
    x"3E803622",
    x"3E80424D",
    x"3E804E77",
    x"3E805AA1",
    x"3E8066CC",
    x"3E8072F6",
    x"3E807F20",
    x"3E808B4A",
    x"3E809774",
    x"3E80A39E",
    x"3E80AFC7",
    x"3E80BBF1",
    x"3E80C81B",
    x"3E80D444",
    x"3E80E06E",
    x"3E80EC97",
    x"3E80F8C0",
    x"3E8104E9",
    x"3E811113",
    x"3E811D3C",
    x"3E812965",
    x"3E81358E",
    x"3E8141B6",
    x"3E814DDF",
    x"3E815A08",
    x"3E816630",
    x"3E817259",
    x"3E817E81",
    x"3E818AAA",
    x"3E8196D2",
    x"3E81A2FA",
    x"3E81AF22",
    x"3E81BB4A",
    x"3E81C772",
    x"3E81D39A",
    x"3E81DFC2",
    x"3E81EBEA",
    x"3E81F811",
    x"3E820439",
    x"3E821060",
    x"3E821C88",
    x"3E8228AF",
    x"3E8234D7",
    x"3E8240FE",
    x"3E824D25",
    x"3E82594C",
    x"3E826573",
    x"3E82719A",
    x"3E827DC0",
    x"3E8289E7",
    x"3E82960E",
    x"3E82A234",
    x"3E82AE5B",
    x"3E82BA81",
    x"3E82C6A8",
    x"3E82D2CE",
    x"3E82DEF4",
    x"3E82EB1A",
    x"3E82F740",
    x"3E830366",
    x"3E830F8C",
    x"3E831BB2",
    x"3E8327D7",
    x"3E8333FD",
    x"3E834022",
    x"3E834C48",
    x"3E83586D",
    x"3E836493",
    x"3E8370B8",
    x"3E837CDD",
    x"3E838902",
    x"3E839527",
    x"3E83A14C",
    x"3E83AD71",
    x"3E83B995",
    x"3E83C5BA",
    x"3E83D1DF",
    x"3E83DE03",
    x"3E83EA28",
    x"3E83F64C",
    x"3E840270",
    x"3E840E94",
    x"3E841AB8",
    x"3E8426DD",
    x"3E843300",
    x"3E843F24",
    x"3E844B48",
    x"3E84576C",
    x"3E84638F",
    x"3E846FB3",
    x"3E847BD6",
    x"3E8487FA",
    x"3E84941D",
    x"3E84A040",
    x"3E84AC64",
    x"3E84B887",
    x"3E84C4AA",
    x"3E84D0CC",
    x"3E84DCEF",
    x"3E84E912",
    x"3E84F535",
    x"3E850157",
    x"3E850D7A",
    x"3E85199C",
    x"3E8525BF",
    x"3E8531E1",
    x"3E853E03",
    x"3E854A25",
    x"3E855647",
    x"3E856269",
    x"3E856E8B",
    x"3E857AAD",
    x"3E8586CE",
    x"3E8592F0",
    x"3E859F12",
    x"3E85AB33",
    x"3E85B755",
    x"3E85C376",
    x"3E85CF97",
    x"3E85DBB8",
    x"3E85E7D9",
    x"3E85F3FA",
    x"3E86001B",
    x"3E860C3C",
    x"3E86185D",
    x"3E86247D",
    x"3E86309E",
    x"3E863CBE",
    x"3E8648DF",
    x"3E8654FF",
    x"3E86611F",
    x"3E866D40",
    x"3E867960",
    x"3E868580",
    x"3E8691A0",
    x"3E869DBF",
    x"3E86A9DF",
    x"3E86B5FF",
    x"3E86C21F",
    x"3E86CE3E",
    x"3E86DA5D",
    x"3E86E67D",
    x"3E86F29C",
    x"3E86FEBB",
    x"3E870ADA",
    x"3E8716F9",
    x"3E872318",
    x"3E872F37",
    x"3E873B56",
    x"3E874775",
    x"3E875393",
    x"3E875FB2",
    x"3E876BD0",
    x"3E8777EF",
    x"3E87840D",
    x"3E87902B",
    x"3E879C49",
    x"3E87A868",
    x"3E87B486",
    x"3E87C0A3",
    x"3E87CCC1",
    x"3E87D8DF",
    x"3E87E4FD",
    x"3E87F11A",
    x"3E87FD38",
    x"3E880955",
    x"3E881572",
    x"3E882190",
    x"3E882DAD",
    x"3E8839CA",
    x"3E8845E7",
    x"3E885204",
    x"3E885E21",
    x"3E886A3D",
    x"3E88765A",
    x"3E888277",
    x"3E888E93",
    x"3E889AB0",
    x"3E88A6CC",
    x"3E88B2E8",
    x"3E88BF04",
    x"3E88CB20",
    x"3E88D73C",
    x"3E88E358",
    x"3E88EF74",
    x"3E88FB90",
    x"3E8907AC",
    x"3E8913C7",
    x"3E891FE3",
    x"3E892BFE",
    x"3E893819",
    x"3E894435",
    x"3E895050",
    x"3E895C6B",
    x"3E896886",
    x"3E8974A1",
    x"3E8980BC",
    x"3E898CD7",
    x"3E8998F1",
    x"3E89A50C",
    x"3E89B126",
    x"3E89BD41",
    x"3E89C95B",
    x"3E89D575",
    x"3E89E190",
    x"3E89EDAA",
    x"3E89F9C4",
    x"3E8A05DE",
    x"3E8A11F7",
    x"3E8A1E11",
    x"3E8A2A2B",
    x"3E8A3645",
    x"3E8A425E",
    x"3E8A4E78",
    x"3E8A5A91",
    x"3E8A66AA",
    x"3E8A72C3",
    x"3E8A7EDC",
    x"3E8A8AF5",
    x"3E8A970E",
    x"3E8AA327",
    x"3E8AAF40",
    x"3E8ABB59",
    x"3E8AC771",
    x"3E8AD38A",
    x"3E8ADFA2",
    x"3E8AEBBB",
    x"3E8AF7D3",
    x"3E8B03EB",
    x"3E8B1003",
    x"3E8B1C1B",
    x"3E8B2833",
    x"3E8B344B",
    x"3E8B4063",
    x"3E8B4C7A",
    x"3E8B5892",
    x"3E8B64AA",
    x"3E8B70C1",
    x"3E8B7CD8",
    x"3E8B88F0",
    x"3E8B9507",
    x"3E8BA11E",
    x"3E8BAD35",
    x"3E8BB94C",
    x"3E8BC563",
    x"3E8BD179",
    x"3E8BDD90",
    x"3E8BE9A7",
    x"3E8BF5BD",
    x"3E8C01D4",
    x"3E8C0DEA",
    x"3E8C1A00",
    x"3E8C2616",
    x"3E8C322C",
    x"3E8C3E42",
    x"3E8C4A58",
    x"3E8C566E",
    x"3E8C6284",
    x"3E8C6E9A",
    x"3E8C7AAF",
    x"3E8C86C5",
    x"3E8C92DA",
    x"3E8C9EEF",
    x"3E8CAB05",
    x"3E8CB71A",
    x"3E8CC32F",
    x"3E8CCF44",
    x"3E8CDB59",
    x"3E8CE76D",
    x"3E8CF382",
    x"3E8CFF97",
    x"3E8D0BAB",
    x"3E8D17C0",
    x"3E8D23D4",
    x"3E8D2FE9",
    x"3E8D3BFD",
    x"3E8D4811",
    x"3E8D5425",
    x"3E8D6039",
    x"3E8D6C4D",
    x"3E8D7861",
    x"3E8D8474",
    x"3E8D9088",
    x"3E8D9C9B",
    x"3E8DA8AF",
    x"3E8DB4C2",
    x"3E8DC0D6",
    x"3E8DCCE9",
    x"3E8DD8FC",
    x"3E8DE50F",
    x"3E8DF122",
    x"3E8DFD35",
    x"3E8E0947",
    x"3E8E155A",
    x"3E8E216D",
    x"3E8E2D7F",
    x"3E8E3992",
    x"3E8E45A4",
    x"3E8E51B6",
    x"3E8E5DC8",
    x"3E8E69DB",
    x"3E8E75ED",
    x"3E8E81FE",
    x"3E8E8E10",
    x"3E8E9A22",
    x"3E8EA634",
    x"3E8EB245",
    x"3E8EBE57",
    x"3E8ECA68",
    x"3E8ED679",
    x"3E8EE28B",
    x"3E8EEE9C",
    x"3E8EFAAD",
    x"3E8F06BE",
    x"3E8F12CF",
    x"3E8F1EDF",
    x"3E8F2AF0",
    x"3E8F3701",
    x"3E8F4311",
    x"3E8F4F22",
    x"3E8F5B32",
    x"3E8F6742",
    x"3E8F7353",
    x"3E8F7F63",
    x"3E8F8B73",
    x"3E8F9783",
    x"3E8FA392",
    x"3E8FAFA2",
    x"3E8FBBB2",
    x"3E8FC7C1",
    x"3E8FD3D1",
    x"3E8FDFE0",
    x"3E8FEBF0",
    x"3E8FF7FF",
    x"3E90040E",
    x"3E90101D",
    x"3E901C2C",
    x"3E90283B",
    x"3E90344A",
    x"3E904059",
    x"3E904C67",
    x"3E905876",
    x"3E906484",
    x"3E907093",
    x"3E907CA1",
    x"3E9088AF",
    x"3E9094BD",
    x"3E90A0CB",
    x"3E90ACD9",
    x"3E90B8E7",
    x"3E90C4F5",
    x"3E90D102",
    x"3E90DD10",
    x"3E90E91D",
    x"3E90F52B",
    x"3E910138",
    x"3E910D45",
    x"3E911953",
    x"3E912560",
    x"3E91316D",
    x"3E913D79",
    x"3E914986",
    x"3E915593",
    x"3E9161A0",
    x"3E916DAC",
    x"3E9179B9",
    x"3E9185C5",
    x"3E9191D1",
    x"3E919DDD",
    x"3E91A9E9",
    x"3E91B5F5",
    x"3E91C201",
    x"3E91CE0D",
    x"3E91DA19",
    x"3E91E625",
    x"3E91F230",
    x"3E91FE3C",
    x"3E920A47",
    x"3E921652",
    x"3E92225E",
    x"3E922E69",
    x"3E923A74",
    x"3E92467F",
    x"3E92528A",
    x"3E925E94",
    x"3E926A9F",
    x"3E9276AA",
    x"3E9282B4",
    x"3E928EBF",
    x"3E929AC9",
    x"3E92A6D3",
    x"3E92B2DD",
    x"3E92BEE7",
    x"3E92CAF1",
    x"3E92D6FB",
    x"3E92E305",
    x"3E92EF0F",
    x"3E92FB18",
    x"3E930722",
    x"3E93132B",
    x"3E931F35",
    x"3E932B3E",
    x"3E933747",
    x"3E934350",
    x"3E934F59",
    x"3E935B62",
    x"3E93676B",
    x"3E937374",
    x"3E937F7D",
    x"3E938B85",
    x"3E93978E",
    x"3E93A396",
    x"3E93AF9E",
    x"3E93BBA6",
    x"3E93C7AF",
    x"3E93D3B7",
    x"3E93DFBF",
    x"3E93EBC6",
    x"3E93F7CE",
    x"3E9403D6",
    x"3E940FDD",
    x"3E941BE5",
    x"3E9427EC",
    x"3E9433F4",
    x"3E943FFB",
    x"3E944C02",
    x"3E945809",
    x"3E946410",
    x"3E947017",
    x"3E947C1E",
    x"3E948824",
    x"3E94942B",
    x"3E94A031",
    x"3E94AC38",
    x"3E94B83E",
    x"3E94C444",
    x"3E94D04B",
    x"3E94DC51",
    x"3E94E857",
    x"3E94F45D",
    x"3E950062",
    x"3E950C68",
    x"3E95186E",
    x"3E952473",
    x"3E953079",
    x"3E953C7E",
    x"3E954883",
    x"3E955488",
    x"3E95608D",
    x"3E956C92",
    x"3E957897",
    x"3E95849C",
    x"3E9590A1",
    x"3E959CA6",
    x"3E95A8AA",
    x"3E95B4AE",
    x"3E95C0B3",
    x"3E95CCB7",
    x"3E95D8BB",
    x"3E95E4BF",
    x"3E95F0C3",
    x"3E95FCC7",
    x"3E9608CB",
    x"3E9614CF",
    x"3E9620D2",
    x"3E962CD6",
    x"3E9638D9",
    x"3E9644DD",
    x"3E9650E0",
    x"3E965CE3",
    x"3E9668E6",
    x"3E9674E9",
    x"3E9680EC",
    x"3E968CEF",
    x"3E9698F2",
    x"3E96A4F4",
    x"3E96B0F7",
    x"3E96BCF9",
    x"3E96C8FC",
    x"3E96D4FE",
    x"3E96E100",
    x"3E96ED02",
    x"3E96F904",
    x"3E970506",
    x"3E971108",
    x"3E971D0A",
    x"3E97290B",
    x"3E97350D",
    x"3E97410E",
    x"3E974D10",
    x"3E975911",
    x"3E976512",
    x"3E977113",
    x"3E977D14",
    x"3E978915",
    x"3E979516",
    x"3E97A117",
    x"3E97AD17",
    x"3E97B918",
    x"3E97C518",
    x"3E97D119",
    x"3E97DD19",
    x"3E97E919",
    x"3E97F519",
    x"3E980119",
    x"3E980D19",
    x"3E981919",
    x"3E982519",
    x"3E983118",
    x"3E983D18",
    x"3E984917",
    x"3E985517",
    x"3E986116",
    x"3E986D15",
    x"3E987914",
    x"3E988513",
    x"3E989112",
    x"3E989D11",
    x"3E98A910",
    x"3E98B50E",
    x"3E98C10D",
    x"3E98CD0B",
    x"3E98D90A",
    x"3E98E508",
    x"3E98F106",
    x"3E98FD04",
    x"3E990902",
    x"3E991500",
    x"3E9920FE",
    x"3E992CFB",
    x"3E9938F9",
    x"3E9944F7",
    x"3E9950F4",
    x"3E995CF1",
    x"3E9968EE",
    x"3E9974EC",
    x"3E9980E9",
    x"3E998CE6",
    x"3E9998E3",
    x"3E99A4DF",
    x"3E99B0DC",
    x"3E99BCD9",
    x"3E99C8D5",
    x"3E99D4D1",
    x"3E99E0CE",
    x"3E99ECCA",
    x"3E99F8C6",
    x"3E9A04C2",
    x"3E9A10BE",
    x"3E9A1CBA",
    x"3E9A28B6",
    x"3E9A34B1",
    x"3E9A40AD",
    x"3E9A4CA8",
    x"3E9A58A4",
    x"3E9A649F",
    x"3E9A709A",
    x"3E9A7C95",
    x"3E9A8890",
    x"3E9A948B",
    x"3E9AA086",
    x"3E9AAC81",
    x"3E9AB87B",
    x"3E9AC476",
    x"3E9AD070",
    x"3E9ADC6B",
    x"3E9AE865",
    x"3E9AF45F",
    x"3E9B0059",
    x"3E9B0C53",
    x"3E9B184D",
    x"3E9B2447",
    x"3E9B3041",
    x"3E9B3C3A",
    x"3E9B4834",
    x"3E9B542D",
    x"3E9B6027",
    x"3E9B6C20",
    x"3E9B7819",
    x"3E9B8412",
    x"3E9B900B",
    x"3E9B9C04",
    x"3E9BA7FD",
    x"3E9BB3F5",
    x"3E9BBFEE",
    x"3E9BCBE6",
    x"3E9BD7DF",
    x"3E9BE3D7",
    x"3E9BEFCF",
    x"3E9BFBC7",
    x"3E9C07BF",
    x"3E9C13B7",
    x"3E9C1FAF",
    x"3E9C2BA7",
    x"3E9C379E",
    x"3E9C4396",
    x"3E9C4F8D",
    x"3E9C5B85",
    x"3E9C677C",
    x"3E9C7373",
    x"3E9C7F6A",
    x"3E9C8B61",
    x"3E9C9758",
    x"3E9CA34F",
    x"3E9CAF46",
    x"3E9CBB3C",
    x"3E9CC733",
    x"3E9CD329",
    x"3E9CDF20",
    x"3E9CEB16",
    x"3E9CF70C",
    x"3E9D0302",
    x"3E9D0EF8",
    x"3E9D1AEE",
    x"3E9D26E3",
    x"3E9D32D9",
    x"3E9D3ECF",
    x"3E9D4AC4",
    x"3E9D56BA",
    x"3E9D62AF",
    x"3E9D6EA4",
    x"3E9D7A99",
    x"3E9D868E",
    x"3E9D9283",
    x"3E9D9E78",
    x"3E9DAA6D",
    x"3E9DB661",
    x"3E9DC256",
    x"3E9DCE4A",
    x"3E9DDA3E",
    x"3E9DE633",
    x"3E9DF227",
    x"3E9DFE1B",
    x"3E9E0A0F",
    x"3E9E1603",
    x"3E9E21F6",
    x"3E9E2DEA",
    x"3E9E39DE",
    x"3E9E45D1",
    x"3E9E51C4",
    x"3E9E5DB8",
    x"3E9E69AB",
    x"3E9E759E",
    x"3E9E8191",
    x"3E9E8D84",
    x"3E9E9977",
    x"3E9EA569",
    x"3E9EB15C",
    x"3E9EBD4F",
    x"3E9EC941",
    x"3E9ED533",
    x"3E9EE126",
    x"3E9EED18",
    x"3E9EF90A",
    x"3E9F04FC",
    x"3E9F10EE",
    x"3E9F1CDF",
    x"3E9F28D1",
    x"3E9F34C3",
    x"3E9F40B4",
    x"3E9F4CA5",
    x"3E9F5897",
    x"3E9F6488",
    x"3E9F7079",
    x"3E9F7C6A",
    x"3E9F885B",
    x"3E9F944C",
    x"3E9FA03C",
    x"3E9FAC2D",
    x"3E9FB81D",
    x"3E9FC40E",
    x"3E9FCFFE",
    x"3E9FDBEE",
    x"3E9FE7DE",
    x"3E9FF3CE",
    x"3E9FFFBE",
    x"3EA00BAE",
    x"3EA0179E",
    x"3EA0238E",
    x"3EA02F7D",
    x"3EA03B6D",
    x"3EA0475C",
    x"3EA0534B",
    x"3EA05F3A",
    x"3EA06B29",
    x"3EA07718",
    x"3EA08307",
    x"3EA08EF6",
    x"3EA09AE5",
    x"3EA0A6D3",
    x"3EA0B2C2",
    x"3EA0BEB0",
    x"3EA0CA9E",
    x"3EA0D68D",
    x"3EA0E27B",
    x"3EA0EE69",
    x"3EA0FA57",
    x"3EA10644",
    x"3EA11232",
    x"3EA11E20",
    x"3EA12A0D",
    x"3EA135FB",
    x"3EA141E8",
    x"3EA14DD5",
    x"3EA159C2",
    x"3EA165AF",
    x"3EA1719C",
    x"3EA17D89",
    x"3EA18976",
    x"3EA19562",
    x"3EA1A14F",
    x"3EA1AD3B",
    x"3EA1B928",
    x"3EA1C514",
    x"3EA1D100",
    x"3EA1DCEC",
    x"3EA1E8D8",
    x"3EA1F4C4",
    x"3EA200B0",
    x"3EA20C9B",
    x"3EA21887",
    x"3EA22472",
    x"3EA2305E",
    x"3EA23C49",
    x"3EA24834",
    x"3EA2541F",
    x"3EA2600A",
    x"3EA26BF5",
    x"3EA277E0",
    x"3EA283CB",
    x"3EA28FB5",
    x"3EA29BA0",
    x"3EA2A78A",
    x"3EA2B374",
    x"3EA2BF5E",
    x"3EA2CB49",
    x"3EA2D733",
    x"3EA2E31C",
    x"3EA2EF06",
    x"3EA2FAF0",
    x"3EA306DA",
    x"3EA312C3",
    x"3EA31EAD",
    x"3EA32A96",
    x"3EA3367F",
    x"3EA34268",
    x"3EA34E51",
    x"3EA35A3A",
    x"3EA36623",
    x"3EA3720C",
    x"3EA37DF4",
    x"3EA389DD",
    x"3EA395C5",
    x"3EA3A1AD",
    x"3EA3AD96",
    x"3EA3B97E",
    x"3EA3C566",
    x"3EA3D14E",
    x"3EA3DD36",
    x"3EA3E91D",
    x"3EA3F505",
    x"3EA400ED",
    x"3EA40CD4",
    x"3EA418BB",
    x"3EA424A3",
    x"3EA4308A",
    x"3EA43C71",
    x"3EA44858",
    x"3EA4543F",
    x"3EA46025",
    x"3EA46C0C",
    x"3EA477F2",
    x"3EA483D9",
    x"3EA48FBF",
    x"3EA49BA6",
    x"3EA4A78C",
    x"3EA4B372",
    x"3EA4BF58",
    x"3EA4CB3E",
    x"3EA4D723",
    x"3EA4E309",
    x"3EA4EEEE",
    x"3EA4FAD4",
    x"3EA506B9",
    x"3EA5129F",
    x"3EA51E84",
    x"3EA52A69",
    x"3EA5364E",
    x"3EA54233",
    x"3EA54E17",
    x"3EA559FC",
    x"3EA565E1",
    x"3EA571C5",
    x"3EA57DA9",
    x"3EA5898E",
    x"3EA59572",
    x"3EA5A156",
    x"3EA5AD3A",
    x"3EA5B91E",
    x"3EA5C501",
    x"3EA5D0E5",
    x"3EA5DCC9",
    x"3EA5E8AC",
    x"3EA5F48F",
    x"3EA60073",
    x"3EA60C56",
    x"3EA61839",
    x"3EA6241C",
    x"3EA62FFF",
    x"3EA63BE2",
    x"3EA647C4",
    x"3EA653A7",
    x"3EA65F89",
    x"3EA66B6C",
    x"3EA6774E",
    x"3EA68330",
    x"3EA68F12",
    x"3EA69AF4",
    x"3EA6A6D6",
    x"3EA6B2B8",
    x"3EA6BE99",
    x"3EA6CA7B",
    x"3EA6D65C",
    x"3EA6E23E",
    x"3EA6EE1F",
    x"3EA6FA00",
    x"3EA705E1",
    x"3EA711C2",
    x"3EA71DA3",
    x"3EA72984",
    x"3EA73564",
    x"3EA74145",
    x"3EA74D25",
    x"3EA75906",
    x"3EA764E6",
    x"3EA770C6",
    x"3EA77CA6",
    x"3EA78886",
    x"3EA79466",
    x"3EA7A046",
    x"3EA7AC25",
    x"3EA7B805",
    x"3EA7C3E4",
    x"3EA7CFC4",
    x"3EA7DBA3",
    x"3EA7E782",
    x"3EA7F361",
    x"3EA7FF40",
    x"3EA80B1F",
    x"3EA816FE",
    x"3EA822DC",
    x"3EA82EBB",
    x"3EA83A99",
    x"3EA84678",
    x"3EA85256",
    x"3EA85E34",
    x"3EA86A12",
    x"3EA875F0",
    x"3EA881CE",
    x"3EA88DAB",
    x"3EA89989",
    x"3EA8A567",
    x"3EA8B144",
    x"3EA8BD21",
    x"3EA8C8FE",
    x"3EA8D4DC",
    x"3EA8E0B9",
    x"3EA8EC95",
    x"3EA8F872",
    x"3EA9044F",
    x"3EA9102C",
    x"3EA91C08",
    x"3EA927E5",
    x"3EA933C1",
    x"3EA93F9D",
    x"3EA94B79",
    x"3EA95755",
    x"3EA96331",
    x"3EA96F0D",
    x"3EA97AE8",
    x"3EA986C4",
    x"3EA992A0",
    x"3EA99E7B",
    x"3EA9AA56",
    x"3EA9B631",
    x"3EA9C20C",
    x"3EA9CDE7",
    x"3EA9D9C2",
    x"3EA9E59D",
    x"3EA9F178",
    x"3EA9FD52",
    x"3EAA092D",
    x"3EAA1507",
    x"3EAA20E1",
    x"3EAA2CBB",
    x"3EAA3895",
    x"3EAA446F",
    x"3EAA5049",
    x"3EAA5C23",
    x"3EAA67FD",
    x"3EAA73D6",
    x"3EAA7FB0",
    x"3EAA8B89",
    x"3EAA9762",
    x"3EAAA33B",
    x"3EAAAF14",
    x"3EAABAED",
    x"3EAAC6C6",
    x"3EAAD29F",
    x"3EAADE77",
    x"3EAAEA50",
    x"3EAAF628",
    x"3EAB0201",
    x"3EAB0DD9",
    x"3EAB19B1",
    x"3EAB2589",
    x"3EAB3161",
    x"3EAB3D39",
    x"3EAB4910",
    x"3EAB54E8",
    x"3EAB60BF",
    x"3EAB6C97",
    x"3EAB786E",
    x"3EAB8445",
    x"3EAB901C",
    x"3EAB9BF3",
    x"3EABA7CA",
    x"3EABB3A1",
    x"3EABBF77",
    x"3EABCB4E",
    x"3EABD724",
    x"3EABE2FB",
    x"3EABEED1",
    x"3EABFAA7",
    x"3EAC067D",
    x"3EAC1253",
    x"3EAC1E29",
    x"3EAC29FF",
    x"3EAC35D4",
    x"3EAC41AA",
    x"3EAC4D7F",
    x"3EAC5954",
    x"3EAC652A",
    x"3EAC70FF",
    x"3EAC7CD4",
    x"3EAC88A9",
    x"3EAC947D",
    x"3EACA052",
    x"3EACAC27",
    x"3EACB7FB",
    x"3EACC3CF",
    x"3EACCFA4",
    x"3EACDB78",
    x"3EACE74C",
    x"3EACF320",
    x"3EACFEF4",
    x"3EAD0AC7",
    x"3EAD169B",
    x"3EAD226F",
    x"3EAD2E42",
    x"3EAD3A15",
    x"3EAD45E9",
    x"3EAD51BC",
    x"3EAD5D8F",
    x"3EAD6962",
    x"3EAD7534",
    x"3EAD8107",
    x"3EAD8CDA",
    x"3EAD98AC",
    x"3EADA47F",
    x"3EADB051",
    x"3EADBC23",
    x"3EADC7F5",
    x"3EADD3C7",
    x"3EADDF99",
    x"3EADEB6B",
    x"3EADF73C",
    x"3EAE030E",
    x"3EAE0EDF",
    x"3EAE1AB1",
    x"3EAE2682",
    x"3EAE3253",
    x"3EAE3E24",
    x"3EAE49F5",
    x"3EAE55C6",
    x"3EAE6197",
    x"3EAE6D67",
    x"3EAE7938",
    x"3EAE8508",
    x"3EAE90D8",
    x"3EAE9CA8",
    x"3EAEA879",
    x"3EAEB449",
    x"3EAEC018",
    x"3EAECBE8",
    x"3EAED7B8",
    x"3EAEE387",
    x"3EAEEF57",
    x"3EAEFB26",
    x"3EAF06F5",
    x"3EAF12C5",
    x"3EAF1E94",
    x"3EAF2A62",
    x"3EAF3631",
    x"3EAF4200",
    x"3EAF4DCF",
    x"3EAF599D",
    x"3EAF656B",
    x"3EAF713A",
    x"3EAF7D08",
    x"3EAF88D6",
    x"3EAF94A4",
    x"3EAFA072",
    x"3EAFAC40",
    x"3EAFB80D",
    x"3EAFC3DB",
    x"3EAFCFA8",
    x"3EAFDB76",
    x"3EAFE743",
    x"3EAFF310",
    x"3EAFFEDD",
    x"3EB00AAA",
    x"3EB01677",
    x"3EB02243",
    x"3EB02E10",
    x"3EB039DC",
    x"3EB045A9",
    x"3EB05175",
    x"3EB05D41",
    x"3EB0690D",
    x"3EB074D9",
    x"3EB080A5",
    x"3EB08C71",
    x"3EB0983C",
    x"3EB0A408",
    x"3EB0AFD3",
    x"3EB0BB9F",
    x"3EB0C76A",
    x"3EB0D335",
    x"3EB0DF00",
    x"3EB0EACB",
    x"3EB0F696",
    x"3EB10260",
    x"3EB10E2B",
    x"3EB119F5",
    x"3EB125C0",
    x"3EB1318A",
    x"3EB13D54",
    x"3EB1491E",
    x"3EB154E8",
    x"3EB160B2",
    x"3EB16C7C",
    x"3EB17845",
    x"3EB1840F",
    x"3EB18FD8",
    x"3EB19BA1",
    x"3EB1A76B",
    x"3EB1B334",
    x"3EB1BEFD",
    x"3EB1CAC5",
    x"3EB1D68E",
    x"3EB1E257",
    x"3EB1EE1F",
    x"3EB1F9E8",
    x"3EB205B0",
    x"3EB21178",
    x"3EB21D41",
    x"3EB22909",
    x"3EB234D0",
    x"3EB24098",
    x"3EB24C60",
    x"3EB25827",
    x"3EB263EF",
    x"3EB26FB6",
    x"3EB27B7E",
    x"3EB28745",
    x"3EB2930C",
    x"3EB29ED3",
    x"3EB2AA99",
    x"3EB2B660",
    x"3EB2C227",
    x"3EB2CDED",
    x"3EB2D9B4",
    x"3EB2E57A",
    x"3EB2F140",
    x"3EB2FD06",
    x"3EB308CC",
    x"3EB31492",
    x"3EB32058",
    x"3EB32C1D",
    x"3EB337E3",
    x"3EB343A8",
    x"3EB34F6E",
    x"3EB35B33",
    x"3EB366F8",
    x"3EB372BD",
    x"3EB37E82",
    x"3EB38A47",
    x"3EB3960B",
    x"3EB3A1D0",
    x"3EB3AD94",
    x"3EB3B959",
    x"3EB3C51D",
    x"3EB3D0E1",
    x"3EB3DCA5",
    x"3EB3E869",
    x"3EB3F42D",
    x"3EB3FFF0",
    x"3EB40BB4",
    x"3EB41777",
    x"3EB4233B",
    x"3EB42EFE",
    x"3EB43AC1",
    x"3EB44684",
    x"3EB45247",
    x"3EB45E0A",
    x"3EB469CD",
    x"3EB4758F",
    x"3EB48152",
    x"3EB48D14",
    x"3EB498D6",
    x"3EB4A499",
    x"3EB4B05B",
    x"3EB4BC1D",
    x"3EB4C7DE",
    x"3EB4D3A0",
    x"3EB4DF62",
    x"3EB4EB23",
    x"3EB4F6E5",
    x"3EB502A6",
    x"3EB50E67",
    x"3EB51A28",
    x"3EB525E9",
    x"3EB531AA",
    x"3EB53D6B",
    x"3EB5492B",
    x"3EB554EC",
    x"3EB560AC",
    x"3EB56C6D",
    x"3EB5782D",
    x"3EB583ED",
    x"3EB58FAD",
    x"3EB59B6D",
    x"3EB5A72D",
    x"3EB5B2EC",
    x"3EB5BEAC",
    x"3EB5CA6B",
    x"3EB5D62B",
    x"3EB5E1EA",
    x"3EB5EDA9",
    x"3EB5F968",
    x"3EB60527",
    x"3EB610E6",
    x"3EB61CA4",
    x"3EB62863",
    x"3EB63421",
    x"3EB63FE0",
    x"3EB64B9E",
    x"3EB6575C",
    x"3EB6631A",
    x"3EB66ED8",
    x"3EB67A96",
    x"3EB68653",
    x"3EB69211",
    x"3EB69DCE",
    x"3EB6A98C",
    x"3EB6B549",
    x"3EB6C106",
    x"3EB6CCC3",
    x"3EB6D880",
    x"3EB6E43D",
    x"3EB6EFFA",
    x"3EB6FBB6",
    x"3EB70773",
    x"3EB7132F",
    x"3EB71EEB",
    x"3EB72AA7",
    x"3EB73663",
    x"3EB7421F",
    x"3EB74DDB",
    x"3EB75997",
    x"3EB76552",
    x"3EB7710E",
    x"3EB77CC9",
    x"3EB78884",
    x"3EB79440",
    x"3EB79FFB",
    x"3EB7ABB6",
    x"3EB7B770",
    x"3EB7C32B",
    x"3EB7CEE6",
    x"3EB7DAA0",
    x"3EB7E65B",
    x"3EB7F215",
    x"3EB7FDCF",
    x"3EB80989",
    x"3EB81543",
    x"3EB820FD",
    x"3EB82CB6",
    x"3EB83870",
    x"3EB8442A",
    x"3EB84FE3",
    x"3EB85B9C",
    x"3EB86755",
    x"3EB8730E",
    x"3EB87EC7",
    x"3EB88A80",
    x"3EB89639",
    x"3EB8A1F1",
    x"3EB8ADAA",
    x"3EB8B962",
    x"3EB8C51B",
    x"3EB8D0D3",
    x"3EB8DC8B",
    x"3EB8E843",
    x"3EB8F3FA",
    x"3EB8FFB2",
    x"3EB90B6A",
    x"3EB91721",
    x"3EB922D9",
    x"3EB92E90",
    x"3EB93A47",
    x"3EB945FE",
    x"3EB951B5",
    x"3EB95D6C",
    x"3EB96923",
    x"3EB974D9",
    x"3EB98090",
    x"3EB98C46",
    x"3EB997FC",
    x"3EB9A3B2",
    x"3EB9AF68",
    x"3EB9BB1E",
    x"3EB9C6D4",
    x"3EB9D28A",
    x"3EB9DE3F",
    x"3EB9E9F5",
    x"3EB9F5AA",
    x"3EBA015F",
    x"3EBA0D15",
    x"3EBA18CA",
    x"3EBA247F",
    x"3EBA3033",
    x"3EBA3BE8",
    x"3EBA479D",
    x"3EBA5351",
    x"3EBA5F05",
    x"3EBA6ABA",
    x"3EBA766E",
    x"3EBA8222",
    x"3EBA8DD6",
    x"3EBA9989",
    x"3EBAA53D",
    x"3EBAB0F1",
    x"3EBABCA4",
    x"3EBAC857",
    x"3EBAD40B",
    x"3EBADFBE",
    x"3EBAEB71",
    x"3EBAF724",
    x"3EBB02D6",
    x"3EBB0E89",
    x"3EBB1A3C",
    x"3EBB25EE",
    x"3EBB31A0",
    x"3EBB3D53",
    x"3EBB4905",
    x"3EBB54B7",
    x"3EBB6069",
    x"3EBB6C1A",
    x"3EBB77CC",
    x"3EBB837E",
    x"3EBB8F2F",
    x"3EBB9AE0",
    x"3EBBA692",
    x"3EBBB243",
    x"3EBBBDF4",
    x"3EBBC9A4",
    x"3EBBD555",
    x"3EBBE106",
    x"3EBBECB6",
    x"3EBBF867",
    x"3EBC0417",
    x"3EBC0FC7",
    x"3EBC1B77",
    x"3EBC2727",
    x"3EBC32D7",
    x"3EBC3E87",
    x"3EBC4A36",
    x"3EBC55E6",
    x"3EBC6195",
    x"3EBC6D45",
    x"3EBC78F4",
    x"3EBC84A3",
    x"3EBC9052",
    x"3EBC9C00",
    x"3EBCA7AF",
    x"3EBCB35E",
    x"3EBCBF0C",
    x"3EBCCABB",
    x"3EBCD669",
    x"3EBCE217",
    x"3EBCEDC5",
    x"3EBCF973",
    x"3EBD0521",
    x"3EBD10CE",
    x"3EBD1C7C",
    x"3EBD2829",
    x"3EBD33D7",
    x"3EBD3F84",
    x"3EBD4B31",
    x"3EBD56DE",
    x"3EBD628B",
    x"3EBD6E38",
    x"3EBD79E4",
    x"3EBD8591",
    x"3EBD913D",
    x"3EBD9CEA",
    x"3EBDA896",
    x"3EBDB442",
    x"3EBDBFEE",
    x"3EBDCB9A",
    x"3EBDD746",
    x"3EBDE2F1",
    x"3EBDEE9D",
    x"3EBDFA48",
    x"3EBE05F3",
    x"3EBE119E",
    x"3EBE1D4A",
    x"3EBE28F4",
    x"3EBE349F",
    x"3EBE404A",
    x"3EBE4BF5",
    x"3EBE579F",
    x"3EBE6349",
    x"3EBE6EF4",
    x"3EBE7A9E",
    x"3EBE8648",
    x"3EBE91F2",
    x"3EBE9D9C",
    x"3EBEA945",
    x"3EBEB4EF",
    x"3EBEC098",
    x"3EBECC42",
    x"3EBED7EB",
    x"3EBEE394",
    x"3EBEEF3D",
    x"3EBEFAE6",
    x"3EBF068F",
    x"3EBF1237",
    x"3EBF1DE0",
    x"3EBF2988",
    x"3EBF3530",
    x"3EBF40D9",
    x"3EBF4C81",
    x"3EBF5829",
    x"3EBF63D0",
    x"3EBF6F78",
    x"3EBF7B20",
    x"3EBF86C7",
    x"3EBF926F",
    x"3EBF9E16",
    x"3EBFA9BD",
    x"3EBFB564",
    x"3EBFC10B",
    x"3EBFCCB2",
    x"3EBFD858",
    x"3EBFE3FF",
    x"3EBFEFA5",
    x"3EBFFB4C",
    x"3EC006F2",
    x"3EC01298",
    x"3EC01E3E",
    x"3EC029E4",
    x"3EC0358A",
    x"3EC0412F",
    x"3EC04CD5",
    x"3EC0587A",
    x"3EC06420",
    x"3EC06FC5",
    x"3EC07B6A",
    x"3EC0870F",
    x"3EC092B4",
    x"3EC09E58",
    x"3EC0A9FD",
    x"3EC0B5A1",
    x"3EC0C146",
    x"3EC0CCEA",
    x"3EC0D88E",
    x"3EC0E432",
    x"3EC0EFD6",
    x"3EC0FB7A",
    x"3EC1071E",
    x"3EC112C1",
    x"3EC11E64",
    x"3EC12A08",
    x"3EC135AB",
    x"3EC1414E",
    x"3EC14CF1",
    x"3EC15894",
    x"3EC16437",
    x"3EC16FD9",
    x"3EC17B7C",
    x"3EC1871E",
    x"3EC192C0",
    x"3EC19E63",
    x"3EC1AA05",
    x"3EC1B5A7",
    x"3EC1C148",
    x"3EC1CCEA",
    x"3EC1D88C",
    x"3EC1E42D",
    x"3EC1EFCE",
    x"3EC1FB70",
    x"3EC20711",
    x"3EC212B2",
    x"3EC21E53",
    x"3EC229F3",
    x"3EC23594",
    x"3EC24135",
    x"3EC24CD5",
    x"3EC25875",
    x"3EC26415",
    x"3EC26FB5",
    x"3EC27B55",
    x"3EC286F5",
    x"3EC29295",
    x"3EC29E34",
    x"3EC2A9D4",
    x"3EC2B573",
    x"3EC2C112",
    x"3EC2CCB2",
    x"3EC2D851",
    x"3EC2E3EF",
    x"3EC2EF8E",
    x"3EC2FB2D",
    x"3EC306CB",
    x"3EC3126A",
    x"3EC31E08",
    x"3EC329A6",
    x"3EC33544",
    x"3EC340E2",
    x"3EC34C80",
    x"3EC3581E",
    x"3EC363BB",
    x"3EC36F59",
    x"3EC37AF6",
    x"3EC38693",
    x"3EC39231",
    x"3EC39DCE",
    x"3EC3A96A",
    x"3EC3B507",
    x"3EC3C0A4",
    x"3EC3CC40",
    x"3EC3D7DD",
    x"3EC3E379",
    x"3EC3EF15",
    x"3EC3FAB1",
    x"3EC4064D",
    x"3EC411E9",
    x"3EC41D85",
    x"3EC42920",
    x"3EC434BC",
    x"3EC44057",
    x"3EC44BF2",
    x"3EC4578D",
    x"3EC46328",
    x"3EC46EC3",
    x"3EC47A5E",
    x"3EC485F9",
    x"3EC49193",
    x"3EC49D2E",
    x"3EC4A8C8",
    x"3EC4B462",
    x"3EC4BFFC",
    x"3EC4CB96",
    x"3EC4D730",
    x"3EC4E2C9",
    x"3EC4EE63",
    x"3EC4F9FD",
    x"3EC50596",
    x"3EC5112F",
    x"3EC51CC8",
    x"3EC52861",
    x"3EC533FA",
    x"3EC53F93",
    x"3EC54B2B",
    x"3EC556C4",
    x"3EC5625C",
    x"3EC56DF4",
    x"3EC5798D",
    x"3EC58525",
    x"3EC590BD",
    x"3EC59C54",
    x"3EC5A7EC",
    x"3EC5B384",
    x"3EC5BF1B",
    x"3EC5CAB2",
    x"3EC5D649",
    x"3EC5E1E1",
    x"3EC5ED77",
    x"3EC5F90E",
    x"3EC604A5",
    x"3EC6103C",
    x"3EC61BD2",
    x"3EC62768",
    x"3EC632FF",
    x"3EC63E95",
    x"3EC64A2B",
    x"3EC655C1",
    x"3EC66156",
    x"3EC66CEC",
    x"3EC67882",
    x"3EC68417",
    x"3EC68FAC",
    x"3EC69B41",
    x"3EC6A6D6",
    x"3EC6B26B",
    x"3EC6BE00",
    x"3EC6C995",
    x"3EC6D529",
    x"3EC6E0BE",
    x"3EC6EC52",
    x"3EC6F7E6",
    x"3EC7037B",
    x"3EC70F0E",
    x"3EC71AA2",
    x"3EC72636",
    x"3EC731CA",
    x"3EC73D5D",
    x"3EC748F0",
    x"3EC75484",
    x"3EC76017",
    x"3EC76BAA",
    x"3EC7773D",
    x"3EC782D0",
    x"3EC78E62",
    x"3EC799F5",
    x"3EC7A587",
    x"3EC7B119",
    x"3EC7BCAC",
    x"3EC7C83E",
    x"3EC7D3CF",
    x"3EC7DF61",
    x"3EC7EAF3",
    x"3EC7F685",
    x"3EC80216",
    x"3EC80DA7",
    x"3EC81938",
    x"3EC824CA",
    x"3EC8305B",
    x"3EC83BEB",
    x"3EC8477C",
    x"3EC8530D",
    x"3EC85E9D",
    x"3EC86A2D",
    x"3EC875BE",
    x"3EC8814E",
    x"3EC88CDE",
    x"3EC8986E",
    x"3EC8A3FD",
    x"3EC8AF8D",
    x"3EC8BB1D",
    x"3EC8C6AC",
    x"3EC8D23B",
    x"3EC8DDCA",
    x"3EC8E959",
    x"3EC8F4E8",
    x"3EC90077",
    x"3EC90C06",
    x"3EC91794",
    x"3EC92323",
    x"3EC92EB1",
    x"3EC93A3F",
    x"3EC945CD",
    x"3EC9515B",
    x"3EC95CE9",
    x"3EC96877",
    x"3EC97404",
    x"3EC97F92",
    x"3EC98B1F",
    x"3EC996AC",
    x"3EC9A239",
    x"3EC9ADC6",
    x"3EC9B953",
    x"3EC9C4E0",
    x"3EC9D06C",
    x"3EC9DBF9",
    x"3EC9E785",
    x"3EC9F312",
    x"3EC9FE9E",
    x"3ECA0A2A",
    x"3ECA15B5",
    x"3ECA2141",
    x"3ECA2CCD",
    x"3ECA3858",
    x"3ECA43E4",
    x"3ECA4F6F",
    x"3ECA5AFA",
    x"3ECA6685",
    x"3ECA7210",
    x"3ECA7D9B",
    x"3ECA8925",
    x"3ECA94B0",
    x"3ECAA03A",
    x"3ECAABC5",
    x"3ECAB74F",
    x"3ECAC2D9",
    x"3ECACE63",
    x"3ECAD9ED",
    x"3ECAE576",
    x"3ECAF100",
    x"3ECAFC89",
    x"3ECB0813",
    x"3ECB139C",
    x"3ECB1F25",
    x"3ECB2AAE",
    x"3ECB3637",
    x"3ECB41BF",
    x"3ECB4D48",
    x"3ECB58D0",
    x"3ECB6459",
    x"3ECB6FE1",
    x"3ECB7B69",
    x"3ECB86F1",
    x"3ECB9279",
    x"3ECB9E00",
    x"3ECBA988",
    x"3ECBB50F",
    x"3ECBC097",
    x"3ECBCC1E",
    x"3ECBD7A5",
    x"3ECBE32C",
    x"3ECBEEB3",
    x"3ECBFA3A",
    x"3ECC05C0",
    x"3ECC1147",
    x"3ECC1CCD",
    x"3ECC2853",
    x"3ECC33DA",
    x"3ECC3F60",
    x"3ECC4AE5",
    x"3ECC566B",
    x"3ECC61F1",
    x"3ECC6D76",
    x"3ECC78FC",
    x"3ECC8481",
    x"3ECC9006",
    x"3ECC9B8B",
    x"3ECCA710",
    x"3ECCB295",
    x"3ECCBE19",
    x"3ECCC99E",
    x"3ECCD522",
    x"3ECCE0A7",
    x"3ECCEC2B",
    x"3ECCF7AF",
    x"3ECD0333",
    x"3ECD0EB6",
    x"3ECD1A3A",
    x"3ECD25BE",
    x"3ECD3141",
    x"3ECD3CC4",
    x"3ECD4847",
    x"3ECD53CA",
    x"3ECD5F4D",
    x"3ECD6AD0",
    x"3ECD7653",
    x"3ECD81D5",
    x"3ECD8D58",
    x"3ECD98DA",
    x"3ECDA45C",
    x"3ECDAFDE",
    x"3ECDBB60",
    x"3ECDC6E2",
    x"3ECDD264",
    x"3ECDDDE5",
    x"3ECDE967",
    x"3ECDF4E8",
    x"3ECE0069",
    x"3ECE0BEA",
    x"3ECE176B",
    x"3ECE22EC",
    x"3ECE2E6D",
    x"3ECE39ED",
    x"3ECE456E",
    x"3ECE50EE",
    x"3ECE5C6E",
    x"3ECE67EE",
    x"3ECE736E",
    x"3ECE7EEE",
    x"3ECE8A6E",
    x"3ECE95ED",
    x"3ECEA16D",
    x"3ECEACEC",
    x"3ECEB86B",
    x"3ECEC3EA",
    x"3ECECF69",
    x"3ECEDAE8",
    x"3ECEE667",
    x"3ECEF1E5",
    x"3ECEFD64",
    x"3ECF08E2",
    x"3ECF1460",
    x"3ECF1FDE",
    x"3ECF2B5C",
    x"3ECF36DA",
    x"3ECF4258",
    x"3ECF4DD5",
    x"3ECF5953",
    x"3ECF64D0",
    x"3ECF704D",
    x"3ECF7BCA",
    x"3ECF8747",
    x"3ECF92C4",
    x"3ECF9E41",
    x"3ECFA9BD",
    x"3ECFB53A",
    x"3ECFC0B6",
    x"3ECFCC32",
    x"3ECFD7AE",
    x"3ECFE32A",
    x"3ECFEEA6",
    x"3ECFFA22",
    x"3ED0059D",
    x"3ED01119",
    x"3ED01C94",
    x"3ED0280F",
    x"3ED0338A",
    x"3ED03F05",
    x"3ED04A80",
    x"3ED055FB",
    x"3ED06175",
    x"3ED06CF0",
    x"3ED0786A",
    x"3ED083E4",
    x"3ED08F5E",
    x"3ED09AD8",
    x"3ED0A652",
    x"3ED0B1CC",
    x"3ED0BD45",
    x"3ED0C8BF",
    x"3ED0D438",
    x"3ED0DFB1",
    x"3ED0EB2A",
    x"3ED0F6A3",
    x"3ED1021C",
    x"3ED10D95",
    x"3ED1190D",
    x"3ED12485",
    x"3ED12FFE",
    x"3ED13B76",
    x"3ED146EE",
    x"3ED15266",
    x"3ED15DDE",
    x"3ED16955",
    x"3ED174CD",
    x"3ED18044",
    x"3ED18BBC",
    x"3ED19733",
    x"3ED1A2AA",
    x"3ED1AE21",
    x"3ED1B998",
    x"3ED1C50E",
    x"3ED1D085",
    x"3ED1DBFB",
    x"3ED1E771",
    x"3ED1F2E8",
    x"3ED1FE5E",
    x"3ED209D3",
    x"3ED21549",
    x"3ED220BF",
    x"3ED22C34",
    x"3ED237AA",
    x"3ED2431F",
    x"3ED24E94",
    x"3ED25A09",
    x"3ED2657E",
    x"3ED270F3",
    x"3ED27C68",
    x"3ED287DC",
    x"3ED29350",
    x"3ED29EC5",
    x"3ED2AA39",
    x"3ED2B5AD",
    x"3ED2C121",
    x"3ED2CC94",
    x"3ED2D808",
    x"3ED2E37C",
    x"3ED2EEEF",
    x"3ED2FA62",
    x"3ED305D5",
    x"3ED31148",
    x"3ED31CBB",
    x"3ED3282E",
    x"3ED333A0",
    x"3ED33F13",
    x"3ED34A85",
    x"3ED355F7",
    x"3ED3616A",
    x"3ED36CDB",
    x"3ED3784D",
    x"3ED383BF",
    x"3ED38F31",
    x"3ED39AA2",
    x"3ED3A613",
    x"3ED3B185",
    x"3ED3BCF6",
    x"3ED3C867",
    x"3ED3D3D7",
    x"3ED3DF48",
    x"3ED3EAB9",
    x"3ED3F629",
    x"3ED40199",
    x"3ED40D0A",
    x"3ED4187A",
    x"3ED423EA",
    x"3ED42F59",
    x"3ED43AC9",
    x"3ED44639",
    x"3ED451A8",
    x"3ED45D17",
    x"3ED46886",
    x"3ED473F5",
    x"3ED47F64",
    x"3ED48AD3",
    x"3ED49642",
    x"3ED4A1B0",
    x"3ED4AD1F",
    x"3ED4B88D",
    x"3ED4C3FB",
    x"3ED4CF69",
    x"3ED4DAD7",
    x"3ED4E645",
    x"3ED4F1B2",
    x"3ED4FD20",
    x"3ED5088D",
    x"3ED513FA",
    x"3ED51F68",
    x"3ED52AD5",
    x"3ED53641",
    x"3ED541AE",
    x"3ED54D1B",
    x"3ED55887",
    x"3ED563F3",
    x"3ED56F60",
    x"3ED57ACC",
    x"3ED58638",
    x"3ED591A4",
    x"3ED59D0F",
    x"3ED5A87B",
    x"3ED5B3E6",
    x"3ED5BF52",
    x"3ED5CABD",
    x"3ED5D628",
    x"3ED5E193",
    x"3ED5ECFD",
    x"3ED5F868",
    x"3ED603D3",
    x"3ED60F3D",
    x"3ED61AA7",
    x"3ED62611",
    x"3ED6317B",
    x"3ED63CE5",
    x"3ED6484F",
    x"3ED653B9",
    x"3ED65F22",
    x"3ED66A8C",
    x"3ED675F5",
    x"3ED6815E",
    x"3ED68CC7",
    x"3ED69830",
    x"3ED6A399",
    x"3ED6AF01",
    x"3ED6BA6A",
    x"3ED6C5D2",
    x"3ED6D13A",
    x"3ED6DCA2",
    x"3ED6E80A",
    x"3ED6F372",
    x"3ED6FEDA",
    x"3ED70A41",
    x"3ED715A9",
    x"3ED72110",
    x"3ED72C77",
    x"3ED737DE",
    x"3ED74345",
    x"3ED74EAC",
    x"3ED75A13",
    x"3ED76579",
    x"3ED770E0",
    x"3ED77C46",
    x"3ED787AC",
    x"3ED79312",
    x"3ED79E78",
    x"3ED7A9DE",
    x"3ED7B543",
    x"3ED7C0A9",
    x"3ED7CC0E",
    x"3ED7D773",
    x"3ED7E2D8",
    x"3ED7EE3D",
    x"3ED7F9A2",
    x"3ED80507",
    x"3ED8106B",
    x"3ED81BD0",
    x"3ED82734",
    x"3ED83298",
    x"3ED83DFC",
    x"3ED84960",
    x"3ED854C4",
    x"3ED86028",
    x"3ED86B8B",
    x"3ED876EF",
    x"3ED88252",
    x"3ED88DB5",
    x"3ED89918",
    x"3ED8A47B",
    x"3ED8AFDE",
    x"3ED8BB40",
    x"3ED8C6A3",
    x"3ED8D205",
    x"3ED8DD67",
    x"3ED8E8CA",
    x"3ED8F42C",
    x"3ED8FF8D",
    x"3ED90AEF",
    x"3ED91651",
    x"3ED921B2",
    x"3ED92D13",
    x"3ED93875",
    x"3ED943D6",
    x"3ED94F37",
    x"3ED95A97",
    x"3ED965F8",
    x"3ED97159",
    x"3ED97CB9",
    x"3ED98819",
    x"3ED99379",
    x"3ED99ED9",
    x"3ED9AA39",
    x"3ED9B599",
    x"3ED9C0F9",
    x"3ED9CC58",
    x"3ED9D7B7",
    x"3ED9E317",
    x"3ED9EE76",
    x"3ED9F9D5",
    x"3EDA0533",
    x"3EDA1092",
    x"3EDA1BF1",
    x"3EDA274F",
    x"3EDA32AD",
    x"3EDA3E0C",
    x"3EDA496A",
    x"3EDA54C8",
    x"3EDA6025",
    x"3EDA6B83",
    x"3EDA76E0",
    x"3EDA823E",
    x"3EDA8D9B",
    x"3EDA98F8",
    x"3EDAA455",
    x"3EDAAFB2",
    x"3EDABB0F",
    x"3EDAC66B",
    x"3EDAD1C8",
    x"3EDADD24",
    x"3EDAE880",
    x"3EDAF3DC",
    x"3EDAFF38",
    x"3EDB0A94",
    x"3EDB15F0",
    x"3EDB214B",
    x"3EDB2CA7",
    x"3EDB3802",
    x"3EDB435D",
    x"3EDB4EB8",
    x"3EDB5A13",
    x"3EDB656E",
    x"3EDB70C8",
    x"3EDB7C23",
    x"3EDB877D",
    x"3EDB92D7",
    x"3EDB9E31",
    x"3EDBA98B",
    x"3EDBB4E5",
    x"3EDBC03F",
    x"3EDBCB98",
    x"3EDBD6F2",
    x"3EDBE24B",
    x"3EDBEDA4",
    x"3EDBF8FD",
    x"3EDC0456",
    x"3EDC0FAF",
    x"3EDC1B08",
    x"3EDC2660",
    x"3EDC31B8",
    x"3EDC3D11",
    x"3EDC4869",
    x"3EDC53C1",
    x"3EDC5F18",
    x"3EDC6A70",
    x"3EDC75C8",
    x"3EDC811F",
    x"3EDC8C76",
    x"3EDC97CE",
    x"3EDCA325",
    x"3EDCAE7C",
    x"3EDCB9D2",
    x"3EDCC529",
    x"3EDCD07F",
    x"3EDCDBD6",
    x"3EDCE72C",
    x"3EDCF282",
    x"3EDCFDD8",
    x"3EDD092E",
    x"3EDD1484",
    x"3EDD1FD9",
    x"3EDD2B2F",
    x"3EDD3684",
    x"3EDD41D9",
    x"3EDD4D2E",
    x"3EDD5883",
    x"3EDD63D8",
    x"3EDD6F2C",
    x"3EDD7A81",
    x"3EDD85D5",
    x"3EDD912A",
    x"3EDD9C7E",
    x"3EDDA7D2",
    x"3EDDB325",
    x"3EDDBE79",
    x"3EDDC9CD",
    x"3EDDD520",
    x"3EDDE073",
    x"3EDDEBC7",
    x"3EDDF71A",
    x"3EDE026C",
    x"3EDE0DBF",
    x"3EDE1912",
    x"3EDE2464",
    x"3EDE2FB7",
    x"3EDE3B09",
    x"3EDE465B",
    x"3EDE51AD",
    x"3EDE5CFF",
    x"3EDE6851",
    x"3EDE73A2",
    x"3EDE7EF3",
    x"3EDE8A45",
    x"3EDE9596",
    x"3EDEA0E7",
    x"3EDEAC38",
    x"3EDEB789",
    x"3EDEC2D9",
    x"3EDECE2A",
    x"3EDED97A",
    x"3EDEE4CA",
    x"3EDEF01A",
    x"3EDEFB6A",
    x"3EDF06BA",
    x"3EDF120A",
    x"3EDF1D59",
    x"3EDF28A9",
    x"3EDF33F8",
    x"3EDF3F47",
    x"3EDF4A96",
    x"3EDF55E5",
    x"3EDF6134",
    x"3EDF6C82",
    x"3EDF77D1",
    x"3EDF831F",
    x"3EDF8E6D",
    x"3EDF99BB",
    x"3EDFA509",
    x"3EDFB057",
    x"3EDFBBA5",
    x"3EDFC6F2",
    x"3EDFD240",
    x"3EDFDD8D",
    x"3EDFE8DA",
    x"3EDFF427",
    x"3EDFFF74",
    x"3EE00AC1",
    x"3EE0160D",
    x"3EE0215A",
    x"3EE02CA6",
    x"3EE037F2",
    x"3EE0433E",
    x"3EE04E8A",
    x"3EE059D6",
    x"3EE06522",
    x"3EE0706D",
    x"3EE07BB8",
    x"3EE08704",
    x"3EE0924F",
    x"3EE09D9A",
    x"3EE0A8E5",
    x"3EE0B42F",
    x"3EE0BF7A",
    x"3EE0CAC4",
    x"3EE0D60E",
    x"3EE0E159",
    x"3EE0ECA3",
    x"3EE0F7ED",
    x"3EE10336",
    x"3EE10E80",
    x"3EE119C9",
    x"3EE12513",
    x"3EE1305C",
    x"3EE13BA5",
    x"3EE146EE",
    x"3EE15237",
    x"3EE15D7F",
    x"3EE168C8",
    x"3EE17410",
    x"3EE17F58",
    x"3EE18AA1",
    x"3EE195E9",
    x"3EE1A130",
    x"3EE1AC78",
    x"3EE1B7C0",
    x"3EE1C307",
    x"3EE1CE4E",
    x"3EE1D996",
    x"3EE1E4DD",
    x"3EE1F023",
    x"3EE1FB6A",
    x"3EE206B1",
    x"3EE211F7",
    x"3EE21D3E",
    x"3EE22884",
    x"3EE233CA",
    x"3EE23F10",
    x"3EE24A56",
    x"3EE2559B",
    x"3EE260E1",
    x"3EE26C26",
    x"3EE2776C",
    x"3EE282B1",
    x"3EE28DF6",
    x"3EE2993A",
    x"3EE2A47F",
    x"3EE2AFC4",
    x"3EE2BB08",
    x"3EE2C64C",
    x"3EE2D191",
    x"3EE2DCD5",
    x"3EE2E819",
    x"3EE2F35C",
    x"3EE2FEA0",
    x"3EE309E3",
    x"3EE31527",
    x"3EE3206A",
    x"3EE32BAD",
    x"3EE336F0",
    x"3EE34233",
    x"3EE34D75",
    x"3EE358B8",
    x"3EE363FA",
    x"3EE36F3D",
    x"3EE37A7F",
    x"3EE385C1",
    x"3EE39102",
    x"3EE39C44",
    x"3EE3A786",
    x"3EE3B2C7",
    x"3EE3BE08",
    x"3EE3C94A",
    x"3EE3D48B",
    x"3EE3DFCB",
    x"3EE3EB0C",
    x"3EE3F64D",
    x"3EE4018D",
    x"3EE40CCE",
    x"3EE4180E",
    x"3EE4234E",
    x"3EE42E8E",
    x"3EE439CE",
    x"3EE4450D",
    x"3EE4504D",
    x"3EE45B8C",
    x"3EE466CB",
    x"3EE4720A",
    x"3EE47D49",
    x"3EE48888",
    x"3EE493C7",
    x"3EE49F05",
    x"3EE4AA44",
    x"3EE4B582",
    x"3EE4C0C0",
    x"3EE4CBFE",
    x"3EE4D73C",
    x"3EE4E27A",
    x"3EE4EDB7",
    x"3EE4F8F5",
    x"3EE50432",
    x"3EE50F6F",
    x"3EE51AAC",
    x"3EE525E9",
    x"3EE53126",
    x"3EE53C62",
    x"3EE5479F",
    x"3EE552DB",
    x"3EE55E17",
    x"3EE56953",
    x"3EE5748F",
    x"3EE57FCB",
    x"3EE58B07",
    x"3EE59642",
    x"3EE5A17E",
    x"3EE5ACB9",
    x"3EE5B7F4",
    x"3EE5C32F",
    x"3EE5CE6A",
    x"3EE5D9A4",
    x"3EE5E4DF",
    x"3EE5F019",
    x"3EE5FB54",
    x"3EE6068E",
    x"3EE611C8",
    x"3EE61D02",
    x"3EE6283B",
    x"3EE63375",
    x"3EE63EAE",
    x"3EE649E7",
    x"3EE65521",
    x"3EE6605A",
    x"3EE66B93",
    x"3EE676CB",
    x"3EE68204",
    x"3EE68D3C",
    x"3EE69875",
    x"3EE6A3AD",
    x"3EE6AEE5",
    x"3EE6BA1D",
    x"3EE6C554",
    x"3EE6D08C",
    x"3EE6DBC4",
    x"3EE6E6FB",
    x"3EE6F232",
    x"3EE6FD69",
    x"3EE708A0",
    x"3EE713D7",
    x"3EE71F0E",
    x"3EE72A44",
    x"3EE7357A",
    x"3EE740B1",
    x"3EE74BE7",
    x"3EE7571D",
    x"3EE76253",
    x"3EE76D88",
    x"3EE778BE",
    x"3EE783F3",
    x"3EE78F28",
    x"3EE79A5D",
    x"3EE7A592",
    x"3EE7B0C7",
    x"3EE7BBFC",
    x"3EE7C731",
    x"3EE7D265",
    x"3EE7DD99",
    x"3EE7E8CD",
    x"3EE7F401",
    x"3EE7FF35",
    x"3EE80A69",
    x"3EE8159C",
    x"3EE820D0",
    x"3EE82C03",
    x"3EE83736",
    x"3EE84269",
    x"3EE84D9C",
    x"3EE858CF",
    x"3EE86402",
    x"3EE86F34",
    x"3EE87A66",
    x"3EE88599",
    x"3EE890CB",
    x"3EE89BFD",
    x"3EE8A72E",
    x"3EE8B260",
    x"3EE8BD91",
    x"3EE8C8C3",
    x"3EE8D3F4",
    x"3EE8DF25",
    x"3EE8EA56",
    x"3EE8F587",
    x"3EE900B7",
    x"3EE90BE8",
    x"3EE91718",
    x"3EE92248",
    x"3EE92D78",
    x"3EE938A8",
    x"3EE943D8",
    x"3EE94F08",
    x"3EE95A37",
    x"3EE96567",
    x"3EE97096",
    x"3EE97BC5",
    x"3EE986F4",
    x"3EE99223",
    x"3EE99D51",
    x"3EE9A880",
    x"3EE9B3AE",
    x"3EE9BEDD",
    x"3EE9CA0B",
    x"3EE9D539",
    x"3EE9E066",
    x"3EE9EB94",
    x"3EE9F6C2",
    x"3EEA01EF",
    x"3EEA0D1C",
    x"3EEA1849",
    x"3EEA2376",
    x"3EEA2EA3",
    x"3EEA39D0",
    x"3EEA44FD",
    x"3EEA5029",
    x"3EEA5B55",
    x"3EEA6681",
    x"3EEA71AD",
    x"3EEA7CD9",
    x"3EEA8805",
    x"3EEA9330",
    x"3EEA9E5C",
    x"3EEAA987",
    x"3EEAB4B2",
    x"3EEABFDD",
    x"3EEACB08",
    x"3EEAD633",
    x"3EEAE15D",
    x"3EEAEC88",
    x"3EEAF7B2",
    x"3EEB02DC",
    x"3EEB0E06",
    x"3EEB1930",
    x"3EEB245A",
    x"3EEB2F84",
    x"3EEB3AAD",
    x"3EEB45D6",
    x"3EEB50FF",
    x"3EEB5C28",
    x"3EEB6751",
    x"3EEB727A",
    x"3EEB7DA3",
    x"3EEB88CB",
    x"3EEB93F3",
    x"3EEB9F1C",
    x"3EEBAA44",
    x"3EEBB56C",
    x"3EEBC093",
    x"3EEBCBBB",
    x"3EEBD6E2",
    x"3EEBE20A",
    x"3EEBED31",
    x"3EEBF858",
    x"3EEC037F",
    x"3EEC0EA5",
    x"3EEC19CC",
    x"3EEC24F3",
    x"3EEC3019",
    x"3EEC3B3F",
    x"3EEC4665",
    x"3EEC518B",
    x"3EEC5CB1",
    x"3EEC67D6",
    x"3EEC72FC",
    x"3EEC7E21",
    x"3EEC8946",
    x"3EEC946B",
    x"3EEC9F90",
    x"3EECAAB5",
    x"3EECB5DA",
    x"3EECC0FE",
    x"3EECCC22",
    x"3EECD747",
    x"3EECE26B",
    x"3EECED8F",
    x"3EECF8B2",
    x"3EED03D6",
    x"3EED0EF9",
    x"3EED1A1D",
    x"3EED2540",
    x"3EED3063",
    x"3EED3B86",
    x"3EED46A9",
    x"3EED51CB",
    x"3EED5CEE",
    x"3EED6810",
    x"3EED7332",
    x"3EED7E54",
    x"3EED8976",
    x"3EED9498",
    x"3EED9FB9",
    x"3EEDAADB",
    x"3EEDB5FC",
    x"3EEDC11D",
    x"3EEDCC3E",
    x"3EEDD75F",
    x"3EEDE280",
    x"3EEDEDA1",
    x"3EEDF8C1",
    x"3EEE03E2",
    x"3EEE0F02",
    x"3EEE1A22",
    x"3EEE2542",
    x"3EEE3061",
    x"3EEE3B81",
    x"3EEE46A0",
    x"3EEE51C0",
    x"3EEE5CDF",
    x"3EEE67FE",
    x"3EEE731D",
    x"3EEE7E3C",
    x"3EEE895A",
    x"3EEE9479",
    x"3EEE9F97",
    x"3EEEAAB5",
    x"3EEEB5D3",
    x"3EEEC0F1",
    x"3EEECC0F",
    x"3EEED72C",
    x"3EEEE24A",
    x"3EEEED67",
    x"3EEEF884",
    x"3EEF03A1",
    x"3EEF0EBE",
    x"3EEF19DB",
    x"3EEF24F7",
    x"3EEF3014",
    x"3EEF3B30",
    x"3EEF464C",
    x"3EEF5168",
    x"3EEF5C84",
    x"3EEF67A0",
    x"3EEF72BC",
    x"3EEF7DD7",
    x"3EEF88F2",
    x"3EEF940D",
    x"3EEF9F28",
    x"3EEFAA43",
    x"3EEFB55E",
    x"3EEFC079",
    x"3EEFCB93",
    x"3EEFD6AD",
    x"3EEFE1C7",
    x"3EEFECE1",
    x"3EEFF7FB",
    x"3EF00315",
    x"3EF00E2E",
    x"3EF01948",
    x"3EF02461",
    x"3EF02F7A",
    x"3EF03A93",
    x"3EF045AC",
    x"3EF050C5",
    x"3EF05BDD",
    x"3EF066F6",
    x"3EF0720E",
    x"3EF07D26",
    x"3EF0883E",
    x"3EF09356",
    x"3EF09E6E",
    x"3EF0A985",
    x"3EF0B49C",
    x"3EF0BFB4",
    x"3EF0CACB",
    x"3EF0D5E2",
    x"3EF0E0F9",
    x"3EF0EC0F",
    x"3EF0F726",
    x"3EF1023C",
    x"3EF10D52",
    x"3EF11868",
    x"3EF1237E",
    x"3EF12E94",
    x"3EF139AA",
    x"3EF144BF",
    x"3EF14FD5",
    x"3EF15AEA",
    x"3EF165FF",
    x"3EF17114",
    x"3EF17C28",
    x"3EF1873D",
    x"3EF19252",
    x"3EF19D66",
    x"3EF1A87A",
    x"3EF1B38E",
    x"3EF1BEA2",
    x"3EF1C9B6",
    x"3EF1D4C9",
    x"3EF1DFDD",
    x"3EF1EAF0",
    x"3EF1F603",
    x"3EF20116",
    x"3EF20C29",
    x"3EF2173C",
    x"3EF2224F",
    x"3EF22D61",
    x"3EF23873",
    x"3EF24385",
    x"3EF24E97",
    x"3EF259A9",
    x"3EF264BB",
    x"3EF26FCD",
    x"3EF27ADE",
    x"3EF285EF",
    x"3EF29100",
    x"3EF29C11",
    x"3EF2A722",
    x"3EF2B233",
    x"3EF2BD43",
    x"3EF2C854",
    x"3EF2D364",
    x"3EF2DE74",
    x"3EF2E984",
    x"3EF2F494",
    x"3EF2FFA4",
    x"3EF30AB3",
    x"3EF315C2",
    x"3EF320D2",
    x"3EF32BE1",
    x"3EF336F0",
    x"3EF341FE",
    x"3EF34D0D",
    x"3EF3581C",
    x"3EF3632A",
    x"3EF36E38",
    x"3EF37946",
    x"3EF38454",
    x"3EF38F62",
    x"3EF39A6F",
    x"3EF3A57D",
    x"3EF3B08A",
    x"3EF3BB97",
    x"3EF3C6A4",
    x"3EF3D1B1",
    x"3EF3DCBE",
    x"3EF3E7CB",
    x"3EF3F2D7",
    x"3EF3FDE3",
    x"3EF408F0",
    x"3EF413FB",
    x"3EF41F07",
    x"3EF42A13",
    x"3EF4351F",
    x"3EF4402A",
    x"3EF44B35",
    x"3EF45640",
    x"3EF4614B",
    x"3EF46C56",
    x"3EF47761",
    x"3EF4826B",
    x"3EF48D76",
    x"3EF49880",
    x"3EF4A38A",
    x"3EF4AE94",
    x"3EF4B99E",
    x"3EF4C4A7",
    x"3EF4CFB1",
    x"3EF4DABA",
    x"3EF4E5C3",
    x"3EF4F0CC",
    x"3EF4FBD5",
    x"3EF506DE",
    x"3EF511E7",
    x"3EF51CEF",
    x"3EF527F8",
    x"3EF53300",
    x"3EF53E08",
    x"3EF54910",
    x"3EF55417",
    x"3EF55F1F",
    x"3EF56A26",
    x"3EF5752E",
    x"3EF58035",
    x"3EF58B3C",
    x"3EF59643",
    x"3EF5A149",
    x"3EF5AC50",
    x"3EF5B756",
    x"3EF5C25C",
    x"3EF5CD62",
    x"3EF5D868",
    x"3EF5E36E",
    x"3EF5EE74",
    x"3EF5F979",
    x"3EF6047F",
    x"3EF60F84",
    x"3EF61A89",
    x"3EF6258E",
    x"3EF63093",
    x"3EF63B97",
    x"3EF6469C",
    x"3EF651A0",
    x"3EF65CA4",
    x"3EF667A8",
    x"3EF672AC",
    x"3EF67DB0",
    x"3EF688B3",
    x"3EF693B7",
    x"3EF69EBA",
    x"3EF6A9BD",
    x"3EF6B4C0",
    x"3EF6BFC3",
    x"3EF6CAC6",
    x"3EF6D5C8",
    x"3EF6E0CB",
    x"3EF6EBCD",
    x"3EF6F6CF",
    x"3EF701D1",
    x"3EF70CD3",
    x"3EF717D4",
    x"3EF722D6",
    x"3EF72DD7",
    x"3EF738D8",
    x"3EF743D9",
    x"3EF74EDA",
    x"3EF759DB",
    x"3EF764DC",
    x"3EF76FDC",
    x"3EF77ADC",
    x"3EF785DC",
    x"3EF790DC",
    x"3EF79BDC",
    x"3EF7A6DC",
    x"3EF7B1DC",
    x"3EF7BCDB",
    x"3EF7C7DA",
    x"3EF7D2D9",
    x"3EF7DDD8",
    x"3EF7E8D7",
    x"3EF7F3D6",
    x"3EF7FED4",
    x"3EF809D3",
    x"3EF814D1",
    x"3EF81FCF",
    x"3EF82ACD",
    x"3EF835CB",
    x"3EF840C8",
    x"3EF84BC6",
    x"3EF856C3",
    x"3EF861C0",
    x"3EF86CBD",
    x"3EF877BA",
    x"3EF882B7",
    x"3EF88DB3",
    x"3EF898B0",
    x"3EF8A3AC",
    x"3EF8AEA8",
    x"3EF8B9A4",
    x"3EF8C4A0",
    x"3EF8CF9C",
    x"3EF8DA97",
    x"3EF8E592",
    x"3EF8F08E",
    x"3EF8FB89",
    x"3EF90684",
    x"3EF9117E",
    x"3EF91C79",
    x"3EF92773",
    x"3EF9326E",
    x"3EF93D68",
    x"3EF94862",
    x"3EF9535C",
    x"3EF95E56",
    x"3EF9694F",
    x"3EF97449",
    x"3EF97F42",
    x"3EF98A3B",
    x"3EF99534",
    x"3EF9A02D",
    x"3EF9AB25",
    x"3EF9B61E",
    x"3EF9C116",
    x"3EF9CC0E",
    x"3EF9D707",
    x"3EF9E1FE",
    x"3EF9ECF6",
    x"3EF9F7EE",
    x"3EFA02E5",
    x"3EFA0DDD",
    x"3EFA18D4",
    x"3EFA23CB",
    x"3EFA2EC2",
    x"3EFA39B8",
    x"3EFA44AF",
    x"3EFA4FA5",
    x"3EFA5A9C",
    x"3EFA6592",
    x"3EFA7088",
    x"3EFA7B7D",
    x"3EFA8673",
    x"3EFA9169",
    x"3EFA9C5E",
    x"3EFAA753",
    x"3EFAB248",
    x"3EFABD3D",
    x"3EFAC832",
    x"3EFAD326",
    x"3EFADE1B",
    x"3EFAE90F",
    x"3EFAF403",
    x"3EFAFEF7",
    x"3EFB09EB",
    x"3EFB14DF",
    x"3EFB1FD2",
    x"3EFB2AC6",
    x"3EFB35B9",
    x"3EFB40AC",
    x"3EFB4B9F",
    x"3EFB5692",
    x"3EFB6184",
    x"3EFB6C77",
    x"3EFB7769",
    x"3EFB825B",
    x"3EFB8D4D",
    x"3EFB983F",
    x"3EFBA331",
    x"3EFBAE22",
    x"3EFBB914",
    x"3EFBC405",
    x"3EFBCEF6",
    x"3EFBD9E7",
    x"3EFBE4D8",
    x"3EFBEFC9",
    x"3EFBFAB9",
    x"3EFC05AA",
    x"3EFC109A",
    x"3EFC1B8A",
    x"3EFC267A",
    x"3EFC3169",
    x"3EFC3C59",
    x"3EFC4748",
    x"3EFC5238",
    x"3EFC5D27",
    x"3EFC6816",
    x"3EFC7305",
    x"3EFC7DF3",
    x"3EFC88E2",
    x"3EFC93D0",
    x"3EFC9EBF",
    x"3EFCA9AD",
    x"3EFCB49B",
    x"3EFCBF88",
    x"3EFCCA76",
    x"3EFCD563",
    x"3EFCE051",
    x"3EFCEB3E",
    x"3EFCF62B",
    x"3EFD0118",
    x"3EFD0C04",
    x"3EFD16F1",
    x"3EFD21DD",
    x"3EFD2CCA",
    x"3EFD37B6",
    x"3EFD42A2",
    x"3EFD4D8D",
    x"3EFD5879",
    x"3EFD6365",
    x"3EFD6E50",
    x"3EFD793B",
    x"3EFD8426",
    x"3EFD8F11",
    x"3EFD99FC",
    x"3EFDA4E6",
    x"3EFDAFD1",
    x"3EFDBABB",
    x"3EFDC5A5",
    x"3EFDD08F",
    x"3EFDDB79",
    x"3EFDE662",
    x"3EFDF14C",
    x"3EFDFC35",
    x"3EFE071E",
    x"3EFE1207",
    x"3EFE1CF0",
    x"3EFE27D9",
    x"3EFE32C2",
    x"3EFE3DAA",
    x"3EFE4892",
    x"3EFE537A",
    x"3EFE5E62",
    x"3EFE694A",
    x"3EFE7432",
    x"3EFE7F19",
    x"3EFE8A01",
    x"3EFE94E8",
    x"3EFE9FCF",
    x"3EFEAAB6",
    x"3EFEB59D",
    x"3EFEC083",
    x"3EFECB6A",
    x"3EFED650",
    x"3EFEE136",
    x"3EFEEC1C",
    x"3EFEF702",
    x"3EFF01E8",
    x"3EFF0CCD",
    x"3EFF17B2",
    x"3EFF2298",
    x"3EFF2D7D",
    x"3EFF3862",
    x"3EFF4346",
    x"3EFF4E2B",
    x"3EFF590F",
    x"3EFF63F4",
    x"3EFF6ED8",
    x"3EFF79BC",
    x"3EFF849F",
    x"3EFF8F83",
    x"3EFF9A67",
    x"3EFFA54A",
    x"3EFFB02D",
    x"3EFFBB10",
    x"3EFFC5F3",
    x"3EFFD0D6",
    x"3EFFDBB8",
    x"3EFFE69B",
    x"3EFFF17D",
    x"3EFFFC5F",
    x"3F0003A1",
    x"3F000912",
    x"3F000E82",
    x"3F0013F3",
    x"3F001964",
    x"3F001ED4",
    x"3F002445",
    x"3F0029B5",
    x"3F002F26",
    x"3F003496",
    x"3F003A06",
    x"3F003F76",
    x"3F0044E6",
    x"3F004A56",
    x"3F004FC6",
    x"3F005536",
    x"3F005AA6",
    x"3F006016",
    x"3F006585",
    x"3F006AF5",
    x"3F007064",
    x"3F0075D4",
    x"3F007B43",
    x"3F0080B2",
    x"3F008621",
    x"3F008B90",
    x"3F0090FF",
    x"3F00966E",
    x"3F009BDD",
    x"3F00A14C",
    x"3F00A6BA",
    x"3F00AC29",
    x"3F00B197",
    x"3F00B706",
    x"3F00BC74",
    x"3F00C1E2",
    x"3F00C751",
    x"3F00CCBF",
    x"3F00D22D",
    x"3F00D79B",
    x"3F00DD09",
    x"3F00E276",
    x"3F00E7E4",
    x"3F00ED52",
    x"3F00F2BF",
    x"3F00F82D",
    x"3F00FD9A",
    x"3F010308",
    x"3F010875",
    x"3F010DE2",
    x"3F01134F",
    x"3F0118BC",
    x"3F011E29",
    x"3F012396",
    x"3F012903",
    x"3F012E70",
    x"3F0133DC",
    x"3F013949",
    x"3F013EB5",
    x"3F014422",
    x"3F01498E",
    x"3F014EFA",
    x"3F015467",
    x"3F0159D3",
    x"3F015F3F",
    x"3F0164AB",
    x"3F016A17",
    x"3F016F82",
    x"3F0174EE",
    x"3F017A5A",
    x"3F017FC5",
    x"3F018531",
    x"3F018A9C",
    x"3F019007",
    x"3F019573",
    x"3F019ADE",
    x"3F01A049",
    x"3F01A5B4",
    x"3F01AB1F",
    x"3F01B08A",
    x"3F01B5F5",
    x"3F01BB5F",
    x"3F01C0CA",
    x"3F01C634",
    x"3F01CB9F",
    x"3F01D109",
    x"3F01D674",
    x"3F01DBDE",
    x"3F01E148",
    x"3F01E6B2",
    x"3F01EC1C",
    x"3F01F186",
    x"3F01F6F0",
    x"3F01FC59",
    x"3F0201C3",
    x"3F02072D",
    x"3F020C96",
    x"3F021200",
    x"3F021769",
    x"3F021CD2",
    x"3F02223C",
    x"3F0227A5",
    x"3F022D0E",
    x"3F023277",
    x"3F0237E0",
    x"3F023D48",
    x"3F0242B1",
    x"3F02481A",
    x"3F024D82",
    x"3F0252EB",
    x"3F025853",
    x"3F025DBC",
    x"3F026324",
    x"3F02688C",
    x"3F026DF4",
    x"3F02735C",
    x"3F0278C4",
    x"3F027E2C",
    x"3F028394",
    x"3F0288FC",
    x"3F028E63",
    x"3F0293CB",
    x"3F029932",
    x"3F029E9A",
    x"3F02A401",
    x"3F02A968",
    x"3F02AED0",
    x"3F02B437",
    x"3F02B99E",
    x"3F02BF05",
    x"3F02C46B",
    x"3F02C9D2",
    x"3F02CF39",
    x"3F02D49F",
    x"3F02DA06",
    x"3F02DF6C",
    x"3F02E4D3",
    x"3F02EA39",
    x"3F02EF9F",
    x"3F02F506",
    x"3F02FA6C",
    x"3F02FFD2",
    x"3F030537",
    x"3F030A9D",
    x"3F031003",
    x"3F031569",
    x"3F031ACE",
    x"3F032034",
    x"3F032599",
    x"3F032AFF",
    x"3F033064",
    x"3F0335C9",
    x"3F033B2E",
    x"3F034093",
    x"3F0345F8",
    x"3F034B5D",
    x"3F0350C2",
    x"3F035627",
    x"3F035B8B",
    x"3F0360F0",
    x"3F036654",
    x"3F036BB9",
    x"3F03711D",
    x"3F037681",
    x"3F037BE5",
    x"3F03814A",
    x"3F0386AE",
    x"3F038C11",
    x"3F039175",
    x"3F0396D9",
    x"3F039C3D",
    x"3F03A1A0",
    x"3F03A704",
    x"3F03AC67",
    x"3F03B1CB",
    x"3F03B72E",
    x"3F03BC91",
    x"3F03C1F4",
    x"3F03C757",
    x"3F03CCBA",
    x"3F03D21D",
    x"3F03D780",
    x"3F03DCE3",
    x"3F03E246",
    x"3F03E7A8",
    x"3F03ED0B",
    x"3F03F26D",
    x"3F03F7CF",
    x"3F03FD32",
    x"3F040294",
    x"3F0407F6",
    x"3F040D58",
    x"3F0412BA",
    x"3F04181C",
    x"3F041D7E",
    x"3F0422DF",
    x"3F042841",
    x"3F042DA2",
    x"3F043304",
    x"3F043865",
    x"3F043DC7",
    x"3F044328",
    x"3F044889",
    x"3F044DEA",
    x"3F04534B",
    x"3F0458AC",
    x"3F045E0D",
    x"3F04636E",
    x"3F0468CE",
    x"3F046E2F",
    x"3F04738F",
    x"3F0478F0",
    x"3F047E50",
    x"3F0483B0",
    x"3F048911",
    x"3F048E71",
    x"3F0493D1",
    x"3F049931",
    x"3F049E91",
    x"3F04A3F0",
    x"3F04A950",
    x"3F04AEB0",
    x"3F04B40F",
    x"3F04B96F",
    x"3F04BECE",
    x"3F04C42D",
    x"3F04C98D",
    x"3F04CEEC",
    x"3F04D44B",
    x"3F04D9AA",
    x"3F04DF09",
    x"3F04E468",
    x"3F04E9C6",
    x"3F04EF25",
    x"3F04F484",
    x"3F04F9E2",
    x"3F04FF41",
    x"3F05049F",
    x"3F0509FD",
    x"3F050F5B",
    x"3F0514BA",
    x"3F051A18",
    x"3F051F75",
    x"3F0524D3",
    x"3F052A31",
    x"3F052F8F",
    x"3F0534EC",
    x"3F053A4A",
    x"3F053FA8",
    x"3F054505",
    x"3F054A62",
    x"3F054FBF",
    x"3F05551D",
    x"3F055A7A",
    x"3F055FD7",
    x"3F056534",
    x"3F056A90",
    x"3F056FED",
    x"3F05754A",
    x"3F057AA6",
    x"3F058003",
    x"3F05855F",
    x"3F058ABC",
    x"3F059018",
    x"3F059574",
    x"3F059AD0",
    x"3F05A02C",
    x"3F05A588",
    x"3F05AAE4",
    x"3F05B040",
    x"3F05B59C",
    x"3F05BAF7",
    x"3F05C053",
    x"3F05C5AE",
    x"3F05CB0A",
    x"3F05D065",
    x"3F05D5C0",
    x"3F05DB1B",
    x"3F05E076",
    x"3F05E5D1",
    x"3F05EB2C",
    x"3F05F087",
    x"3F05F5E2",
    x"3F05FB3C",
    x"3F060097",
    x"3F0605F1",
    x"3F060B4C",
    x"3F0610A6",
    x"3F061600",
    x"3F061B5B",
    x"3F0620B5",
    x"3F06260F",
    x"3F062B69",
    x"3F0630C2",
    x"3F06361C",
    x"3F063B76",
    x"3F0640CF",
    x"3F064629",
    x"3F064B82",
    x"3F0650DC",
    x"3F065635",
    x"3F065B8E",
    x"3F0660E7",
    x"3F066640",
    x"3F066B99",
    x"3F0670F2",
    x"3F06764B",
    x"3F067BA4",
    x"3F0680FC",
    x"3F068655",
    x"3F068BAD",
    x"3F069106",
    x"3F06965E",
    x"3F069BB6",
    x"3F06A10E",
    x"3F06A667",
    x"3F06ABBF",
    x"3F06B116",
    x"3F06B66E",
    x"3F06BBC6",
    x"3F06C11E",
    x"3F06C675",
    x"3F06CBCD",
    x"3F06D124",
    x"3F06D67B",
    x"3F06DBD3",
    x"3F06E12A",
    x"3F06E681",
    x"3F06EBD8",
    x"3F06F12F",
    x"3F06F686",
    x"3F06FBDD",
    x"3F070133",
    x"3F07068A",
    x"3F070BE0",
    x"3F071137",
    x"3F07168D",
    x"3F071BE3",
    x"3F07213A",
    x"3F072690",
    x"3F072BE6",
    x"3F07313C",
    x"3F073692",
    x"3F073BE7",
    x"3F07413D",
    x"3F074693",
    x"3F074BE8",
    x"3F07513E",
    x"3F075693",
    x"3F075BE8",
    x"3F07613E",
    x"3F076693",
    x"3F076BE8",
    x"3F07713D",
    x"3F077692",
    x"3F077BE6",
    x"3F07813B",
    x"3F078690",
    x"3F078BE4",
    x"3F079139",
    x"3F07968D",
    x"3F079BE2",
    x"3F07A136",
    x"3F07A68A",
    x"3F07ABDE",
    x"3F07B132",
    x"3F07B686",
    x"3F07BBDA",
    x"3F07C12E",
    x"3F07C681",
    x"3F07CBD5",
    x"3F07D128",
    x"3F07D67C",
    x"3F07DBCF",
    x"3F07E122",
    x"3F07E676",
    x"3F07EBC9",
    x"3F07F11C",
    x"3F07F66F",
    x"3F07FBC1",
    x"3F080114",
    x"3F080667",
    x"3F080BB9",
    x"3F08110C",
    x"3F08165E",
    x"3F081BB1",
    x"3F082103",
    x"3F082655",
    x"3F082BA7",
    x"3F0830F9",
    x"3F08364B",
    x"3F083B9D",
    x"3F0840EF",
    x"3F084641",
    x"3F084B92",
    x"3F0850E4",
    x"3F085635",
    x"3F085B87",
    x"3F0860D8",
    x"3F086629",
    x"3F086B7A",
    x"3F0870CB",
    x"3F08761C",
    x"3F087B6D",
    x"3F0880BE",
    x"3F08860F",
    x"3F088B5F",
    x"3F0890B0",
    x"3F089600",
    x"3F089B51",
    x"3F08A0A1",
    x"3F08A5F1",
    x"3F08AB41",
    x"3F08B091",
    x"3F08B5E1",
    x"3F08BB31",
    x"3F08C081",
    x"3F08C5D1",
    x"3F08CB20",
    x"3F08D070",
    x"3F08D5BF",
    x"3F08DB0F",
    x"3F08E05E",
    x"3F08E5AD",
    x"3F08EAFD",
    x"3F08F04C",
    x"3F08F59B",
    x"3F08FAEA",
    x"3F090038",
    x"3F090587",
    x"3F090AD6",
    x"3F091024",
    x"3F091573",
    x"3F091AC1",
    x"3F092010",
    x"3F09255E",
    x"3F092AAC",
    x"3F092FFA",
    x"3F093548",
    x"3F093A96",
    x"3F093FE4",
    x"3F094531",
    x"3F094A7F",
    x"3F094FCD",
    x"3F09551A",
    x"3F095A68",
    x"3F095FB5",
    x"3F096502",
    x"3F096A4F",
    x"3F096F9C",
    x"3F0974E9",
    x"3F097A36",
    x"3F097F83",
    x"3F0984D0",
    x"3F098A1D",
    x"3F098F69",
    x"3F0994B6",
    x"3F099A02",
    x"3F099F4E",
    x"3F09A49B",
    x"3F09A9E7",
    x"3F09AF33",
    x"3F09B47F",
    x"3F09B9CB",
    x"3F09BF17",
    x"3F09C463",
    x"3F09C9AE",
    x"3F09CEFA",
    x"3F09D445",
    x"3F09D991",
    x"3F09DEDC",
    x"3F09E427",
    x"3F09E973",
    x"3F09EEBE",
    x"3F09F409",
    x"3F09F954",
    x"3F09FE9E",
    x"3F0A03E9",
    x"3F0A0934",
    x"3F0A0E7E",
    x"3F0A13C9",
    x"3F0A1913",
    x"3F0A1E5E",
    x"3F0A23A8",
    x"3F0A28F2",
    x"3F0A2E3C",
    x"3F0A3386",
    x"3F0A38D0",
    x"3F0A3E1A",
    x"3F0A4364",
    x"3F0A48AD",
    x"3F0A4DF7",
    x"3F0A5341",
    x"3F0A588A",
    x"3F0A5DD3",
    x"3F0A631D",
    x"3F0A6866",
    x"3F0A6DAF",
    x"3F0A72F8",
    x"3F0A7841",
    x"3F0A7D8A",
    x"3F0A82D2",
    x"3F0A881B",
    x"3F0A8D64",
    x"3F0A92AC",
    x"3F0A97F5",
    x"3F0A9D3D",
    x"3F0AA285",
    x"3F0AA7CD",
    x"3F0AAD16",
    x"3F0AB25E",
    x"3F0AB7A5",
    x"3F0ABCED",
    x"3F0AC235",
    x"3F0AC77D",
    x"3F0ACCC4",
    x"3F0AD20C",
    x"3F0AD753",
    x"3F0ADC9B",
    x"3F0AE1E2",
    x"3F0AE729",
    x"3F0AEC70",
    x"3F0AF1B7",
    x"3F0AF6FE",
    x"3F0AFC45",
    x"3F0B018C",
    x"3F0B06D2",
    x"3F0B0C19",
    x"3F0B115F",
    x"3F0B16A6",
    x"3F0B1BEC",
    x"3F0B2132",
    x"3F0B2679",
    x"3F0B2BBF",
    x"3F0B3105",
    x"3F0B364B",
    x"3F0B3B90",
    x"3F0B40D6",
    x"3F0B461C",
    x"3F0B4B61",
    x"3F0B50A7",
    x"3F0B55EC",
    x"3F0B5B32",
    x"3F0B6077",
    x"3F0B65BC",
    x"3F0B6B01",
    x"3F0B7046",
    x"3F0B758B",
    x"3F0B7AD0",
    x"3F0B8015",
    x"3F0B8559",
    x"3F0B8A9E",
    x"3F0B8FE2",
    x"3F0B9527",
    x"3F0B9A6B",
    x"3F0B9FAF",
    x"3F0BA4F4",
    x"3F0BAA38",
    x"3F0BAF7C",
    x"3F0BB4BF",
    x"3F0BBA03",
    x"3F0BBF47",
    x"3F0BC48B",
    x"3F0BC9CE",
    x"3F0BCF12",
    x"3F0BD455",
    x"3F0BD998",
    x"3F0BDEDC",
    x"3F0BE41F",
    x"3F0BE962",
    x"3F0BEEA5",
    x"3F0BF3E8",
    x"3F0BF92B",
    x"3F0BFE6D",
    x"3F0C03B0",
    x"3F0C08F2",
    x"3F0C0E35",
    x"3F0C1377",
    x"3F0C18BA",
    x"3F0C1DFC",
    x"3F0C233E",
    x"3F0C2880",
    x"3F0C2DC2",
    x"3F0C3304",
    x"3F0C3846",
    x"3F0C3D87",
    x"3F0C42C9",
    x"3F0C480B",
    x"3F0C4D4C",
    x"3F0C528D",
    x"3F0C57CF",
    x"3F0C5D10",
    x"3F0C6251",
    x"3F0C6792",
    x"3F0C6CD3",
    x"3F0C7214",
    x"3F0C7755",
    x"3F0C7C95",
    x"3F0C81D6",
    x"3F0C8716",
    x"3F0C8C57",
    x"3F0C9197",
    x"3F0C96D7",
    x"3F0C9C18",
    x"3F0CA158",
    x"3F0CA698",
    x"3F0CABD8",
    x"3F0CB118",
    x"3F0CB657",
    x"3F0CBB97",
    x"3F0CC0D7",
    x"3F0CC616",
    x"3F0CCB56",
    x"3F0CD095",
    x"3F0CD5D4",
    x"3F0CDB13",
    x"3F0CE052",
    x"3F0CE591",
    x"3F0CEAD0",
    x"3F0CF00F",
    x"3F0CF54E",
    x"3F0CFA8D",
    x"3F0CFFCB",
    x"3F0D050A",
    x"3F0D0A48",
    x"3F0D0F86",
    x"3F0D14C5",
    x"3F0D1A03",
    x"3F0D1F41",
    x"3F0D247F",
    x"3F0D29BD",
    x"3F0D2EFA",
    x"3F0D3438",
    x"3F0D3976",
    x"3F0D3EB3",
    x"3F0D43F1",
    x"3F0D492E",
    x"3F0D4E6C",
    x"3F0D53A9",
    x"3F0D58E6",
    x"3F0D5E23",
    x"3F0D6360",
    x"3F0D689D",
    x"3F0D6DDA",
    x"3F0D7316",
    x"3F0D7853",
    x"3F0D7D8F",
    x"3F0D82CC",
    x"3F0D8808",
    x"3F0D8D45",
    x"3F0D9281",
    x"3F0D97BD",
    x"3F0D9CF9",
    x"3F0DA235",
    x"3F0DA771",
    x"3F0DACAC",
    x"3F0DB1E8",
    x"3F0DB724",
    x"3F0DBC5F",
    x"3F0DC19B",
    x"3F0DC6D6",
    x"3F0DCC11",
    x"3F0DD14C",
    x"3F0DD687",
    x"3F0DDBC2",
    x"3F0DE0FD",
    x"3F0DE638",
    x"3F0DEB73",
    x"3F0DF0AE",
    x"3F0DF5E8",
    x"3F0DFB23",
    x"3F0E005D",
    x"3F0E0597",
    x"3F0E0AD2",
    x"3F0E100C",
    x"3F0E1546",
    x"3F0E1A80",
    x"3F0E1FBA",
    x"3F0E24F3",
    x"3F0E2A2D",
    x"3F0E2F67",
    x"3F0E34A0",
    x"3F0E39DA",
    x"3F0E3F13",
    x"3F0E444C",
    x"3F0E4986",
    x"3F0E4EBF",
    x"3F0E53F8",
    x"3F0E5931",
    x"3F0E5E6A",
    x"3F0E63A2",
    x"3F0E68DB",
    x"3F0E6E14",
    x"3F0E734C",
    x"3F0E7885",
    x"3F0E7DBD",
    x"3F0E82F5",
    x"3F0E882D",
    x"3F0E8D65",
    x"3F0E929D",
    x"3F0E97D5",
    x"3F0E9D0D",
    x"3F0EA245",
    x"3F0EA77D",
    x"3F0EACB4",
    x"3F0EB1EC",
    x"3F0EB723",
    x"3F0EBC5A",
    x"3F0EC192",
    x"3F0EC6C9",
    x"3F0ECC00",
    x"3F0ED137",
    x"3F0ED66E",
    x"3F0EDBA4",
    x"3F0EE0DB",
    x"3F0EE612",
    x"3F0EEB48",
    x"3F0EF07F",
    x"3F0EF5B5",
    x"3F0EFAEB",
    x"3F0F0022",
    x"3F0F0558",
    x"3F0F0A8E",
    x"3F0F0FC4",
    x"3F0F14FA",
    x"3F0F1A2F",
    x"3F0F1F65",
    x"3F0F249B",
    x"3F0F29D0",
    x"3F0F2F05",
    x"3F0F343B",
    x"3F0F3970",
    x"3F0F3EA5",
    x"3F0F43DA",
    x"3F0F490F",
    x"3F0F4E44",
    x"3F0F5379",
    x"3F0F58AE",
    x"3F0F5DE2",
    x"3F0F6317",
    x"3F0F684B",
    x"3F0F6D80",
    x"3F0F72B4",
    x"3F0F77E8",
    x"3F0F7D1C",
    x"3F0F8250",
    x"3F0F8784",
    x"3F0F8CB8",
    x"3F0F91EC",
    x"3F0F9720",
    x"3F0F9C53",
    x"3F0FA187",
    x"3F0FA6BA",
    x"3F0FABEE",
    x"3F0FB121",
    x"3F0FB654",
    x"3F0FBB87",
    x"3F0FC0BA",
    x"3F0FC5ED",
    x"3F0FCB20",
    x"3F0FD053",
    x"3F0FD585",
    x"3F0FDAB8",
    x"3F0FDFEA",
    x"3F0FE51D",
    x"3F0FEA4F",
    x"3F0FEF81",
    x"3F0FF4B3",
    x"3F0FF9E5",
    x"3F0FFF17",
    x"3F100449",
    x"3F10097B",
    x"3F100EAD",
    x"3F1013DE",
    x"3F101910",
    x"3F101E41",
    x"3F102373",
    x"3F1028A4",
    x"3F102DD5",
    x"3F103306",
    x"3F103837",
    x"3F103D68",
    x"3F104299",
    x"3F1047CA",
    x"3F104CFA",
    x"3F10522B",
    x"3F10575B",
    x"3F105C8C",
    x"3F1061BC",
    x"3F1066EC",
    x"3F106C1C",
    x"3F10714C",
    x"3F10767C",
    x"3F107BAC",
    x"3F1080DC",
    x"3F10860C",
    x"3F108B3B",
    x"3F10906B",
    x"3F10959A",
    x"3F109ACA",
    x"3F109FF9",
    x"3F10A528",
    x"3F10AA57",
    x"3F10AF86",
    x"3F10B4B5",
    x"3F10B9E4",
    x"3F10BF13",
    x"3F10C441",
    x"3F10C970",
    x"3F10CE9E",
    x"3F10D3CD",
    x"3F10D8FB",
    x"3F10DE29",
    x"3F10E357",
    x"3F10E885",
    x"3F10EDB3",
    x"3F10F2E1",
    x"3F10F80F",
    x"3F10FD3D",
    x"3F11026A",
    x"3F110798",
    x"3F110CC5",
    x"3F1111F3",
    x"3F111720",
    x"3F111C4D",
    x"3F11217A",
    x"3F1126A7",
    x"3F112BD4",
    x"3F113101",
    x"3F11362E",
    x"3F113B5A",
    x"3F114087",
    x"3F1145B3",
    x"3F114AE0",
    x"3F11500C",
    x"3F115538",
    x"3F115A64",
    x"3F115F90",
    x"3F1164BC",
    x"3F1169E8",
    x"3F116F14",
    x"3F117440",
    x"3F11796B",
    x"3F117E97",
    x"3F1183C2",
    x"3F1188ED",
    x"3F118E19",
    x"3F119344",
    x"3F11986F",
    x"3F119D9A",
    x"3F11A2C5",
    x"3F11A7F0",
    x"3F11AD1A",
    x"3F11B245",
    x"3F11B76F",
    x"3F11BC9A",
    x"3F11C1C4",
    x"3F11C6EF",
    x"3F11CC19",
    x"3F11D143",
    x"3F11D66D",
    x"3F11DB97",
    x"3F11E0C1",
    x"3F11E5EA",
    x"3F11EB14",
    x"3F11F03E",
    x"3F11F567",
    x"3F11FA91",
    x"3F11FFBA",
    x"3F1204E3",
    x"3F120A0C",
    x"3F120F35",
    x"3F12145E",
    x"3F121987",
    x"3F121EB0",
    x"3F1223D9",
    x"3F122901",
    x"3F122E2A",
    x"3F123352",
    x"3F12387A",
    x"3F123DA3",
    x"3F1242CB",
    x"3F1247F3",
    x"3F124D1B",
    x"3F125243",
    x"3F12576B",
    x"3F125C92",
    x"3F1261BA",
    x"3F1266E2",
    x"3F126C09",
    x"3F127130",
    x"3F127658",
    x"3F127B7F",
    x"3F1280A6",
    x"3F1285CD",
    x"3F128AF4",
    x"3F12901B",
    x"3F129542",
    x"3F129A68",
    x"3F129F8F",
    x"3F12A4B5",
    x"3F12A9DC",
    x"3F12AF02",
    x"3F12B428",
    x"3F12B94E",
    x"3F12BE74",
    x"3F12C39A",
    x"3F12C8C0",
    x"3F12CDE6",
    x"3F12D30C",
    x"3F12D831",
    x"3F12DD57",
    x"3F12E27C",
    x"3F12E7A2",
    x"3F12ECC7",
    x"3F12F1EC",
    x"3F12F711",
    x"3F12FC36",
    x"3F13015B",
    x"3F130680",
    x"3F130BA5",
    x"3F1310C9",
    x"3F1315EE",
    x"3F131B12",
    x"3F132037",
    x"3F13255B",
    x"3F132A7F",
    x"3F132FA3",
    x"3F1334C7",
    x"3F1339EB",
    x"3F133F0F",
    x"3F134433",
    x"3F134956",
    x"3F134E7A",
    x"3F13539D",
    x"3F1358C1",
    x"3F135DE4",
    x"3F136307",
    x"3F13682A",
    x"3F136D4D",
    x"3F137270",
    x"3F137793",
    x"3F137CB6",
    x"3F1381D9",
    x"3F1386FB",
    x"3F138C1E",
    x"3F139140",
    x"3F139663",
    x"3F139B85",
    x"3F13A0A7",
    x"3F13A5C9",
    x"3F13AAEB",
    x"3F13B00D",
    x"3F13B52F",
    x"3F13BA50",
    x"3F13BF72",
    x"3F13C493",
    x"3F13C9B5",
    x"3F13CED6",
    x"3F13D3F8",
    x"3F13D919",
    x"3F13DE3A",
    x"3F13E35B",
    x"3F13E87C",
    x"3F13ED9C",
    x"3F13F2BD",
    x"3F13F7DE",
    x"3F13FCFE",
    x"3F14021F",
    x"3F14073F",
    x"3F140C5F",
    x"3F141180",
    x"3F1416A0",
    x"3F141BC0",
    x"3F1420E0",
    x"3F142600",
    x"3F142B1F",
    x"3F14303F",
    x"3F14355E",
    x"3F143A7E",
    x"3F143F9D",
    x"3F1444BD",
    x"3F1449DC",
    x"3F144EFB",
    x"3F14541A",
    x"3F145939",
    x"3F145E58",
    x"3F146377",
    x"3F146895",
    x"3F146DB4",
    x"3F1472D2",
    x"3F1477F1",
    x"3F147D0F",
    x"3F14822D",
    x"3F14874B",
    x"3F148C69",
    x"3F149187",
    x"3F1496A5",
    x"3F149BC3",
    x"3F14A0E1",
    x"3F14A5FE",
    x"3F14AB1C",
    x"3F14B039",
    x"3F14B557",
    x"3F14BA74",
    x"3F14BF91",
    x"3F14C4AE",
    x"3F14C9CB",
    x"3F14CEE8",
    x"3F14D405",
    x"3F14D921",
    x"3F14DE3E",
    x"3F14E35A",
    x"3F14E877",
    x"3F14ED93",
    x"3F14F2B0",
    x"3F14F7CC",
    x"3F14FCE8",
    x"3F150204",
    x"3F150720",
    x"3F150C3B",
    x"3F151157",
    x"3F151673",
    x"3F151B8E",
    x"3F1520AA",
    x"3F1525C5",
    x"3F152AE0",
    x"3F152FFC",
    x"3F153517",
    x"3F153A32",
    x"3F153F4D",
    x"3F154467",
    x"3F154982",
    x"3F154E9D",
    x"3F1553B7",
    x"3F1558D2",
    x"3F155DEC",
    x"3F156306",
    x"3F156821",
    x"3F156D3B",
    x"3F157255",
    x"3F15776F",
    x"3F157C88",
    x"3F1581A2",
    x"3F1586BC",
    x"3F158BD5",
    x"3F1590EF",
    x"3F159608",
    x"3F159B21",
    x"3F15A03B",
    x"3F15A554",
    x"3F15AA6D",
    x"3F15AF86",
    x"3F15B49F",
    x"3F15B9B7",
    x"3F15BED0",
    x"3F15C3E9",
    x"3F15C901",
    x"3F15CE19",
    x"3F15D332",
    x"3F15D84A",
    x"3F15DD62",
    x"3F15E27A",
    x"3F15E792",
    x"3F15ECAA",
    x"3F15F1C2",
    x"3F15F6D9",
    x"3F15FBF1",
    x"3F160108",
    x"3F160620",
    x"3F160B37",
    x"3F16104E",
    x"3F161565",
    x"3F161A7C",
    x"3F161F93",
    x"3F1624AA",
    x"3F1629C1",
    x"3F162ED8",
    x"3F1633EE",
    x"3F163905",
    x"3F163E1B",
    x"3F164331",
    x"3F164847",
    x"3F164D5E",
    x"3F165274",
    x"3F16578A",
    x"3F165C9F",
    x"3F1661B5",
    x"3F1666CB",
    x"3F166BE0",
    x"3F1670F6",
    x"3F16760B",
    x"3F167B21",
    x"3F168036",
    x"3F16854B",
    x"3F168A60",
    x"3F168F75",
    x"3F16948A",
    x"3F16999F",
    x"3F169EB3",
    x"3F16A3C8",
    x"3F16A8DC",
    x"3F16ADF1",
    x"3F16B305",
    x"3F16B819",
    x"3F16BD2D",
    x"3F16C241",
    x"3F16C755",
    x"3F16CC69",
    x"3F16D17D",
    x"3F16D691",
    x"3F16DBA4",
    x"3F16E0B8",
    x"3F16E5CB",
    x"3F16EADE",
    x"3F16EFF2",
    x"3F16F505",
    x"3F16FA18",
    x"3F16FF2B",
    x"3F17043E",
    x"3F170950",
    x"3F170E63",
    x"3F171376",
    x"3F171888",
    x"3F171D9B",
    x"3F1722AD",
    x"3F1727BF",
    x"3F172CD1",
    x"3F1731E3",
    x"3F1736F5",
    x"3F173C07",
    x"3F174119",
    x"3F17462B",
    x"3F174B3C",
    x"3F17504E",
    x"3F17555F",
    x"3F175A70",
    x"3F175F82",
    x"3F176493",
    x"3F1769A4",
    x"3F176EB5",
    x"3F1773C6",
    x"3F1778D6",
    x"3F177DE7",
    x"3F1782F8",
    x"3F178808",
    x"3F178D18",
    x"3F179229",
    x"3F179739",
    x"3F179C49",
    x"3F17A159",
    x"3F17A669",
    x"3F17AB79",
    x"3F17B089",
    x"3F17B598",
    x"3F17BAA8",
    x"3F17BFB7",
    x"3F17C4C7",
    x"3F17C9D6",
    x"3F17CEE5",
    x"3F17D3F4",
    x"3F17D903",
    x"3F17DE12",
    x"3F17E321",
    x"3F17E830",
    x"3F17ED3F",
    x"3F17F24D",
    x"3F17F75C",
    x"3F17FC6A",
    x"3F180178",
    x"3F180687",
    x"3F180B95",
    x"3F1810A3",
    x"3F1815B1",
    x"3F181ABE",
    x"3F181FCC",
    x"3F1824DA",
    x"3F1829E7",
    x"3F182EF5",
    x"3F183402",
    x"3F183910",
    x"3F183E1D",
    x"3F18432A",
    x"3F184837",
    x"3F184D44",
    x"3F185251",
    x"3F18575D",
    x"3F185C6A",
    x"3F186177",
    x"3F186683",
    x"3F186B8F",
    x"3F18709C",
    x"3F1875A8",
    x"3F187AB4",
    x"3F187FC0",
    x"3F1884CC",
    x"3F1889D8",
    x"3F188EE3",
    x"3F1893EF",
    x"3F1898FB",
    x"3F189E06",
    x"3F18A311",
    x"3F18A81D",
    x"3F18AD28",
    x"3F18B233",
    x"3F18B73E",
    x"3F18BC49",
    x"3F18C154",
    x"3F18C65E",
    x"3F18CB69",
    x"3F18D073",
    x"3F18D57E",
    x"3F18DA88",
    x"3F18DF92",
    x"3F18E49D",
    x"3F18E9A7",
    x"3F18EEB1",
    x"3F18F3BB",
    x"3F18F8C4",
    x"3F18FDCE",
    x"3F1902D8",
    x"3F1907E1",
    x"3F190CEB",
    x"3F1911F4",
    x"3F1916FD",
    x"3F191C06",
    x"3F19210F",
    x"3F192618",
    x"3F192B21",
    x"3F19302A",
    x"3F193533",
    x"3F193A3B",
    x"3F193F44",
    x"3F19444C",
    x"3F194955",
    x"3F194E5D",
    x"3F195365",
    x"3F19586D",
    x"3F195D75",
    x"3F19627D",
    x"3F196784",
    x"3F196C8C",
    x"3F197194",
    x"3F19769B",
    x"3F197BA3",
    x"3F1980AA",
    x"3F1985B1",
    x"3F198AB8",
    x"3F198FBF",
    x"3F1994C6",
    x"3F1999CD",
    x"3F199ED4",
    x"3F19A3DA",
    x"3F19A8E1",
    x"3F19ADE7",
    x"3F19B2EE",
    x"3F19B7F4",
    x"3F19BCFA",
    x"3F19C200",
    x"3F19C706",
    x"3F19CC0C",
    x"3F19D112",
    x"3F19D618",
    x"3F19DB1E",
    x"3F19E023",
    x"3F19E529",
    x"3F19EA2E",
    x"3F19EF33",
    x"3F19F438",
    x"3F19F93D",
    x"3F19FE42",
    x"3F1A0347",
    x"3F1A084C",
    x"3F1A0D51",
    x"3F1A1255",
    x"3F1A175A",
    x"3F1A1C5E",
    x"3F1A2163",
    x"3F1A2667",
    x"3F1A2B6B",
    x"3F1A306F",
    x"3F1A3573",
    x"3F1A3A77",
    x"3F1A3F7B",
    x"3F1A447E",
    x"3F1A4982",
    x"3F1A4E86",
    x"3F1A5389",
    x"3F1A588C",
    x"3F1A5D8F",
    x"3F1A6293",
    x"3F1A6796",
    x"3F1A6C99",
    x"3F1A719B",
    x"3F1A769E",
    x"3F1A7BA1",
    x"3F1A80A3",
    x"3F1A85A6",
    x"3F1A8AA8",
    x"3F1A8FAB",
    x"3F1A94AD",
    x"3F1A99AF",
    x"3F1A9EB1",
    x"3F1AA3B3",
    x"3F1AA8B5",
    x"3F1AADB6",
    x"3F1AB2B8",
    x"3F1AB7BA",
    x"3F1ABCBB",
    x"3F1AC1BC",
    x"3F1AC6BE",
    x"3F1ACBBF",
    x"3F1AD0C0",
    x"3F1AD5C1",
    x"3F1ADAC2",
    x"3F1ADFC3",
    x"3F1AE4C3",
    x"3F1AE9C4",
    x"3F1AEEC4",
    x"3F1AF3C5",
    x"3F1AF8C5",
    x"3F1AFDC5",
    x"3F1B02C6",
    x"3F1B07C6",
    x"3F1B0CC6",
    x"3F1B11C5",
    x"3F1B16C5",
    x"3F1B1BC5",
    x"3F1B20C4",
    x"3F1B25C4",
    x"3F1B2AC3",
    x"3F1B2FC3",
    x"3F1B34C2",
    x"3F1B39C1",
    x"3F1B3EC0",
    x"3F1B43BF",
    x"3F1B48BE",
    x"3F1B4DBD",
    x"3F1B52BB",
    x"3F1B57BA",
    x"3F1B5CB8",
    x"3F1B61B7",
    x"3F1B66B5",
    x"3F1B6BB3",
    x"3F1B70B1",
    x"3F1B75AF",
    x"3F1B7AAD",
    x"3F1B7FAB",
    x"3F1B84A9",
    x"3F1B89A6",
    x"3F1B8EA4",
    x"3F1B93A1",
    x"3F1B989E",
    x"3F1B9D9C",
    x"3F1BA299",
    x"3F1BA796",
    x"3F1BAC93",
    x"3F1BB190",
    x"3F1BB68D",
    x"3F1BBB89",
    x"3F1BC086",
    x"3F1BC582",
    x"3F1BCA7F",
    x"3F1BCF7B",
    x"3F1BD477",
    x"3F1BD973",
    x"3F1BDE6F",
    x"3F1BE36B",
    x"3F1BE867",
    x"3F1BED63",
    x"3F1BF25F",
    x"3F1BF75A",
    x"3F1BFC56",
    x"3F1C0151",
    x"3F1C064C",
    x"3F1C0B47",
    x"3F1C1042",
    x"3F1C153D",
    x"3F1C1A38",
    x"3F1C1F33",
    x"3F1C242E",
    x"3F1C2929",
    x"3F1C2E23",
    x"3F1C331D",
    x"3F1C3818",
    x"3F1C3D12",
    x"3F1C420C",
    x"3F1C4706",
    x"3F1C4C00",
    x"3F1C50FA",
    x"3F1C55F4",
    x"3F1C5AEE",
    x"3F1C5FE7",
    x"3F1C64E1",
    x"3F1C69DA",
    x"3F1C6ED3",
    x"3F1C73CC",
    x"3F1C78C6",
    x"3F1C7DBF",
    x"3F1C82B8",
    x"3F1C87B0",
    x"3F1C8CA9",
    x"3F1C91A2",
    x"3F1C969A",
    x"3F1C9B93",
    x"3F1CA08B",
    x"3F1CA583",
    x"3F1CAA7C",
    x"3F1CAF74",
    x"3F1CB46C",
    x"3F1CB963",
    x"3F1CBE5B",
    x"3F1CC353",
    x"3F1CC84B",
    x"3F1CCD42",
    x"3F1CD239",
    x"3F1CD731",
    x"3F1CDC28",
    x"3F1CE11F",
    x"3F1CE616",
    x"3F1CEB0D",
    x"3F1CF004",
    x"3F1CF4FB",
    x"3F1CF9F1",
    x"3F1CFEE8",
    x"3F1D03DE",
    x"3F1D08D5",
    x"3F1D0DCB",
    x"3F1D12C1",
    x"3F1D17B7",
    x"3F1D1CAD",
    x"3F1D21A3",
    x"3F1D2699",
    x"3F1D2B8F",
    x"3F1D3084",
    x"3F1D357A",
    x"3F1D3A6F",
    x"3F1D3F65",
    x"3F1D445A",
    x"3F1D494F",
    x"3F1D4E44",
    x"3F1D5339",
    x"3F1D582E",
    x"3F1D5D23",
    x"3F1D6217",
    x"3F1D670C",
    x"3F1D6C00",
    x"3F1D70F5",
    x"3F1D75E9",
    x"3F1D7ADD",
    x"3F1D7FD1",
    x"3F1D84C5",
    x"3F1D89B9",
    x"3F1D8EAD",
    x"3F1D93A1",
    x"3F1D9894",
    x"3F1D9D88",
    x"3F1DA27B",
    x"3F1DA76F",
    x"3F1DAC62",
    x"3F1DB155",
    x"3F1DB648",
    x"3F1DBB3B",
    x"3F1DC02E",
    x"3F1DC521",
    x"3F1DCA13",
    x"3F1DCF06",
    x"3F1DD3F8",
    x"3F1DD8EB",
    x"3F1DDDDD",
    x"3F1DE2CF",
    x"3F1DE7C1",
    x"3F1DECB3",
    x"3F1DF1A5",
    x"3F1DF697",
    x"3F1DFB89",
    x"3F1E007B",
    x"3F1E056C",
    x"3F1E0A5D",
    x"3F1E0F4F",
    x"3F1E1440",
    x"3F1E1931",
    x"3F1E1E22",
    x"3F1E2313",
    x"3F1E2804",
    x"3F1E2CF5",
    x"3F1E31E6",
    x"3F1E36D6",
    x"3F1E3BC7",
    x"3F1E40B7",
    x"3F1E45A7",
    x"3F1E4A98",
    x"3F1E4F88",
    x"3F1E5478",
    x"3F1E5968",
    x"3F1E5E57",
    x"3F1E6347",
    x"3F1E6837",
    x"3F1E6D26",
    x"3F1E7216",
    x"3F1E7705",
    x"3F1E7BF4",
    x"3F1E80E3",
    x"3F1E85D2",
    x"3F1E8AC1",
    x"3F1E8FB0",
    x"3F1E949F",
    x"3F1E998E",
    x"3F1E9E7C",
    x"3F1EA36B",
    x"3F1EA859",
    x"3F1EAD47",
    x"3F1EB236",
    x"3F1EB724",
    x"3F1EBC12",
    x"3F1EC100",
    x"3F1EC5ED",
    x"3F1ECADB",
    x"3F1ECFC9",
    x"3F1ED4B6",
    x"3F1ED9A4",
    x"3F1EDE91",
    x"3F1EE37E",
    x"3F1EE86C",
    x"3F1EED59",
    x"3F1EF245",
    x"3F1EF732",
    x"3F1EFC1F",
    x"3F1F010C",
    x"3F1F05F8",
    x"3F1F0AE5",
    x"3F1F0FD1",
    x"3F1F14BD",
    x"3F1F19AA",
    x"3F1F1E96",
    x"3F1F2382",
    x"3F1F286E",
    x"3F1F2D59",
    x"3F1F3245",
    x"3F1F3731",
    x"3F1F3C1C",
    x"3F1F4108",
    x"3F1F45F3",
    x"3F1F4ADE",
    x"3F1F4FC9",
    x"3F1F54B4",
    x"3F1F599F",
    x"3F1F5E8A",
    x"3F1F6375",
    x"3F1F6860",
    x"3F1F6D4A",
    x"3F1F7235",
    x"3F1F771F",
    x"3F1F7C09",
    x"3F1F80F3",
    x"3F1F85DD",
    x"3F1F8AC7",
    x"3F1F8FB1",
    x"3F1F949B",
    x"3F1F9985",
    x"3F1F9E6E",
    x"3F1FA358",
    x"3F1FA841",
    x"3F1FAD2B",
    x"3F1FB214",
    x"3F1FB6FD",
    x"3F1FBBE6",
    x"3F1FC0CF",
    x"3F1FC5B8",
    x"3F1FCAA0",
    x"3F1FCF89",
    x"3F1FD472",
    x"3F1FD95A",
    x"3F1FDE42",
    x"3F1FE32B",
    x"3F1FE813",
    x"3F1FECFB",
    x"3F1FF1E3",
    x"3F1FF6CB",
    x"3F1FFBB2",
    x"3F20009A",
    x"3F200582",
    x"3F200A69",
    x"3F200F50",
    x"3F201438",
    x"3F20191F",
    x"3F201E06",
    x"3F2022ED",
    x"3F2027D4",
    x"3F202CBB",
    x"3F2031A1",
    x"3F203688",
    x"3F203B6F",
    x"3F204055",
    x"3F20453B",
    x"3F204A21",
    x"3F204F08",
    x"3F2053EE",
    x"3F2058D4",
    x"3F205DB9",
    x"3F20629F",
    x"3F206785",
    x"3F206C6A",
    x"3F207150",
    x"3F207635",
    x"3F207B1A",
    x"3F208000",
    x"3F2084E5",
    x"3F2089CA",
    x"3F208EAE",
    x"3F209393",
    x"3F209878",
    x"3F209D5C",
    x"3F20A241",
    x"3F20A725",
    x"3F20AC0A",
    x"3F20B0EE",
    x"3F20B5D2",
    x"3F20BAB6",
    x"3F20BF9A",
    x"3F20C47E",
    x"3F20C961",
    x"3F20CE45",
    x"3F20D328",
    x"3F20D80C",
    x"3F20DCEF",
    x"3F20E1D2",
    x"3F20E6B5",
    x"3F20EB99",
    x"3F20F07B",
    x"3F20F55E",
    x"3F20FA41",
    x"3F20FF24",
    x"3F210406",
    x"3F2108E9",
    x"3F210DCB",
    x"3F2112AD",
    x"3F21178F",
    x"3F211C71",
    x"3F212153",
    x"3F212635",
    x"3F212B17",
    x"3F212FF9",
    x"3F2134DA",
    x"3F2139BC",
    x"3F213E9D",
    x"3F21437E",
    x"3F214860",
    x"3F214D41",
    x"3F215222",
    x"3F215703",
    x"3F215BE3",
    x"3F2160C4",
    x"3F2165A5",
    x"3F216A85",
    x"3F216F66",
    x"3F217446",
    x"3F217926",
    x"3F217E06",
    x"3F2182E6",
    x"3F2187C6",
    x"3F218CA6",
    x"3F219186",
    x"3F219665",
    x"3F219B45",
    x"3F21A024",
    x"3F21A504",
    x"3F21A9E3",
    x"3F21AEC2",
    x"3F21B3A1",
    x"3F21B880",
    x"3F21BD5F",
    x"3F21C23E",
    x"3F21C71C",
    x"3F21CBFB",
    x"3F21D0D9",
    x"3F21D5B8",
    x"3F21DA96",
    x"3F21DF74",
    x"3F21E452",
    x"3F21E930",
    x"3F21EE0E",
    x"3F21F2EC",
    x"3F21F7C9",
    x"3F21FCA7",
    x"3F220185",
    x"3F220662",
    x"3F220B3F",
    x"3F22101C",
    x"3F2214FA",
    x"3F2219D7",
    x"3F221EB3",
    x"3F222390",
    x"3F22286D",
    x"3F222D4A",
    x"3F223226",
    x"3F223702",
    x"3F223BDF",
    x"3F2240BB",
    x"3F224597",
    x"3F224A73",
    x"3F224F4F",
    x"3F22542B",
    x"3F225907",
    x"3F225DE2",
    x"3F2262BE",
    x"3F226799",
    x"3F226C74",
    x"3F227150",
    x"3F22762B",
    x"3F227B06",
    x"3F227FE1",
    x"3F2284BC",
    x"3F228996",
    x"3F228E71",
    x"3F22934C",
    x"3F229826",
    x"3F229D00",
    x"3F22A1DB",
    x"3F22A6B5",
    x"3F22AB8F",
    x"3F22B069",
    x"3F22B543",
    x"3F22BA1D",
    x"3F22BEF6",
    x"3F22C3D0",
    x"3F22C8A9",
    x"3F22CD83",
    x"3F22D25C",
    x"3F22D735",
    x"3F22DC0E",
    x"3F22E0E7",
    x"3F22E5C0",
    x"3F22EA99",
    x"3F22EF72",
    x"3F22F44A",
    x"3F22F923",
    x"3F22FDFB",
    x"3F2302D3",
    x"3F2307AB",
    x"3F230C84",
    x"3F23115C",
    x"3F231633",
    x"3F231B0B",
    x"3F231FE3",
    x"3F2324BB",
    x"3F232992",
    x"3F232E6A",
    x"3F233341",
    x"3F233818",
    x"3F233CEF",
    x"3F2341C6",
    x"3F23469D",
    x"3F234B74",
    x"3F23504B",
    x"3F235521",
    x"3F2359F8",
    x"3F235ECE",
    x"3F2363A5",
    x"3F23687B",
    x"3F236D51",
    x"3F237227",
    x"3F2376FD",
    x"3F237BD3",
    x"3F2380A8",
    x"3F23857E",
    x"3F238A54",
    x"3F238F29",
    x"3F2393FE",
    x"3F2398D4",
    x"3F239DA9",
    x"3F23A27E",
    x"3F23A753",
    x"3F23AC28",
    x"3F23B0FC",
    x"3F23B5D1",
    x"3F23BAA6",
    x"3F23BF7A",
    x"3F23C44F",
    x"3F23C923",
    x"3F23CDF7",
    x"3F23D2CB",
    x"3F23D79F",
    x"3F23DC73",
    x"3F23E147",
    x"3F23E61A",
    x"3F23EAEE",
    x"3F23EFC1",
    x"3F23F495",
    x"3F23F968",
    x"3F23FE3B",
    x"3F24030E",
    x"3F2407E1",
    x"3F240CB4",
    x"3F241187",
    x"3F24165A",
    x"3F241B2C",
    x"3F241FFF",
    x"3F2424D1",
    x"3F2429A3",
    x"3F242E75",
    x"3F243348",
    x"3F24381A",
    x"3F243CEB",
    x"3F2441BD",
    x"3F24468F",
    x"3F244B60",
    x"3F245032",
    x"3F245503",
    x"3F2459D5",
    x"3F245EA6",
    x"3F246377",
    x"3F246848",
    x"3F246D19",
    x"3F2471EA",
    x"3F2476BA",
    x"3F247B8B",
    x"3F24805B",
    x"3F24852C",
    x"3F2489FC",
    x"3F248ECC",
    x"3F24939C",
    x"3F24986D",
    x"3F249D3C",
    x"3F24A20C",
    x"3F24A6DC",
    x"3F24ABAC",
    x"3F24B07B",
    x"3F24B54A",
    x"3F24BA1A",
    x"3F24BEE9",
    x"3F24C3B8",
    x"3F24C887",
    x"3F24CD56",
    x"3F24D225",
    x"3F24D6F4",
    x"3F24DBC2",
    x"3F24E091",
    x"3F24E55F",
    x"3F24EA2D",
    x"3F24EEFC",
    x"3F24F3CA",
    x"3F24F898",
    x"3F24FD66",
    x"3F250234",
    x"3F250701",
    x"3F250BCF",
    x"3F25109C",
    x"3F25156A",
    x"3F251A37",
    x"3F251F04",
    x"3F2523D2",
    x"3F25289F",
    x"3F252D6C",
    x"3F253238",
    x"3F253705",
    x"3F253BD2",
    x"3F25409E",
    x"3F25456B",
    x"3F254A37",
    x"3F254F03",
    x"3F2553CF",
    x"3F25589B",
    x"3F255D67",
    x"3F256233",
    x"3F2566FF",
    x"3F256BCB",
    x"3F257096",
    x"3F257562",
    x"3F257A2D",
    x"3F257EF8",
    x"3F2583C3",
    x"3F25888E",
    x"3F258D59",
    x"3F259224",
    x"3F2596EF",
    x"3F259BB9",
    x"3F25A084",
    x"3F25A54E",
    x"3F25AA19",
    x"3F25AEE3",
    x"3F25B3AD",
    x"3F25B877",
    x"3F25BD41",
    x"3F25C20B",
    x"3F25C6D5",
    x"3F25CB9E",
    x"3F25D068",
    x"3F25D531",
    x"3F25D9FB",
    x"3F25DEC4",
    x"3F25E38D",
    x"3F25E856",
    x"3F25ED1F",
    x"3F25F1E8",
    x"3F25F6B1",
    x"3F25FB79",
    x"3F260042",
    x"3F26050A",
    x"3F2609D3",
    x"3F260E9B",
    x"3F261363",
    x"3F26182B",
    x"3F261CF3",
    x"3F2621BB",
    x"3F262682",
    x"3F262B4A",
    x"3F263012",
    x"3F2634D9",
    x"3F2639A0",
    x"3F263E68",
    x"3F26432F",
    x"3F2647F6",
    x"3F264CBD",
    x"3F265184",
    x"3F26564A",
    x"3F265B11",
    x"3F265FD8",
    x"3F26649E",
    x"3F266964",
    x"3F266E2B",
    x"3F2672F1",
    x"3F2677B7",
    x"3F267C7D",
    x"3F268143",
    x"3F268608",
    x"3F268ACE",
    x"3F268F93",
    x"3F269459",
    x"3F26991E",
    x"3F269DE3",
    x"3F26A2A9",
    x"3F26A76E",
    x"3F26AC33",
    x"3F26B0F7",
    x"3F26B5BC",
    x"3F26BA81",
    x"3F26BF45",
    x"3F26C40A",
    x"3F26C8CE",
    x"3F26CD92",
    x"3F26D256",
    x"3F26D71A",
    x"3F26DBDE",
    x"3F26E0A2",
    x"3F26E566",
    x"3F26EA2A",
    x"3F26EEED",
    x"3F26F3B0",
    x"3F26F874",
    x"3F26FD37",
    x"3F2701FA",
    x"3F2706BD",
    x"3F270B80",
    x"3F271043",
    x"3F271506",
    x"3F2719C8",
    x"3F271E8B",
    x"3F27234D",
    x"3F272810",
    x"3F272CD2",
    x"3F273194",
    x"3F273656",
    x"3F273B18",
    x"3F273FDA",
    x"3F27449B",
    x"3F27495D",
    x"3F274E1E",
    x"3F2752E0",
    x"3F2757A1",
    x"3F275C62",
    x"3F276123",
    x"3F2765E5",
    x"3F276AA5",
    x"3F276F66",
    x"3F277427",
    x"3F2778E8",
    x"3F277DA8",
    x"3F278268",
    x"3F278729",
    x"3F278BE9",
    x"3F2790A9",
    x"3F279569",
    x"3F279A29",
    x"3F279EE9",
    x"3F27A3A8",
    x"3F27A868",
    x"3F27AD28",
    x"3F27B1E7",
    x"3F27B6A6",
    x"3F27BB65",
    x"3F27C025",
    x"3F27C4E4",
    x"3F27C9A2",
    x"3F27CE61",
    x"3F27D320",
    x"3F27D7DE",
    x"3F27DC9D",
    x"3F27E15B",
    x"3F27E61A",
    x"3F27EAD8",
    x"3F27EF96",
    x"3F27F454",
    x"3F27F912",
    x"3F27FDD0",
    x"3F28028D",
    x"3F28074B",
    x"3F280C08",
    x"3F2810C6",
    x"3F281583",
    x"3F281A40",
    x"3F281EFD",
    x"3F2823BA",
    x"3F282877",
    x"3F282D34",
    x"3F2831F0",
    x"3F2836AD",
    x"3F283B69",
    x"3F284026",
    x"3F2844E2",
    x"3F28499E",
    x"3F284E5A",
    x"3F285316",
    x"3F2857D2",
    x"3F285C8E",
    x"3F286149",
    x"3F286605",
    x"3F286AC0",
    x"3F286F7C",
    x"3F287437",
    x"3F2878F2",
    x"3F287DAD",
    x"3F288268",
    x"3F288723",
    x"3F288BDE",
    x"3F289098",
    x"3F289553",
    x"3F289A0D",
    x"3F289EC8",
    x"3F28A382",
    x"3F28A83C",
    x"3F28ACF6",
    x"3F28B1B0",
    x"3F28B66A",
    x"3F28BB23",
    x"3F28BFDD",
    x"3F28C497",
    x"3F28C950",
    x"3F28CE09",
    x"3F28D2C3",
    x"3F28D77C",
    x"3F28DC35",
    x"3F28E0EE",
    x"3F28E5A6",
    x"3F28EA5F",
    x"3F28EF18",
    x"3F28F3D0",
    x"3F28F889",
    x"3F28FD41",
    x"3F2901F9",
    x"3F2906B1",
    x"3F290B69",
    x"3F291021",
    x"3F2914D9",
    x"3F291991",
    x"3F291E48",
    x"3F292300",
    x"3F2927B7",
    x"3F292C6E",
    x"3F293125",
    x"3F2935DD",
    x"3F293A93",
    x"3F293F4A",
    x"3F294401",
    x"3F2948B8",
    x"3F294D6E",
    x"3F295225",
    x"3F2956DB",
    x"3F295B91",
    x"3F296048",
    x"3F2964FE",
    x"3F2969B4",
    x"3F296E69",
    x"3F29731F",
    x"3F2977D5",
    x"3F297C8A",
    x"3F298140",
    x"3F2985F5",
    x"3F298AAA",
    x"3F298F60",
    x"3F299415",
    x"3F2998CA",
    x"3F299D7E",
    x"3F29A233",
    x"3F29A6E8",
    x"3F29AB9C",
    x"3F29B051",
    x"3F29B505",
    x"3F29B9B9",
    x"3F29BE6D",
    x"3F29C321",
    x"3F29C7D5",
    x"3F29CC89",
    x"3F29D13D",
    x"3F29D5F0",
    x"3F29DAA4",
    x"3F29DF57",
    x"3F29E40B",
    x"3F29E8BE",
    x"3F29ED71",
    x"3F29F224",
    x"3F29F6D7",
    x"3F29FB89",
    x"3F2A003C",
    x"3F2A04EF",
    x"3F2A09A1",
    x"3F2A0E54",
    x"3F2A1306",
    x"3F2A17B8",
    x"3F2A1C6A",
    x"3F2A211C",
    x"3F2A25CE",
    x"3F2A2A80",
    x"3F2A2F31",
    x"3F2A33E3",
    x"3F2A3894",
    x"3F2A3D46",
    x"3F2A41F7",
    x"3F2A46A8",
    x"3F2A4B59",
    x"3F2A500A",
    x"3F2A54BB",
    x"3F2A596C",
    x"3F2A5E1C",
    x"3F2A62CD",
    x"3F2A677D",
    x"3F2A6C2E",
    x"3F2A70DE",
    x"3F2A758E",
    x"3F2A7A3E",
    x"3F2A7EEE",
    x"3F2A839E",
    x"3F2A884D",
    x"3F2A8CFD",
    x"3F2A91AC",
    x"3F2A965C",
    x"3F2A9B0B",
    x"3F2A9FBA",
    x"3F2AA469",
    x"3F2AA918",
    x"3F2AADC7",
    x"3F2AB276",
    x"3F2AB725",
    x"3F2ABBD3",
    x"3F2AC082",
    x"3F2AC530",
    x"3F2AC9DE",
    x"3F2ACE8D",
    x"3F2AD33B",
    x"3F2AD7E9",
    x"3F2ADC96",
    x"3F2AE144",
    x"3F2AE5F2",
    x"3F2AEA9F",
    x"3F2AEF4D",
    x"3F2AF3FA",
    x"3F2AF8A7",
    x"3F2AFD55",
    x"3F2B0202",
    x"3F2B06AF",
    x"3F2B0B5B",
    x"3F2B1008",
    x"3F2B14B5",
    x"3F2B1961",
    x"3F2B1E0E",
    x"3F2B22BA",
    x"3F2B2766",
    x"3F2B2C12",
    x"3F2B30BE",
    x"3F2B356A",
    x"3F2B3A16",
    x"3F2B3EC2",
    x"3F2B436D",
    x"3F2B4819",
    x"3F2B4CC4",
    x"3F2B516F",
    x"3F2B561B",
    x"3F2B5AC6",
    x"3F2B5F71",
    x"3F2B641B",
    x"3F2B68C6",
    x"3F2B6D71",
    x"3F2B721B",
    x"3F2B76C6",
    x"3F2B7B70",
    x"3F2B801A",
    x"3F2B84C5",
    x"3F2B896F",
    x"3F2B8E19",
    x"3F2B92C2",
    x"3F2B976C",
    x"3F2B9C16",
    x"3F2BA0BF",
    x"3F2BA569",
    x"3F2BAA12",
    x"3F2BAEBB",
    x"3F2BB364",
    x"3F2BB80D",
    x"3F2BBCB6",
    x"3F2BC15F",
    x"3F2BC608",
    x"3F2BCAB0",
    x"3F2BCF59",
    x"3F2BD401",
    x"3F2BD8AA",
    x"3F2BDD52",
    x"3F2BE1FA",
    x"3F2BE6A2",
    x"3F2BEB4A",
    x"3F2BEFF1",
    x"3F2BF499",
    x"3F2BF941",
    x"3F2BFDE8",
    x"3F2C028F",
    x"3F2C0737",
    x"3F2C0BDE",
    x"3F2C1085",
    x"3F2C152C",
    x"3F2C19D3",
    x"3F2C1E79",
    x"3F2C2320",
    x"3F2C27C7",
    x"3F2C2C6D",
    x"3F2C3113",
    x"3F2C35B9",
    x"3F2C3A60",
    x"3F2C3F06",
    x"3F2C43AB",
    x"3F2C4851",
    x"3F2C4CF7",
    x"3F2C519D",
    x"3F2C5642",
    x"3F2C5AE7",
    x"3F2C5F8D",
    x"3F2C6432",
    x"3F2C68D7",
    x"3F2C6D7C",
    x"3F2C7221",
    x"3F2C76C5",
    x"3F2C7B6A",
    x"3F2C800F",
    x"3F2C84B3",
    x"3F2C8957",
    x"3F2C8DFC",
    x"3F2C92A0",
    x"3F2C9744",
    x"3F2C9BE8",
    x"3F2CA08C",
    x"3F2CA52F",
    x"3F2CA9D3",
    x"3F2CAE76",
    x"3F2CB31A",
    x"3F2CB7BD",
    x"3F2CBC60",
    x"3F2CC103",
    x"3F2CC5A6",
    x"3F2CCA49",
    x"3F2CCEEC",
    x"3F2CD38F",
    x"3F2CD831",
    x"3F2CDCD4",
    x"3F2CE176",
    x"3F2CE618",
    x"3F2CEABB",
    x"3F2CEF5D",
    x"3F2CF3FF",
    x"3F2CF8A0",
    x"3F2CFD42",
    x"3F2D01E4",
    x"3F2D0685",
    x"3F2D0B27",
    x"3F2D0FC8",
    x"3F2D1469",
    x"3F2D190A",
    x"3F2D1DAB",
    x"3F2D224C",
    x"3F2D26ED",
    x"3F2D2B8E",
    x"3F2D302E",
    x"3F2D34CF",
    x"3F2D396F",
    x"3F2D3E10",
    x"3F2D42B0",
    x"3F2D4750",
    x"3F2D4BF0",
    x"3F2D5090",
    x"3F2D552F",
    x"3F2D59CF",
    x"3F2D5E6F",
    x"3F2D630E",
    x"3F2D67AD",
    x"3F2D6C4D",
    x"3F2D70EC",
    x"3F2D758B",
    x"3F2D7A2A",
    x"3F2D7EC9",
    x"3F2D8367",
    x"3F2D8806",
    x"3F2D8CA4",
    x"3F2D9143",
    x"3F2D95E1",
    x"3F2D9A7F",
    x"3F2D9F1D",
    x"3F2DA3BB",
    x"3F2DA859",
    x"3F2DACF7",
    x"3F2DB195",
    x"3F2DB632",
    x"3F2DBAD0",
    x"3F2DBF6D",
    x"3F2DC40A",
    x"3F2DC8A7",
    x"3F2DCD44",
    x"3F2DD1E1",
    x"3F2DD67E",
    x"3F2DDB1B",
    x"3F2DDFB8",
    x"3F2DE454",
    x"3F2DE8F0",
    x"3F2DED8D",
    x"3F2DF229",
    x"3F2DF6C5",
    x"3F2DFB61",
    x"3F2DFFFD",
    x"3F2E0499",
    x"3F2E0934",
    x"3F2E0DD0",
    x"3F2E126B",
    x"3F2E1707",
    x"3F2E1BA2",
    x"3F2E203D",
    x"3F2E24D8",
    x"3F2E2973",
    x"3F2E2E0E",
    x"3F2E32A9",
    x"3F2E3743",
    x"3F2E3BDE",
    x"3F2E4078",
    x"3F2E4513",
    x"3F2E49AD",
    x"3F2E4E47",
    x"3F2E52E1",
    x"3F2E577B",
    x"3F2E5C15",
    x"3F2E60AE",
    x"3F2E6548",
    x"3F2E69E1",
    x"3F2E6E7B",
    x"3F2E7314",
    x"3F2E77AD",
    x"3F2E7C46",
    x"3F2E80DF",
    x"3F2E8578",
    x"3F2E8A11",
    x"3F2E8EA9",
    x"3F2E9342",
    x"3F2E97DA",
    x"3F2E9C73",
    x"3F2EA10B",
    x"3F2EA5A3",
    x"3F2EAA3B",
    x"3F2EAED3",
    x"3F2EB36B",
    x"3F2EB802",
    x"3F2EBC9A",
    x"3F2EC131",
    x"3F2EC5C9",
    x"3F2ECA60",
    x"3F2ECEF7",
    x"3F2ED38E",
    x"3F2ED825",
    x"3F2EDCBC",
    x"3F2EE153",
    x"3F2EE5E9",
    x"3F2EEA80",
    x"3F2EEF16",
    x"3F2EF3AD",
    x"3F2EF843",
    x"3F2EFCD9",
    x"3F2F016F",
    x"3F2F0605",
    x"3F2F0A9B",
    x"3F2F0F30",
    x"3F2F13C6",
    x"3F2F185B",
    x"3F2F1CF1",
    x"3F2F2186",
    x"3F2F261B",
    x"3F2F2AB0",
    x"3F2F2F45",
    x"3F2F33DA",
    x"3F2F386F",
    x"3F2F3D03",
    x"3F2F4198",
    x"3F2F462C",
    x"3F2F4AC1",
    x"3F2F4F55",
    x"3F2F53E9",
    x"3F2F587D",
    x"3F2F5D11",
    x"3F2F61A5",
    x"3F2F6638",
    x"3F2F6ACC",
    x"3F2F6F5F",
    x"3F2F73F3",
    x"3F2F7886",
    x"3F2F7D19",
    x"3F2F81AC",
    x"3F2F863F",
    x"3F2F8AD2",
    x"3F2F8F65",
    x"3F2F93F7",
    x"3F2F988A",
    x"3F2F9D1C",
    x"3F2FA1AF",
    x"3F2FA641",
    x"3F2FAAD3",
    x"3F2FAF65",
    x"3F2FB3F7",
    x"3F2FB888",
    x"3F2FBD1A",
    x"3F2FC1AC",
    x"3F2FC63D",
    x"3F2FCACF",
    x"3F2FCF60",
    x"3F2FD3F1",
    x"3F2FD882",
    x"3F2FDD13",
    x"3F2FE1A4",
    x"3F2FE634",
    x"3F2FEAC5",
    x"3F2FEF56",
    x"3F2FF3E6",
    x"3F2FF876",
    x"3F2FFD06",
    x"3F300196",
    x"3F300626",
    x"3F300AB6",
    x"3F300F46",
    x"3F3013D6",
    x"3F301865",
    x"3F301CF5",
    x"3F302184",
    x"3F302613",
    x"3F302AA2",
    x"3F302F31",
    x"3F3033C0",
    x"3F30384F",
    x"3F303CDE",
    x"3F30416C",
    x"3F3045FB",
    x"3F304A89",
    x"3F304F18",
    x"3F3053A6",
    x"3F305834",
    x"3F305CC2",
    x"3F306150",
    x"3F3065DD",
    x"3F306A6B",
    x"3F306EF9",
    x"3F307386",
    x"3F307813",
    x"3F307CA1",
    x"3F30812E",
    x"3F3085BB",
    x"3F308A48",
    x"3F308ED4",
    x"3F309361",
    x"3F3097EE",
    x"3F309C7A",
    x"3F30A106",
    x"3F30A593",
    x"3F30AA1F",
    x"3F30AEAB",
    x"3F30B337",
    x"3F30B7C3",
    x"3F30BC4E",
    x"3F30C0DA",
    x"3F30C566",
    x"3F30C9F1",
    x"3F30CE7C",
    x"3F30D307",
    x"3F30D792",
    x"3F30DC1D",
    x"3F30E0A8",
    x"3F30E533",
    x"3F30E9BE",
    x"3F30EE48",
    x"3F30F2D3",
    x"3F30F75D",
    x"3F30FBE7",
    x"3F310071",
    x"3F3104FB",
    x"3F310985",
    x"3F310E0F",
    x"3F311299",
    x"3F311722",
    x"3F311BAC",
    x"3F312035",
    x"3F3124BF",
    x"3F312948",
    x"3F312DD1",
    x"3F31325A",
    x"3F3136E3",
    x"3F313B6B",
    x"3F313FF4",
    x"3F31447D",
    x"3F314905",
    x"3F314D8D",
    x"3F315215",
    x"3F31569E",
    x"3F315B26",
    x"3F315FAD",
    x"3F316435",
    x"3F3168BD",
    x"3F316D44",
    x"3F3171CC",
    x"3F317653",
    x"3F317ADB",
    x"3F317F62",
    x"3F3183E9",
    x"3F318870",
    x"3F318CF6",
    x"3F31917D",
    x"3F319604",
    x"3F319A8A",
    x"3F319F11",
    x"3F31A397",
    x"3F31A81D",
    x"3F31ACA3",
    x"3F31B129",
    x"3F31B5AF",
    x"3F31BA35",
    x"3F31BEBA",
    x"3F31C340",
    x"3F31C7C5",
    x"3F31CC4B",
    x"3F31D0D0",
    x"3F31D555",
    x"3F31D9DA",
    x"3F31DE5F",
    x"3F31E2E4",
    x"3F31E768",
    x"3F31EBED",
    x"3F31F071",
    x"3F31F4F6",
    x"3F31F97A",
    x"3F31FDFE",
    x"3F320282",
    x"3F320706",
    x"3F320B8A",
    x"3F32100E",
    x"3F321491",
    x"3F321915",
    x"3F321D98",
    x"3F32221B",
    x"3F32269E",
    x"3F322B22",
    x"3F322FA5",
    x"3F323427",
    x"3F3238AA",
    x"3F323D2D",
    x"3F3241AF",
    x"3F324632",
    x"3F324AB4",
    x"3F324F36",
    x"3F3253B8",
    x"3F32583A",
    x"3F325CBC",
    x"3F32613E",
    x"3F3265C0",
    x"3F326A41",
    x"3F326EC3",
    x"3F327344",
    x"3F3277C5",
    x"3F327C46",
    x"3F3280C7",
    x"3F328548",
    x"3F3289C9",
    x"3F328E4A",
    x"3F3292CA",
    x"3F32974B",
    x"3F329BCB",
    x"3F32A04C",
    x"3F32A4CC",
    x"3F32A94C",
    x"3F32ADCC",
    x"3F32B24C",
    x"3F32B6CB",
    x"3F32BB4B",
    x"3F32BFCA",
    x"3F32C44A",
    x"3F32C8C9",
    x"3F32CD48",
    x"3F32D1C7",
    x"3F32D646",
    x"3F32DAC5",
    x"3F32DF44",
    x"3F32E3C3",
    x"3F32E841",
    x"3F32ECC0",
    x"3F32F13E",
    x"3F32F5BC",
    x"3F32FA3A",
    x"3F32FEB8",
    x"3F330336",
    x"3F3307B4",
    x"3F330C32",
    x"3F3310AF",
    x"3F33152D",
    x"3F3319AA",
    x"3F331E27",
    x"3F3322A5",
    x"3F332722",
    x"3F332B9F",
    x"3F33301B",
    x"3F333498",
    x"3F333915",
    x"3F333D91",
    x"3F33420E",
    x"3F33468A",
    x"3F334B06",
    x"3F334F82",
    x"3F3353FE",
    x"3F33587A",
    x"3F335CF6",
    x"3F336171",
    x"3F3365ED",
    x"3F336A68",
    x"3F336EE4",
    x"3F33735F",
    x"3F3377DA",
    x"3F337C55",
    x"3F3380D0",
    x"3F33854B",
    x"3F3389C5",
    x"3F338E40",
    x"3F3392BA",
    x"3F339735",
    x"3F339BAF",
    x"3F33A029",
    x"3F33A4A3",
    x"3F33A91D",
    x"3F33AD97",
    x"3F33B210",
    x"3F33B68A",
    x"3F33BB03",
    x"3F33BF7D",
    x"3F33C3F6",
    x"3F33C86F",
    x"3F33CCE8",
    x"3F33D161",
    x"3F33D5DA",
    x"3F33DA53",
    x"3F33DECB",
    x"3F33E344",
    x"3F33E7BC",
    x"3F33EC34",
    x"3F33F0AD",
    x"3F33F525",
    x"3F33F99D",
    x"3F33FE14",
    x"3F34028C",
    x"3F340704",
    x"3F340B7B",
    x"3F340FF3",
    x"3F34146A",
    x"3F3418E1",
    x"3F341D58",
    x"3F3421CF",
    x"3F342646",
    x"3F342ABD",
    x"3F342F34",
    x"3F3433AA",
    x"3F343821",
    x"3F343C97",
    x"3F34410D",
    x"3F344583",
    x"3F3449F9",
    x"3F344E6F",
    x"3F3452E5",
    x"3F34575B",
    x"3F345BD0",
    x"3F346046",
    x"3F3464BB",
    x"3F346930",
    x"3F346DA5",
    x"3F34721A",
    x"3F34768F",
    x"3F347B04",
    x"3F347F79",
    x"3F3483ED",
    x"3F348862",
    x"3F348CD6",
    x"3F34914B",
    x"3F3495BF",
    x"3F349A33",
    x"3F349EA7",
    x"3F34A31B",
    x"3F34A78E",
    x"3F34AC02",
    x"3F34B075",
    x"3F34B4E9",
    x"3F34B95C",
    x"3F34BDCF",
    x"3F34C242",
    x"3F34C6B5",
    x"3F34CB28",
    x"3F34CF9B",
    x"3F34D40D",
    x"3F34D880",
    x"3F34DCF2",
    x"3F34E165",
    x"3F34E5D7",
    x"3F34EA49",
    x"3F34EEBB",
    x"3F34F32D",
    x"3F34F79F",
    x"3F34FC10",
    x"3F350082",
    x"3F3504F3",
    x"3F350965",
    x"3F350DD6",
    x"3F351247",
    x"3F3516B8",
    x"3F351B29",
    x"3F351F9A",
    x"3F35240A",
    x"3F35287B",
    x"3F352CEB",
    x"3F35315C",
    x"3F3535CC",
    x"3F353A3C",
    x"3F353EAC",
    x"3F35431C",
    x"3F35478C",
    x"3F354BFB",
    x"3F35506B",
    x"3F3554DA",
    x"3F35594A",
    x"3F355DB9",
    x"3F356228",
    x"3F356697",
    x"3F356B06",
    x"3F356F75",
    x"3F3573E4",
    x"3F357852",
    x"3F357CC1",
    x"3F35812F",
    x"3F35859D",
    x"3F358A0B",
    x"3F358E79",
    x"3F3592E7",
    x"3F359755",
    x"3F359BC3",
    x"3F35A031",
    x"3F35A49E",
    x"3F35A90B",
    x"3F35AD79",
    x"3F35B1E6",
    x"3F35B653",
    x"3F35BAC0",
    x"3F35BF2D",
    x"3F35C39A",
    x"3F35C806",
    x"3F35CC73",
    x"3F35D0DF",
    x"3F35D54B",
    x"3F35D9B8",
    x"3F35DE24",
    x"3F35E290",
    x"3F35E6FB",
    x"3F35EB67",
    x"3F35EFD3",
    x"3F35F43E",
    x"3F35F8AA",
    x"3F35FD15",
    x"3F360180",
    x"3F3605EB",
    x"3F360A56",
    x"3F360EC1",
    x"3F36132C",
    x"3F361797",
    x"3F361C01",
    x"3F36206C",
    x"3F3624D6",
    x"3F362940",
    x"3F362DAA",
    x"3F363214",
    x"3F36367E",
    x"3F363AE8",
    x"3F363F52",
    x"3F3643BB",
    x"3F364825",
    x"3F364C8E",
    x"3F3650F7",
    x"3F365560",
    x"3F3659C9",
    x"3F365E32",
    x"3F36629B",
    x"3F366704",
    x"3F366B6C",
    x"3F366FD5",
    x"3F36743D",
    x"3F3678A5",
    x"3F367D0D",
    x"3F368175",
    x"3F3685DD",
    x"3F368A45",
    x"3F368EAD",
    x"3F369314",
    x"3F36977C",
    x"3F369BE3",
    x"3F36A04A",
    x"3F36A4B2",
    x"3F36A919",
    x"3F36AD7F",
    x"3F36B1E6",
    x"3F36B64D",
    x"3F36BAB4",
    x"3F36BF1A",
    x"3F36C380",
    x"3F36C7E7",
    x"3F36CC4D",
    x"3F36D0B3",
    x"3F36D519",
    x"3F36D97F",
    x"3F36DDE4",
    x"3F36E24A",
    x"3F36E6AF",
    x"3F36EB15",
    x"3F36EF7A",
    x"3F36F3DF",
    x"3F36F844",
    x"3F36FCA9",
    x"3F37010E",
    x"3F370573",
    x"3F3709D7",
    x"3F370E3C",
    x"3F3712A0",
    x"3F371704",
    x"3F371B69",
    x"3F371FCD",
    x"3F372431",
    x"3F372894",
    x"3F372CF8",
    x"3F37315C",
    x"3F3735BF",
    x"3F373A23",
    x"3F373E86",
    x"3F3742E9",
    x"3F37474C",
    x"3F374BAF",
    x"3F375012",
    x"3F375475",
    x"3F3758D7",
    x"3F375D3A",
    x"3F37619C",
    x"3F3765FE",
    x"3F376A61",
    x"3F376EC3",
    x"3F377325",
    x"3F377787",
    x"3F377BE8",
    x"3F37804A",
    x"3F3784AB",
    x"3F37890D",
    x"3F378D6E",
    x"3F3791CF",
    x"3F379630",
    x"3F379A91",
    x"3F379EF2",
    x"3F37A353",
    x"3F37A7B4",
    x"3F37AC14",
    x"3F37B074",
    x"3F37B4D5",
    x"3F37B935",
    x"3F37BD95",
    x"3F37C1F5",
    x"3F37C655",
    x"3F37CAB5",
    x"3F37CF14",
    x"3F37D374",
    x"3F37D7D3",
    x"3F37DC32",
    x"3F37E092",
    x"3F37E4F1",
    x"3F37E950",
    x"3F37EDAF",
    x"3F37F20D",
    x"3F37F66C",
    x"3F37FACA",
    x"3F37FF29",
    x"3F380387",
    x"3F3807E5",
    x"3F380C43",
    x"3F3810A1",
    x"3F3814FF",
    x"3F38195D",
    x"3F381DBB",
    x"3F382218",
    x"3F382676",
    x"3F382AD3",
    x"3F382F30",
    x"3F38338D",
    x"3F3837EA",
    x"3F383C47",
    x"3F3840A4",
    x"3F384500",
    x"3F38495D",
    x"3F384DB9",
    x"3F385216",
    x"3F385672",
    x"3F385ACE",
    x"3F385F2A",
    x"3F386386",
    x"3F3867E1",
    x"3F386C3D",
    x"3F387099",
    x"3F3874F4",
    x"3F38794F",
    x"3F387DAB",
    x"3F388206",
    x"3F388661",
    x"3F388ABB",
    x"3F388F16",
    x"3F389371",
    x"3F3897CB",
    x"3F389C26",
    x"3F38A080",
    x"3F38A4DA",
    x"3F38A934",
    x"3F38AD8E",
    x"3F38B1E8",
    x"3F38B642",
    x"3F38BA9C",
    x"3F38BEF5",
    x"3F38C34F",
    x"3F38C7A8",
    x"3F38CC01",
    x"3F38D05A",
    x"3F38D4B3",
    x"3F38D90C",
    x"3F38DD65",
    x"3F38E1BD",
    x"3F38E616",
    x"3F38EA6E",
    x"3F38EEC7",
    x"3F38F31F",
    x"3F38F777",
    x"3F38FBCF",
    x"3F390027",
    x"3F39047E",
    x"3F3908D6",
    x"3F390D2E",
    x"3F391185",
    x"3F3915DC",
    x"3F391A33",
    x"3F391E8B",
    x"3F3922E1",
    x"3F392738",
    x"3F392B8F",
    x"3F392FE6",
    x"3F39343C",
    x"3F393893",
    x"3F393CE9",
    x"3F39413F",
    x"3F394595",
    x"3F3949EB",
    x"3F394E41",
    x"3F395297",
    x"3F3956EC",
    x"3F395B42",
    x"3F395F97",
    x"3F3963ED",
    x"3F396842",
    x"3F396C97",
    x"3F3970EC",
    x"3F397541",
    x"3F397995",
    x"3F397DEA",
    x"3F39823E",
    x"3F398693",
    x"3F398AE7",
    x"3F398F3B",
    x"3F39938F",
    x"3F3997E3",
    x"3F399C37",
    x"3F39A08B",
    x"3F39A4DF",
    x"3F39A932",
    x"3F39AD85",
    x"3F39B1D9",
    x"3F39B62C",
    x"3F39BA7F",
    x"3F39BED2",
    x"3F39C325",
    x"3F39C777",
    x"3F39CBCA",
    x"3F39D01D",
    x"3F39D46F",
    x"3F39D8C1",
    x"3F39DD13",
    x"3F39E165",
    x"3F39E5B7",
    x"3F39EA09",
    x"3F39EE5B",
    x"3F39F2AC",
    x"3F39F6FE",
    x"3F39FB4F",
    x"3F39FFA1",
    x"3F3A03F2",
    x"3F3A0843",
    x"3F3A0C94",
    x"3F3A10E4",
    x"3F3A1535",
    x"3F3A1986",
    x"3F3A1DD6",
    x"3F3A2227",
    x"3F3A2677",
    x"3F3A2AC7",
    x"3F3A2F17",
    x"3F3A3367",
    x"3F3A37B7",
    x"3F3A3C06",
    x"3F3A4056",
    x"3F3A44A6",
    x"3F3A48F5",
    x"3F3A4D44",
    x"3F3A5193",
    x"3F3A55E2",
    x"3F3A5A31",
    x"3F3A5E80",
    x"3F3A62CF",
    x"3F3A671D",
    x"3F3A6B6C",
    x"3F3A6FBA",
    x"3F3A7408",
    x"3F3A7856",
    x"3F3A7CA4",
    x"3F3A80F2",
    x"3F3A8540",
    x"3F3A898E",
    x"3F3A8DDB",
    x"3F3A9229",
    x"3F3A9676",
    x"3F3A9AC3",
    x"3F3A9F10",
    x"3F3AA35D",
    x"3F3AA7AA",
    x"3F3AABF7",
    x"3F3AB044",
    x"3F3AB490",
    x"3F3AB8DD",
    x"3F3ABD29",
    x"3F3AC175",
    x"3F3AC5C1",
    x"3F3ACA0D",
    x"3F3ACE59",
    x"3F3AD2A5",
    x"3F3AD6F1",
    x"3F3ADB3C",
    x"3F3ADF88",
    x"3F3AE3D3",
    x"3F3AE81E",
    x"3F3AEC69",
    x"3F3AF0B4",
    x"3F3AF4FF",
    x"3F3AF94A",
    x"3F3AFD94",
    x"3F3B01DF",
    x"3F3B0629",
    x"3F3B0A74",
    x"3F3B0EBE",
    x"3F3B1308",
    x"3F3B1752",
    x"3F3B1B9C",
    x"3F3B1FE5",
    x"3F3B242F",
    x"3F3B2879",
    x"3F3B2CC2",
    x"3F3B310B",
    x"3F3B3554",
    x"3F3B399E",
    x"3F3B3DE6",
    x"3F3B422F",
    x"3F3B4678",
    x"3F3B4AC1",
    x"3F3B4F09",
    x"3F3B5351",
    x"3F3B579A",
    x"3F3B5BE2",
    x"3F3B602A",
    x"3F3B6472",
    x"3F3B68BA",
    x"3F3B6D01",
    x"3F3B7149",
    x"3F3B7590",
    x"3F3B79D8",
    x"3F3B7E1F",
    x"3F3B8266",
    x"3F3B86AD",
    x"3F3B8AF4",
    x"3F3B8F3B",
    x"3F3B9382",
    x"3F3B97C8",
    x"3F3B9C0F",
    x"3F3BA055",
    x"3F3BA49B",
    x"3F3BA8E1",
    x"3F3BAD27",
    x"3F3BB16D",
    x"3F3BB5B3",
    x"3F3BB9F9",
    x"3F3BBE3E",
    x"3F3BC284",
    x"3F3BC6C9",
    x"3F3BCB0E",
    x"3F3BCF53",
    x"3F3BD398",
    x"3F3BD7DD",
    x"3F3BDC22",
    x"3F3BE067",
    x"3F3BE4AB",
    x"3F3BE8F0",
    x"3F3BED34",
    x"3F3BF178",
    x"3F3BF5BC",
    x"3F3BFA00",
    x"3F3BFE44",
    x"3F3C0288",
    x"3F3C06CB",
    x"3F3C0B0F",
    x"3F3C0F52",
    x"3F3C1396",
    x"3F3C17D9",
    x"3F3C1C1C",
    x"3F3C205F",
    x"3F3C24A2",
    x"3F3C28E4",
    x"3F3C2D27",
    x"3F3C316A",
    x"3F3C35AC",
    x"3F3C39EE",
    x"3F3C3E30",
    x"3F3C4272",
    x"3F3C46B4",
    x"3F3C4AF6",
    x"3F3C4F38",
    x"3F3C5379",
    x"3F3C57BB",
    x"3F3C5BFC",
    x"3F3C603E",
    x"3F3C647F",
    x"3F3C68C0",
    x"3F3C6D01",
    x"3F3C7141",
    x"3F3C7582",
    x"3F3C79C3",
    x"3F3C7E03",
    x"3F3C8244",
    x"3F3C8684",
    x"3F3C8AC4",
    x"3F3C8F04",
    x"3F3C9344",
    x"3F3C9784",
    x"3F3C9BC3",
    x"3F3CA003",
    x"3F3CA442",
    x"3F3CA881",
    x"3F3CACC1",
    x"3F3CB100",
    x"3F3CB53F",
    x"3F3CB97E",
    x"3F3CBDBC",
    x"3F3CC1FB",
    x"3F3CC63A",
    x"3F3CCA78",
    x"3F3CCEB6",
    x"3F3CD2F4",
    x"3F3CD733",
    x"3F3CDB70",
    x"3F3CDFAE",
    x"3F3CE3EC",
    x"3F3CE82A",
    x"3F3CEC67",
    x"3F3CF0A5",
    x"3F3CF4E2",
    x"3F3CF91F",
    x"3F3CFD5C",
    x"3F3D0199",
    x"3F3D05D6",
    x"3F3D0A12",
    x"3F3D0E4F",
    x"3F3D128C",
    x"3F3D16C8",
    x"3F3D1B04",
    x"3F3D1F40",
    x"3F3D237C",
    x"3F3D27B8",
    x"3F3D2BF4",
    x"3F3D3030",
    x"3F3D346B",
    x"3F3D38A7",
    x"3F3D3CE2",
    x"3F3D411D",
    x"3F3D4558",
    x"3F3D4993",
    x"3F3D4DCE",
    x"3F3D5209",
    x"3F3D5644",
    x"3F3D5A7E",
    x"3F3D5EB9",
    x"3F3D62F3",
    x"3F3D672D",
    x"3F3D6B67",
    x"3F3D6FA1",
    x"3F3D73DB",
    x"3F3D7815",
    x"3F3D7C4E",
    x"3F3D8088",
    x"3F3D84C1",
    x"3F3D88FB",
    x"3F3D8D34",
    x"3F3D916D",
    x"3F3D95A6",
    x"3F3D99DF",
    x"3F3D9E17",
    x"3F3DA250",
    x"3F3DA688",
    x"3F3DAAC1",
    x"3F3DAEF9",
    x"3F3DB331",
    x"3F3DB769",
    x"3F3DBBA1",
    x"3F3DBFD9",
    x"3F3DC411",
    x"3F3DC848",
    x"3F3DCC80",
    x"3F3DD0B7",
    x"3F3DD4EE",
    x"3F3DD925",
    x"3F3DDD5C",
    x"3F3DE193",
    x"3F3DE5CA",
    x"3F3DEA01",
    x"3F3DEE37",
    x"3F3DF26E",
    x"3F3DF6A4",
    x"3F3DFADA",
    x"3F3DFF10",
    x"3F3E0346",
    x"3F3E077C",
    x"3F3E0BB2",
    x"3F3E0FE7",
    x"3F3E141D",
    x"3F3E1852",
    x"3F3E1C88",
    x"3F3E20BD",
    x"3F3E24F2",
    x"3F3E2927",
    x"3F3E2D5C",
    x"3F3E3190",
    x"3F3E35C5",
    x"3F3E39F9",
    x"3F3E3E2E",
    x"3F3E4262",
    x"3F3E4696",
    x"3F3E4ACA",
    x"3F3E4EFE",
    x"3F3E5332",
    x"3F3E5766",
    x"3F3E5B99",
    x"3F3E5FCD",
    x"3F3E6400",
    x"3F3E6833",
    x"3F3E6C66",
    x"3F3E7099",
    x"3F3E74CC",
    x"3F3E78FF",
    x"3F3E7D31",
    x"3F3E8164",
    x"3F3E8596",
    x"3F3E89C9",
    x"3F3E8DFB",
    x"3F3E922D",
    x"3F3E965F",
    x"3F3E9A91",
    x"3F3E9EC3",
    x"3F3EA2F4",
    x"3F3EA726",
    x"3F3EAB57",
    x"3F3EAF88",
    x"3F3EB3B9",
    x"3F3EB7EA",
    x"3F3EBC1B",
    x"3F3EC04C",
    x"3F3EC47D",
    x"3F3EC8AD",
    x"3F3ECCDE",
    x"3F3ED10E",
    x"3F3ED53F",
    x"3F3ED96F",
    x"3F3EDD9F",
    x"3F3EE1CF",
    x"3F3EE5FE",
    x"3F3EEA2E",
    x"3F3EEE5E",
    x"3F3EF28D",
    x"3F3EF6BC",
    x"3F3EFAEB",
    x"3F3EFF1B",
    x"3F3F034A",
    x"3F3F0778",
    x"3F3F0BA7",
    x"3F3F0FD6",
    x"3F3F1404",
    x"3F3F1833",
    x"3F3F1C61",
    x"3F3F208F",
    x"3F3F24BD",
    x"3F3F28EB",
    x"3F3F2D19",
    x"3F3F3147",
    x"3F3F3574",
    x"3F3F39A2",
    x"3F3F3DCF",
    x"3F3F41FC",
    x"3F3F4629",
    x"3F3F4A56",
    x"3F3F4E83",
    x"3F3F52B0",
    x"3F3F56DD",
    x"3F3F5B09",
    x"3F3F5F36",
    x"3F3F6362",
    x"3F3F678E",
    x"3F3F6BBA",
    x"3F3F6FE6",
    x"3F3F7412",
    x"3F3F783E",
    x"3F3F7C6A",
    x"3F3F8095",
    x"3F3F84C0",
    x"3F3F88EC",
    x"3F3F8D17",
    x"3F3F9142",
    x"3F3F956D",
    x"3F3F9998",
    x"3F3F9DC2",
    x"3F3FA1ED",
    x"3F3FA617",
    x"3F3FAA42",
    x"3F3FAE6C",
    x"3F3FB296",
    x"3F3FB6C0",
    x"3F3FBAEA",
    x"3F3FBF14",
    x"3F3FC33E",
    x"3F3FC767",
    x"3F3FCB91",
    x"3F3FCFBA",
    x"3F3FD3E3",
    x"3F3FD80C",
    x"3F3FDC35",
    x"3F3FE05E",
    x"3F3FE487",
    x"3F3FE8AF",
    x"3F3FECD8",
    x"3F3FF100",
    x"3F3FF529",
    x"3F3FF951",
    x"3F3FFD79",
    x"3F4001A1",
    x"3F4005C8",
    x"3F4009F0",
    x"3F400E18",
    x"3F40123F",
    x"3F401667",
    x"3F401A8E",
    x"3F401EB5",
    x"3F4022DC",
    x"3F402703",
    x"3F402B2A",
    x"3F402F50",
    x"3F403377",
    x"3F40379D",
    x"3F403BC4",
    x"3F403FEA",
    x"3F404410",
    x"3F404836",
    x"3F404C5C",
    x"3F405081",
    x"3F4054A7",
    x"3F4058CD",
    x"3F405CF2",
    x"3F406117",
    x"3F40653C",
    x"3F406961",
    x"3F406D86",
    x"3F4071AB",
    x"3F4075D0",
    x"3F4079F4",
    x"3F407E19",
    x"3F40823D",
    x"3F408661",
    x"3F408A85",
    x"3F408EA9",
    x"3F4092CD",
    x"3F4096F1",
    x"3F409B15",
    x"3F409F38",
    x"3F40A35C",
    x"3F40A77F",
    x"3F40ABA2",
    x"3F40AFC5",
    x"3F40B3E8",
    x"3F40B80B",
    x"3F40BC2E",
    x"3F40C050",
    x"3F40C473",
    x"3F40C895",
    x"3F40CCB7",
    x"3F40D0DA",
    x"3F40D4FC",
    x"3F40D91E",
    x"3F40DD3F",
    x"3F40E161",
    x"3F40E583",
    x"3F40E9A4",
    x"3F40EDC5",
    x"3F40F1E7",
    x"3F40F608",
    x"3F40FA29",
    x"3F40FE49",
    x"3F41026A",
    x"3F41068B",
    x"3F410AAB",
    x"3F410ECC",
    x"3F4112EC",
    x"3F41170C",
    x"3F411B2C",
    x"3F411F4C",
    x"3F41236C",
    x"3F41278C",
    x"3F412BAB",
    x"3F412FCB",
    x"3F4133EA",
    x"3F413809",
    x"3F413C28",
    x"3F414047",
    x"3F414466",
    x"3F414885",
    x"3F414CA4",
    x"3F4150C2",
    x"3F4154E1",
    x"3F4158FF",
    x"3F415D1D",
    x"3F41613B",
    x"3F416559",
    x"3F416977",
    x"3F416D95",
    x"3F4171B2",
    x"3F4175D0",
    x"3F4179ED",
    x"3F417E0A",
    x"3F418228",
    x"3F418645",
    x"3F418A61",
    x"3F418E7E",
    x"3F41929B",
    x"3F4196B7",
    x"3F419AD4",
    x"3F419EF0",
    x"3F41A30C",
    x"3F41A728",
    x"3F41AB44",
    x"3F41AF60",
    x"3F41B37C",
    x"3F41B798",
    x"3F41BBB3",
    x"3F41BFCF",
    x"3F41C3EA",
    x"3F41C805",
    x"3F41CC20",
    x"3F41D03B",
    x"3F41D456",
    x"3F41D870",
    x"3F41DC8B",
    x"3F41E0A5",
    x"3F41E4C0",
    x"3F41E8DA",
    x"3F41ECF4",
    x"3F41F10E",
    x"3F41F528",
    x"3F41F942",
    x"3F41FD5B",
    x"3F420175",
    x"3F42058E",
    x"3F4209A7",
    x"3F420DC1",
    x"3F4211DA",
    x"3F4215F3",
    x"3F421A0B",
    x"3F421E24",
    x"3F42223D",
    x"3F422655",
    x"3F422A6E",
    x"3F422E86",
    x"3F42329E",
    x"3F4236B6",
    x"3F423ACE",
    x"3F423EE5",
    x"3F4242FD",
    x"3F424715",
    x"3F424B2C",
    x"3F424F43",
    x"3F42535B",
    x"3F425772",
    x"3F425B89",
    x"3F425F9F",
    x"3F4263B6",
    x"3F4267CD",
    x"3F426BE3",
    x"3F426FFA",
    x"3F427410",
    x"3F427826",
    x"3F427C3C",
    x"3F428052",
    x"3F428468",
    x"3F42887D",
    x"3F428C93",
    x"3F4290A8",
    x"3F4294BD",
    x"3F4298D3",
    x"3F429CE8",
    x"3F42A0FD",
    x"3F42A511",
    x"3F42A926",
    x"3F42AD3B",
    x"3F42B14F",
    x"3F42B564",
    x"3F42B978",
    x"3F42BD8C",
    x"3F42C1A0",
    x"3F42C5B4",
    x"3F42C9C8",
    x"3F42CDDB",
    x"3F42D1EF",
    x"3F42D602",
    x"3F42DA16",
    x"3F42DE29",
    x"3F42E23C",
    x"3F42E64F",
    x"3F42EA62",
    x"3F42EE74",
    x"3F42F287",
    x"3F42F69A",
    x"3F42FAAC",
    x"3F42FEBE",
    x"3F4302D0",
    x"3F4306E2",
    x"3F430AF4",
    x"3F430F06",
    x"3F431318",
    x"3F431729",
    x"3F431B3B",
    x"3F431F4C",
    x"3F43235D",
    x"3F43276E",
    x"3F432B7F",
    x"3F432F90",
    x"3F4333A1",
    x"3F4337B1",
    x"3F433BC2",
    x"3F433FD2",
    x"3F4343E2",
    x"3F4347F3",
    x"3F434C03",
    x"3F435012",
    x"3F435422",
    x"3F435832",
    x"3F435C41",
    x"3F436051",
    x"3F436460",
    x"3F43686F",
    x"3F436C7F",
    x"3F43708D",
    x"3F43749C",
    x"3F4378AB",
    x"3F437CBA",
    x"3F4380C8",
    x"3F4384D6",
    x"3F4388E5",
    x"3F438CF3",
    x"3F439101",
    x"3F43950F",
    x"3F43991D",
    x"3F439D2A",
    x"3F43A138",
    x"3F43A545",
    x"3F43A953",
    x"3F43AD60",
    x"3F43B16D",
    x"3F43B57A",
    x"3F43B987",
    x"3F43BD93",
    x"3F43C1A0",
    x"3F43C5AC",
    x"3F43C9B9",
    x"3F43CDC5",
    x"3F43D1D1",
    x"3F43D5DD",
    x"3F43D9E9",
    x"3F43DDF5",
    x"3F43E200",
    x"3F43E60C",
    x"3F43EA17",
    x"3F43EE23",
    x"3F43F22E",
    x"3F43F639",
    x"3F43FA44",
    x"3F43FE4F",
    x"3F44025A",
    x"3F440664",
    x"3F440A6F",
    x"3F440E79",
    x"3F441283",
    x"3F44168D",
    x"3F441A97",
    x"3F441EA1",
    x"3F4422AB",
    x"3F4426B5",
    x"3F442ABE",
    x"3F442EC8",
    x"3F4432D1",
    x"3F4436DA",
    x"3F443AE3",
    x"3F443EEC",
    x"3F4442F5",
    x"3F4446FE",
    x"3F444B06",
    x"3F444F0F",
    x"3F445317",
    x"3F44571F",
    x"3F445B27",
    x"3F445F2F",
    x"3F446337",
    x"3F44673F",
    x"3F446B47",
    x"3F446F4E",
    x"3F447356",
    x"3F44775D",
    x"3F447B64",
    x"3F447F6B",
    x"3F448372",
    x"3F448779",
    x"3F448B80",
    x"3F448F86",
    x"3F44938D",
    x"3F449793",
    x"3F449B99",
    x"3F449F9F",
    x"3F44A3A5",
    x"3F44A7AB",
    x"3F44ABB1",
    x"3F44AFB6",
    x"3F44B3BC",
    x"3F44B7C1",
    x"3F44BBC7",
    x"3F44BFCC",
    x"3F44C3D1",
    x"3F44C7D6",
    x"3F44CBDB",
    x"3F44CFDF",
    x"3F44D3E4",
    x"3F44D7E8",
    x"3F44DBED",
    x"3F44DFF1",
    x"3F44E3F5",
    x"3F44E7F9",
    x"3F44EBFD",
    x"3F44F000",
    x"3F44F404",
    x"3F44F807",
    x"3F44FC0B",
    x"3F45000E",
    x"3F450411",
    x"3F450814",
    x"3F450C17",
    x"3F45101A",
    x"3F45141D",
    x"3F45181F",
    x"3F451C22",
    x"3F452024",
    x"3F452426",
    x"3F452828",
    x"3F452C2A",
    x"3F45302C",
    x"3F45342E",
    x"3F45382F",
    x"3F453C31",
    x"3F454032",
    x"3F454433",
    x"3F454834",
    x"3F454C35",
    x"3F455036",
    x"3F455437",
    x"3F455838",
    x"3F455C38",
    x"3F456039",
    x"3F456439",
    x"3F456839",
    x"3F456C39",
    x"3F457039",
    x"3F457439",
    x"3F457839",
    x"3F457C38",
    x"3F458038",
    x"3F458437",
    x"3F458836",
    x"3F458C35",
    x"3F459034",
    x"3F459433",
    x"3F459832",
    x"3F459C31",
    x"3F45A02F",
    x"3F45A42D",
    x"3F45A82C",
    x"3F45AC2A",
    x"3F45B028",
    x"3F45B426",
    x"3F45B824",
    x"3F45BC21",
    x"3F45C01F",
    x"3F45C41C",
    x"3F45C819",
    x"3F45CC17",
    x"3F45D014",
    x"3F45D411",
    x"3F45D80E",
    x"3F45DC0A",
    x"3F45E007",
    x"3F45E403",
    x"3F45E800",
    x"3F45EBFC",
    x"3F45EFF8",
    x"3F45F3F4",
    x"3F45F7F0",
    x"3F45FBEC",
    x"3F45FFE7",
    x"3F4603E3",
    x"3F4607DE",
    x"3F460BDA",
    x"3F460FD5",
    x"3F4613D0",
    x"3F4617CB",
    x"3F461BC6",
    x"3F461FC0",
    x"3F4623BB",
    x"3F4627B5",
    x"3F462BB0",
    x"3F462FAA",
    x"3F4633A4",
    x"3F46379E",
    x"3F463B98",
    x"3F463F91",
    x"3F46438B",
    x"3F464785",
    x"3F464B7E",
    x"3F464F77",
    x"3F465370",
    x"3F465769",
    x"3F465B62",
    x"3F465F5B",
    x"3F466354",
    x"3F46674C",
    x"3F466B45",
    x"3F466F3D",
    x"3F467335",
    x"3F46772D",
    x"3F467B25",
    x"3F467F1D",
    x"3F468315",
    x"3F46870C",
    x"3F468B04",
    x"3F468EFB",
    x"3F4692F2",
    x"3F4696E9",
    x"3F469AE0",
    x"3F469ED7",
    x"3F46A2CE",
    x"3F46A6C5",
    x"3F46AABB",
    x"3F46AEB1",
    x"3F46B2A8",
    x"3F46B69E",
    x"3F46BA94",
    x"3F46BE8A",
    x"3F46C280",
    x"3F46C675",
    x"3F46CA6B",
    x"3F46CE60",
    x"3F46D256",
    x"3F46D64B",
    x"3F46DA40",
    x"3F46DE35",
    x"3F46E22A",
    x"3F46E61E",
    x"3F46EA13",
    x"3F46EE07",
    x"3F46F1FC",
    x"3F46F5F0",
    x"3F46F9E4",
    x"3F46FDD8",
    x"3F4701CC",
    x"3F4705C0",
    x"3F4709B3",
    x"3F470DA7",
    x"3F47119A",
    x"3F47158D",
    x"3F471981",
    x"3F471D74",
    x"3F472167",
    x"3F472559",
    x"3F47294C",
    x"3F472D3F",
    x"3F473131",
    x"3F473523",
    x"3F473916",
    x"3F473D08",
    x"3F4740FA",
    x"3F4744EB",
    x"3F4748DD",
    x"3F474CCF",
    x"3F4750C0",
    x"3F4754B2",
    x"3F4758A3",
    x"3F475C94",
    x"3F476085",
    x"3F476476",
    x"3F476866",
    x"3F476C57",
    x"3F477048",
    x"3F477438",
    x"3F477828",
    x"3F477C18",
    x"3F478008",
    x"3F4783F8",
    x"3F4787E8",
    x"3F478BD8",
    x"3F478FC7",
    x"3F4793B7",
    x"3F4797A6",
    x"3F479B95",
    x"3F479F84",
    x"3F47A373",
    x"3F47A762",
    x"3F47AB51",
    x"3F47AF3F",
    x"3F47B32E",
    x"3F47B71C",
    x"3F47BB0A",
    x"3F47BEF9",
    x"3F47C2E7",
    x"3F47C6D4",
    x"3F47CAC2",
    x"3F47CEB0",
    x"3F47D29D",
    x"3F47D68B",
    x"3F47DA78",
    x"3F47DE65",
    x"3F47E252",
    x"3F47E63F",
    x"3F47EA2C",
    x"3F47EE18",
    x"3F47F205",
    x"3F47F5F1",
    x"3F47F9DE",
    x"3F47FDCA",
    x"3F4801B6",
    x"3F4805A2",
    x"3F48098E",
    x"3F480D79",
    x"3F481165",
    x"3F481550",
    x"3F48193C",
    x"3F481D27",
    x"3F482112",
    x"3F4824FD",
    x"3F4828E8",
    x"3F482CD3",
    x"3F4830BD",
    x"3F4834A8",
    x"3F483892",
    x"3F483C7C",
    x"3F484067",
    x"3F484451",
    x"3F48483A",
    x"3F484C24",
    x"3F48500E",
    x"3F4853F7",
    x"3F4857E1",
    x"3F485BCA",
    x"3F485FB3",
    x"3F48639C",
    x"3F486785",
    x"3F486B6E",
    x"3F486F57",
    x"3F48733F",
    x"3F487728",
    x"3F487B10",
    x"3F487EF8",
    x"3F4882E0",
    x"3F4886C8",
    x"3F488AB0",
    x"3F488E98",
    x"3F48927F",
    x"3F489667",
    x"3F489A4E",
    x"3F489E36",
    x"3F48A21D",
    x"3F48A604",
    x"3F48A9EA",
    x"3F48ADD1",
    x"3F48B1B8",
    x"3F48B59E",
    x"3F48B985",
    x"3F48BD6B",
    x"3F48C151",
    x"3F48C537",
    x"3F48C91D",
    x"3F48CD03",
    x"3F48D0E9",
    x"3F48D4CE",
    x"3F48D8B3",
    x"3F48DC99",
    x"3F48E07E",
    x"3F48E463",
    x"3F48E848",
    x"3F48EC2D",
    x"3F48F011",
    x"3F48F3F6",
    x"3F48F7DA",
    x"3F48FBBF",
    x"3F48FFA3",
    x"3F490387",
    x"3F49076B",
    x"3F490B4F",
    x"3F490F33",
    x"3F491316",
    x"3F4916FA",
    x"3F491ADD",
    x"3F491EC0",
    x"3F4922A3",
    x"3F492686",
    x"3F492A69",
    x"3F492E4C",
    x"3F49322F",
    x"3F493611",
    x"3F4939F4",
    x"3F493DD6",
    x"3F4941B8",
    x"3F49459A",
    x"3F49497C",
    x"3F494D5E",
    x"3F49513F",
    x"3F495521",
    x"3F495902",
    x"3F495CE4",
    x"3F4960C5",
    x"3F4964A6",
    x"3F496887",
    x"3F496C68",
    x"3F497048",
    x"3F497429",
    x"3F497809",
    x"3F497BEA",
    x"3F497FCA",
    x"3F4983AA",
    x"3F49878A",
    x"3F498B6A",
    x"3F498F4A",
    x"3F499329",
    x"3F499709",
    x"3F499AE8",
    x"3F499EC7",
    x"3F49A2A6",
    x"3F49A685",
    x"3F49AA64",
    x"3F49AE43",
    x"3F49B222",
    x"3F49B600",
    x"3F49B9DF",
    x"3F49BDBD",
    x"3F49C19B",
    x"3F49C579",
    x"3F49C957",
    x"3F49CD35",
    x"3F49D112",
    x"3F49D4F0",
    x"3F49D8CD",
    x"3F49DCAB",
    x"3F49E088",
    x"3F49E465",
    x"3F49E842",
    x"3F49EC1F",
    x"3F49EFFB",
    x"3F49F3D8",
    x"3F49F7B4",
    x"3F49FB91",
    x"3F49FF6D",
    x"3F4A0349",
    x"3F4A0725",
    x"3F4A0B01",
    x"3F4A0EDC",
    x"3F4A12B8",
    x"3F4A1693",
    x"3F4A1A6F",
    x"3F4A1E4A",
    x"3F4A2225",
    x"3F4A2600",
    x"3F4A29DB",
    x"3F4A2DB6",
    x"3F4A3190",
    x"3F4A356B",
    x"3F4A3945",
    x"3F4A3D1F",
    x"3F4A40F9",
    x"3F4A44D3",
    x"3F4A48AD",
    x"3F4A4C87",
    x"3F4A5061",
    x"3F4A543A",
    x"3F4A5814",
    x"3F4A5BED",
    x"3F4A5FC6",
    x"3F4A639F",
    x"3F4A6778",
    x"3F4A6B51",
    x"3F4A6F29",
    x"3F4A7302",
    x"3F4A76DA",
    x"3F4A7AB3",
    x"3F4A7E8B",
    x"3F4A8263",
    x"3F4A863B",
    x"3F4A8A13",
    x"3F4A8DEA",
    x"3F4A91C2",
    x"3F4A9599",
    x"3F4A9971",
    x"3F4A9D48",
    x"3F4AA11F",
    x"3F4AA4F6",
    x"3F4AA8CD",
    x"3F4AACA4",
    x"3F4AB07A",
    x"3F4AB451",
    x"3F4AB827",
    x"3F4ABBFD",
    x"3F4ABFD3",
    x"3F4AC3A9",
    x"3F4AC77F",
    x"3F4ACB55",
    x"3F4ACF2A",
    x"3F4AD300",
    x"3F4AD6D5",
    x"3F4ADAAB",
    x"3F4ADE80",
    x"3F4AE255",
    x"3F4AE62A",
    x"3F4AE9FE",
    x"3F4AEDD3",
    x"3F4AF1A8",
    x"3F4AF57C",
    x"3F4AF950",
    x"3F4AFD24",
    x"3F4B00F8",
    x"3F4B04CC",
    x"3F4B08A0",
    x"3F4B0C74",
    x"3F4B1047",
    x"3F4B141B",
    x"3F4B17EE",
    x"3F4B1BC1",
    x"3F4B1F94",
    x"3F4B2367",
    x"3F4B273A",
    x"3F4B2B0D",
    x"3F4B2EDF",
    x"3F4B32B2",
    x"3F4B3684",
    x"3F4B3A56",
    x"3F4B3E28",
    x"3F4B41FA",
    x"3F4B45CC",
    x"3F4B499E",
    x"3F4B4D6F",
    x"3F4B5141",
    x"3F4B5512",
    x"3F4B58E3",
    x"3F4B5CB4",
    x"3F4B6085",
    x"3F4B6456",
    x"3F4B6827",
    x"3F4B6BF7",
    x"3F4B6FC8",
    x"3F4B7398",
    x"3F4B7768",
    x"3F4B7B39",
    x"3F4B7F09",
    x"3F4B82D8",
    x"3F4B86A8",
    x"3F4B8A78",
    x"3F4B8E47",
    x"3F4B9217",
    x"3F4B95E6",
    x"3F4B99B5",
    x"3F4B9D84",
    x"3F4BA153",
    x"3F4BA522",
    x"3F4BA8F0",
    x"3F4BACBF",
    x"3F4BB08D",
    x"3F4BB45B",
    x"3F4BB82A",
    x"3F4BBBF8",
    x"3F4BBFC6",
    x"3F4BC393",
    x"3F4BC761",
    x"3F4BCB2F",
    x"3F4BCEFC",
    x"3F4BD2C9",
    x"3F4BD696",
    x"3F4BDA63",
    x"3F4BDE30",
    x"3F4BE1FD",
    x"3F4BE5CA",
    x"3F4BE996",
    x"3F4BED63",
    x"3F4BF12F",
    x"3F4BF4FB",
    x"3F4BF8C7",
    x"3F4BFC93",
    x"3F4C005F",
    x"3F4C042B",
    x"3F4C07F6",
    x"3F4C0BC2",
    x"3F4C0F8D",
    x"3F4C1358",
    x"3F4C1723",
    x"3F4C1AEE",
    x"3F4C1EB9",
    x"3F4C2284",
    x"3F4C264E",
    x"3F4C2A19",
    x"3F4C2DE3",
    x"3F4C31AD",
    x"3F4C3578",
    x"3F4C3942",
    x"3F4C3D0B",
    x"3F4C40D5",
    x"3F4C449F",
    x"3F4C4868",
    x"3F4C4C32",
    x"3F4C4FFB",
    x"3F4C53C4",
    x"3F4C578D",
    x"3F4C5B56",
    x"3F4C5F1E",
    x"3F4C62E7",
    x"3F4C66B0",
    x"3F4C6A78",
    x"3F4C6E40",
    x"3F4C7208",
    x"3F4C75D0",
    x"3F4C7998",
    x"3F4C7D60",
    x"3F4C8128",
    x"3F4C84EF",
    x"3F4C88B6",
    x"3F4C8C7E",
    x"3F4C9045",
    x"3F4C940C",
    x"3F4C97D3",
    x"3F4C9B99",
    x"3F4C9F60",
    x"3F4CA327",
    x"3F4CA6ED",
    x"3F4CAAB3",
    x"3F4CAE79",
    x"3F4CB23F",
    x"3F4CB605",
    x"3F4CB9CB",
    x"3F4CBD91",
    x"3F4CC156",
    x"3F4CC51C",
    x"3F4CC8E1",
    x"3F4CCCA6",
    x"3F4CD06B",
    x"3F4CD430",
    x"3F4CD7F5",
    x"3F4CDBBA",
    x"3F4CDF7E",
    x"3F4CE343",
    x"3F4CE707",
    x"3F4CEACB",
    x"3F4CEE8F",
    x"3F4CF253",
    x"3F4CF617",
    x"3F4CF9DB",
    x"3F4CFD9E",
    x"3F4D0162",
    x"3F4D0525",
    x"3F4D08E8",
    x"3F4D0CAB",
    x"3F4D106E",
    x"3F4D1431",
    x"3F4D17F4",
    x"3F4D1BB6",
    x"3F4D1F79",
    x"3F4D233B",
    x"3F4D26FD",
    x"3F4D2ABF",
    x"3F4D2E81",
    x"3F4D3243",
    x"3F4D3605",
    x"3F4D39C6",
    x"3F4D3D88",
    x"3F4D4149",
    x"3F4D450A",
    x"3F4D48CB",
    x"3F4D4C8C",
    x"3F4D504D",
    x"3F4D540E",
    x"3F4D57CE",
    x"3F4D5B8F",
    x"3F4D5F4F",
    x"3F4D6310",
    x"3F4D66D0",
    x"3F4D6A90",
    x"3F4D6E4F",
    x"3F4D720F",
    x"3F4D75CF",
    x"3F4D798E",
    x"3F4D7D4E",
    x"3F4D810D",
    x"3F4D84CC",
    x"3F4D888B",
    x"3F4D8C4A",
    x"3F4D9009",
    x"3F4D93C7",
    x"3F4D9786",
    x"3F4D9B44",
    x"3F4D9F02",
    x"3F4DA2C0",
    x"3F4DA67E",
    x"3F4DAA3C",
    x"3F4DADFA",
    x"3F4DB1B8",
    x"3F4DB575",
    x"3F4DB932",
    x"3F4DBCF0",
    x"3F4DC0AD",
    x"3F4DC46A",
    x"3F4DC827",
    x"3F4DCBE3",
    x"3F4DCFA0",
    x"3F4DD35D",
    x"3F4DD719",
    x"3F4DDAD5",
    x"3F4DDE91",
    x"3F4DE24D",
    x"3F4DE609",
    x"3F4DE9C5",
    x"3F4DED81",
    x"3F4DF13C",
    x"3F4DF4F8",
    x"3F4DF8B3",
    x"3F4DFC6E",
    x"3F4E0029",
    x"3F4E03E4",
    x"3F4E079F",
    x"3F4E0B59",
    x"3F4E0F14",
    x"3F4E12CE",
    x"3F4E1689",
    x"3F4E1A43",
    x"3F4E1DFD",
    x"3F4E21B7",
    x"3F4E2570",
    x"3F4E292A",
    x"3F4E2CE4",
    x"3F4E309D",
    x"3F4E3456",
    x"3F4E380F",
    x"3F4E3BC8",
    x"3F4E3F81",
    x"3F4E433A",
    x"3F4E46F3",
    x"3F4E4AAB",
    x"3F4E4E64",
    x"3F4E521C",
    x"3F4E55D4",
    x"3F4E598C",
    x"3F4E5D44",
    x"3F4E60FC",
    x"3F4E64B4",
    x"3F4E686B",
    x"3F4E6C23",
    x"3F4E6FDA",
    x"3F4E7391",
    x"3F4E7748",
    x"3F4E7AFF",
    x"3F4E7EB6",
    x"3F4E826C",
    x"3F4E8623",
    x"3F4E89D9",
    x"3F4E8D90",
    x"3F4E9146",
    x"3F4E94FC",
    x"3F4E98B2",
    x"3F4E9C68",
    x"3F4EA01D",
    x"3F4EA3D3",
    x"3F4EA788",
    x"3F4EAB3E",
    x"3F4EAEF3",
    x"3F4EB2A8",
    x"3F4EB65D",
    x"3F4EBA12",
    x"3F4EBDC6",
    x"3F4EC17B",
    x"3F4EC52F",
    x"3F4EC8E4",
    x"3F4ECC98",
    x"3F4ED04C",
    x"3F4ED400",
    x"3F4ED7B3",
    x"3F4EDB67",
    x"3F4EDF1B",
    x"3F4EE2CE",
    x"3F4EE681",
    x"3F4EEA35",
    x"3F4EEDE8",
    x"3F4EF19B",
    x"3F4EF54D",
    x"3F4EF900",
    x"3F4EFCB3",
    x"3F4F0065",
    x"3F4F0417",
    x"3F4F07CA",
    x"3F4F0B7C",
    x"3F4F0F2E",
    x"3F4F12DF",
    x"3F4F1691",
    x"3F4F1A43",
    x"3F4F1DF4",
    x"3F4F21A5",
    x"3F4F2557",
    x"3F4F2908",
    x"3F4F2CB9",
    x"3F4F3069",
    x"3F4F341A",
    x"3F4F37CB",
    x"3F4F3B7B",
    x"3F4F3F2B",
    x"3F4F42DC",
    x"3F4F468C",
    x"3F4F4A3C",
    x"3F4F4DEB",
    x"3F4F519B",
    x"3F4F554B",
    x"3F4F58FA",
    x"3F4F5CA9",
    x"3F4F6059",
    x"3F4F6408",
    x"3F4F67B7",
    x"3F4F6B65",
    x"3F4F6F14",
    x"3F4F72C3",
    x"3F4F7671",
    x"3F4F7A1F",
    x"3F4F7DCE",
    x"3F4F817C",
    x"3F4F852A",
    x"3F4F88D7",
    x"3F4F8C85",
    x"3F4F9033",
    x"3F4F93E0",
    x"3F4F978D",
    x"3F4F9B3B",
    x"3F4F9EE8",
    x"3F4FA295",
    x"3F4FA642",
    x"3F4FA9EE",
    x"3F4FAD9B",
    x"3F4FB147",
    x"3F4FB4F4",
    x"3F4FB8A0",
    x"3F4FBC4C",
    x"3F4FBFF8",
    x"3F4FC3A4",
    x"3F4FC74F",
    x"3F4FCAFB",
    x"3F4FCEA6",
    x"3F4FD252",
    x"3F4FD5FD",
    x"3F4FD9A8",
    x"3F4FDD53",
    x"3F4FE0FE",
    x"3F4FE4A8",
    x"3F4FE853",
    x"3F4FEBFD",
    x"3F4FEFA8",
    x"3F4FF352",
    x"3F4FF6FC",
    x"3F4FFAA6",
    x"3F4FFE50",
    x"3F5001F9",
    x"3F5005A3",
    x"3F50094C",
    x"3F500CF6",
    x"3F50109F",
    x"3F501448",
    x"3F5017F1",
    x"3F501B9A",
    x"3F501F42",
    x"3F5022EB",
    x"3F502693",
    x"3F502A3B",
    x"3F502DE4",
    x"3F50318C",
    x"3F503534",
    x"3F5038DB",
    x"3F503C83",
    x"3F50402B",
    x"3F5043D2",
    x"3F504779",
    x"3F504B21",
    x"3F504EC8",
    x"3F50526F",
    x"3F505615",
    x"3F5059BC",
    x"3F505D63",
    x"3F506109",
    x"3F5064AF",
    x"3F506856",
    x"3F506BFC",
    x"3F506FA1",
    x"3F507347",
    x"3F5076ED",
    x"3F507A92",
    x"3F507E38",
    x"3F5081DD",
    x"3F508582",
    x"3F508927",
    x"3F508CCC",
    x"3F509071",
    x"3F509416",
    x"3F5097BA",
    x"3F509B5F",
    x"3F509F03",
    x"3F50A2A7",
    x"3F50A64B",
    x"3F50A9EF",
    x"3F50AD93",
    x"3F50B137",
    x"3F50B4DA",
    x"3F50B87E",
    x"3F50BC21",
    x"3F50BFC4",
    x"3F50C367",
    x"3F50C70A",
    x"3F50CAAD",
    x"3F50CE4F",
    x"3F50D1F2",
    x"3F50D594",
    x"3F50D937",
    x"3F50DCD9",
    x"3F50E07B",
    x"3F50E41D",
    x"3F50E7BE",
    x"3F50EB60",
    x"3F50EF02",
    x"3F50F2A3",
    x"3F50F644",
    x"3F50F9E5",
    x"3F50FD86",
    x"3F510127",
    x"3F5104C8",
    x"3F510869",
    x"3F510C09",
    x"3F510FAA",
    x"3F51134A",
    x"3F5116EA",
    x"3F511A8A",
    x"3F511E2A",
    x"3F5121CA",
    x"3F512569",
    x"3F512909",
    x"3F512CA8",
    x"3F513047",
    x"3F5133E7",
    x"3F513786",
    x"3F513B25",
    x"3F513EC3",
    x"3F514262",
    x"3F514600",
    x"3F51499F",
    x"3F514D3D",
    x"3F5150DB",
    x"3F515479",
    x"3F515817",
    x"3F515BB5",
    x"3F515F52",
    x"3F5162F0",
    x"3F51668D",
    x"3F516A2A",
    x"3F516DC8",
    x"3F517165",
    x"3F517501",
    x"3F51789E",
    x"3F517C3B",
    x"3F517FD7",
    x"3F518374",
    x"3F518710",
    x"3F518AAC",
    x"3F518E48",
    x"3F5191E4",
    x"3F51957F",
    x"3F51991B",
    x"3F519CB7",
    x"3F51A052",
    x"3F51A3ED",
    x"3F51A788",
    x"3F51AB23",
    x"3F51AEBE",
    x"3F51B259",
    x"3F51B5F3",
    x"3F51B98E",
    x"3F51BD28",
    x"3F51C0C2",
    x"3F51C45C",
    x"3F51C7F6",
    x"3F51CB90",
    x"3F51CF2A",
    x"3F51D2C3",
    x"3F51D65D",
    x"3F51D9F6",
    x"3F51DD8F",
    x"3F51E129",
    x"3F51E4C1",
    x"3F51E85A",
    x"3F51EBF3",
    x"3F51EF8C",
    x"3F51F324",
    x"3F51F6BC",
    x"3F51FA54",
    x"3F51FDED",
    x"3F520184",
    x"3F52051C",
    x"3F5208B4",
    x"3F520C4C",
    x"3F520FE3",
    x"3F52137A",
    x"3F521711",
    x"3F521AA8",
    x"3F521E3F",
    x"3F5221D6",
    x"3F52256D",
    x"3F522903",
    x"3F522C9A",
    x"3F523030",
    x"3F5233C6",
    x"3F52375C",
    x"3F523AF2",
    x"3F523E88",
    x"3F52421E",
    x"3F5245B3",
    x"3F524949",
    x"3F524CDE",
    x"3F525073",
    x"3F525408",
    x"3F52579D",
    x"3F525B32",
    x"3F525EC6",
    x"3F52625B",
    x"3F5265EF",
    x"3F526983",
    x"3F526D18",
    x"3F5270AC",
    x"3F52743F",
    x"3F5277D3",
    x"3F527B67",
    x"3F527EFA",
    x"3F52828E",
    x"3F528621",
    x"3F5289B4",
    x"3F528D47",
    x"3F5290DA",
    x"3F52946D",
    x"3F5297FF",
    x"3F529B92",
    x"3F529F24",
    x"3F52A2B6",
    x"3F52A649",
    x"3F52A9DA",
    x"3F52AD6C",
    x"3F52B0FE",
    x"3F52B490",
    x"3F52B821",
    x"3F52BBB2",
    x"3F52BF44",
    x"3F52C2D5",
    x"3F52C666",
    x"3F52C9F7",
    x"3F52CD87",
    x"3F52D118",
    x"3F52D4A8",
    x"3F52D839",
    x"3F52DBC9",
    x"3F52DF59",
    x"3F52E2E9",
    x"3F52E679",
    x"3F52EA08",
    x"3F52ED98",
    x"3F52F127",
    x"3F52F4B7",
    x"3F52F846",
    x"3F52FBD5",
    x"3F52FF64",
    x"3F5302F3",
    x"3F530681",
    x"3F530A10",
    x"3F530D9E",
    x"3F53112D",
    x"3F5314BB",
    x"3F531849",
    x"3F531BD7",
    x"3F531F65",
    x"3F5322F2",
    x"3F532680",
    x"3F532A0D",
    x"3F532D9A",
    x"3F533128",
    x"3F5334B5",
    x"3F533841",
    x"3F533BCE",
    x"3F533F5B",
    x"3F5342E7",
    x"3F534674",
    x"3F534A00",
    x"3F534D8C",
    x"3F535118",
    x"3F5354A4",
    x"3F535830",
    x"3F535BBB",
    x"3F535F47",
    x"3F5362D2",
    x"3F53665E",
    x"3F5369E9",
    x"3F536D74",
    x"3F5370FF",
    x"3F537489",
    x"3F537814",
    x"3F537B9E",
    x"3F537F29",
    x"3F5382B3",
    x"3F53863D",
    x"3F5389C7",
    x"3F538D51",
    x"3F5390DB",
    x"3F539464",
    x"3F5397EE",
    x"3F539B77",
    x"3F539F00",
    x"3F53A289",
    x"3F53A612",
    x"3F53A99B",
    x"3F53AD24",
    x"3F53B0AC",
    x"3F53B435",
    x"3F53B7BD",
    x"3F53BB45",
    x"3F53BECD",
    x"3F53C255",
    x"3F53C5DD",
    x"3F53C965",
    x"3F53CCEC",
    x"3F53D074",
    x"3F53D3FB",
    x"3F53D782",
    x"3F53DB09",
    x"3F53DE90",
    x"3F53E217",
    x"3F53E59D",
    x"3F53E924",
    x"3F53ECAA",
    x"3F53F031",
    x"3F53F3B7",
    x"3F53F73D",
    x"3F53FAC3",
    x"3F53FE48",
    x"3F5401CE",
    x"3F540553",
    x"3F5408D9",
    x"3F540C5E",
    x"3F540FE3",
    x"3F541368",
    x"3F5416ED",
    x"3F541A72",
    x"3F541DF6",
    x"3F54217B",
    x"3F5424FF",
    x"3F542883",
    x"3F542C08",
    x"3F542F8C",
    x"3F54330F",
    x"3F543693",
    x"3F543A17",
    x"3F543D9A",
    x"3F54411D",
    x"3F5444A1",
    x"3F544824",
    x"3F544BA7",
    x"3F544F2A",
    x"3F5452AC",
    x"3F54562F",
    x"3F5459B1",
    x"3F545D33",
    x"3F5460B6",
    x"3F546438",
    x"3F5467BA",
    x"3F546B3B",
    x"3F546EBD",
    x"3F54723F",
    x"3F5475C0",
    x"3F547941",
    x"3F547CC3",
    x"3F548044",
    x"3F5483C4",
    x"3F548745",
    x"3F548AC6",
    x"3F548E46",
    x"3F5491C7",
    x"3F549547",
    x"3F5498C7",
    x"3F549C47",
    x"3F549FC7",
    x"3F54A347",
    x"3F54A6C6",
    x"3F54AA46",
    x"3F54ADC5",
    x"3F54B144",
    x"3F54B4C4",
    x"3F54B843",
    x"3F54BBC1",
    x"3F54BF40",
    x"3F54C2BF",
    x"3F54C63D",
    x"3F54C9BC",
    x"3F54CD3A",
    x"3F54D0B8",
    x"3F54D436",
    x"3F54D7B4",
    x"3F54DB31",
    x"3F54DEAF",
    x"3F54E22C",
    x"3F54E5AA",
    x"3F54E927",
    x"3F54ECA4",
    x"3F54F021",
    x"3F54F39E",
    x"3F54F71A",
    x"3F54FA97",
    x"3F54FE13",
    x"3F55018F",
    x"3F55050C",
    x"3F550888",
    x"3F550C04",
    x"3F550F7F",
    x"3F5512FB",
    x"3F551676",
    x"3F5519F2",
    x"3F551D6D",
    x"3F5520E8",
    x"3F552463",
    x"3F5527DE",
    x"3F552B59",
    x"3F552ED4",
    x"3F55324E",
    x"3F5535C8",
    x"3F553943",
    x"3F553CBD",
    x"3F554037",
    x"3F5543B1",
    x"3F55472A",
    x"3F554AA4",
    x"3F554E1D",
    x"3F555197",
    x"3F555510",
    x"3F555889",
    x"3F555C02",
    x"3F555F7B",
    x"3F5562F3",
    x"3F55666C",
    x"3F5569E4",
    x"3F556D5D",
    x"3F5570D5",
    x"3F55744D",
    x"3F5577C5",
    x"3F557B3D",
    x"3F557EB4",
    x"3F55822C",
    x"3F5585A3",
    x"3F55891A",
    x"3F558C92",
    x"3F559009",
    x"3F55937F",
    x"3F5596F6",
    x"3F559A6D",
    x"3F559DE3",
    x"3F55A15A",
    x"3F55A4D0",
    x"3F55A846",
    x"3F55ABBC",
    x"3F55AF32",
    x"3F55B2A8",
    x"3F55B61D",
    x"3F55B993",
    x"3F55BD08",
    x"3F55C07D",
    x"3F55C3F2",
    x"3F55C767",
    x"3F55CADC",
    x"3F55CE51",
    x"3F55D1C5",
    x"3F55D53A",
    x"3F55D8AE",
    x"3F55DC22",
    x"3F55DF96",
    x"3F55E30A",
    x"3F55E67E",
    x"3F55E9F2",
    x"3F55ED65",
    x"3F55F0D9",
    x"3F55F44C",
    x"3F55F7BF",
    x"3F55FB32",
    x"3F55FEA5",
    x"3F560218",
    x"3F56058B",
    x"3F5608FD",
    x"3F560C70",
    x"3F560FE2",
    x"3F561354",
    x"3F5616C6",
    x"3F561A38",
    x"3F561DA9",
    x"3F56211B",
    x"3F56248D",
    x"3F5627FE",
    x"3F562B6F",
    x"3F562EE0",
    x"3F563251",
    x"3F5635C2",
    x"3F563933",
    x"3F563CA3",
    x"3F564014",
    x"3F564384",
    x"3F5646F4",
    x"3F564A64",
    x"3F564DD4",
    x"3F565144",
    x"3F5654B4",
    x"3F565823",
    x"3F565B93",
    x"3F565F02",
    x"3F566271",
    x"3F5665E0",
    x"3F56694F",
    x"3F566CBE",
    x"3F56702C",
    x"3F56739B",
    x"3F567709",
    x"3F567A78",
    x"3F567DE6",
    x"3F568154",
    x"3F5684C2",
    x"3F56882F",
    x"3F568B9D",
    x"3F568F0A",
    x"3F569278",
    x"3F5695E5",
    x"3F569952",
    x"3F569CBF",
    x"3F56A02C",
    x"3F56A399",
    x"3F56A705",
    x"3F56AA72",
    x"3F56ADDE",
    x"3F56B14A",
    x"3F56B4B6",
    x"3F56B822",
    x"3F56BB8E",
    x"3F56BEF9",
    x"3F56C265",
    x"3F56C5D0",
    x"3F56C93C",
    x"3F56CCA7",
    x"3F56D012",
    x"3F56D37D",
    x"3F56D6E8",
    x"3F56DA52",
    x"3F56DDBD",
    x"3F56E127",
    x"3F56E491",
    x"3F56E7FB",
    x"3F56EB65",
    x"3F56EECF",
    x"3F56F239",
    x"3F56F5A3",
    x"3F56F90C",
    x"3F56FC75",
    x"3F56FFDF",
    x"3F570348",
    x"3F5706B1",
    x"3F570A19",
    x"3F570D82",
    x"3F5710EB",
    x"3F571453",
    x"3F5717BB",
    x"3F571B24",
    x"3F571E8C",
    x"3F5721F3",
    x"3F57255B",
    x"3F5728C3",
    x"3F572C2A",
    x"3F572F92",
    x"3F5732F9",
    x"3F573660",
    x"3F5739C7",
    x"3F573D2E",
    x"3F574095",
    x"3F5743FB",
    x"3F574762",
    x"3F574AC8",
    x"3F574E2F",
    x"3F575195",
    x"3F5754FB",
    x"3F575860",
    x"3F575BC6",
    x"3F575F2C",
    x"3F576291",
    x"3F5765F6",
    x"3F57695C",
    x"3F576CC1",
    x"3F577026",
    x"3F57738A",
    x"3F5776EF",
    x"3F577A54",
    x"3F577DB8",
    x"3F57811C",
    x"3F578480",
    x"3F5787E4",
    x"3F578B48",
    x"3F578EAC",
    x"3F579210",
    x"3F579573",
    x"3F5798D7",
    x"3F579C3A",
    x"3F579F9D",
    x"3F57A300",
    x"3F57A663",
    x"3F57A9C6",
    x"3F57AD28",
    x"3F57B08B",
    x"3F57B3ED",
    x"3F57B74F",
    x"3F57BAB1",
    x"3F57BE13",
    x"3F57C175",
    x"3F57C4D7",
    x"3F57C838",
    x"3F57CB9A",
    x"3F57CEFB",
    x"3F57D25C",
    x"3F57D5BD",
    x"3F57D91E",
    x"3F57DC7F",
    x"3F57DFDF",
    x"3F57E340",
    x"3F57E6A0",
    x"3F57EA01",
    x"3F57ED61",
    x"3F57F0C1",
    x"3F57F421",
    x"3F57F780",
    x"3F57FAE0",
    x"3F57FE3F",
    x"3F58019F",
    x"3F5804FE",
    x"3F58085D",
    x"3F580BBC",
    x"3F580F1B",
    x"3F581279",
    x"3F5815D8",
    x"3F581936",
    x"3F581C95",
    x"3F581FF3",
    x"3F582351",
    x"3F5826AF",
    x"3F582A0D",
    x"3F582D6A",
    x"3F5830C8",
    x"3F583425",
    x"3F583782",
    x"3F583AE0",
    x"3F583E3D",
    x"3F584199",
    x"3F5844F6",
    x"3F584853",
    x"3F584BAF",
    x"3F584F0C",
    x"3F585268",
    x"3F5855C4",
    x"3F585920",
    x"3F585C7C",
    x"3F585FD7",
    x"3F586333",
    x"3F58668E",
    x"3F5869EA",
    x"3F586D45",
    x"3F5870A0",
    x"3F5873FB",
    x"3F587756",
    x"3F587AB0",
    x"3F587E0B",
    x"3F588165",
    x"3F5884BF",
    x"3F58881A",
    x"3F588B74",
    x"3F588ECD",
    x"3F589227",
    x"3F589581",
    x"3F5898DA",
    x"3F589C34",
    x"3F589F8D",
    x"3F58A2E6",
    x"3F58A63F",
    x"3F58A998",
    x"3F58ACF0",
    x"3F58B049",
    x"3F58B3A1",
    x"3F58B6FA",
    x"3F58BA52",
    x"3F58BDAA",
    x"3F58C102",
    x"3F58C45A",
    x"3F58C7B1",
    x"3F58CB09",
    x"3F58CE60",
    x"3F58D1B7",
    x"3F58D50E",
    x"3F58D865",
    x"3F58DBBC",
    x"3F58DF13",
    x"3F58E26A",
    x"3F58E5C0",
    x"3F58E916",
    x"3F58EC6D",
    x"3F58EFC3",
    x"3F58F319",
    x"3F58F66F",
    x"3F58F9C4",
    x"3F58FD1A",
    x"3F59006F",
    x"3F5903C5",
    x"3F59071A",
    x"3F590A6F",
    x"3F590DC4",
    x"3F591118",
    x"3F59146D",
    x"3F5917C2",
    x"3F591B16",
    x"3F591E6A",
    x"3F5921BE",
    x"3F592512",
    x"3F592866",
    x"3F592BBA",
    x"3F592F0E",
    x"3F593261",
    x"3F5935B4",
    x"3F593908",
    x"3F593C5B",
    x"3F593FAE",
    x"3F594300",
    x"3F594653",
    x"3F5949A6",
    x"3F594CF8",
    x"3F59504A",
    x"3F59539C",
    x"3F5956EE",
    x"3F595A40",
    x"3F595D92",
    x"3F5960E4",
    x"3F596435",
    x"3F596787",
    x"3F596AD8",
    x"3F596E29",
    x"3F59717A",
    x"3F5974CB",
    x"3F59781C",
    x"3F597B6C",
    x"3F597EBD",
    x"3F59820D",
    x"3F59855D",
    x"3F5988AD",
    x"3F598BFD",
    x"3F598F4D",
    x"3F59929D",
    x"3F5995EC",
    x"3F59993C",
    x"3F599C8B",
    x"3F599FDA",
    x"3F59A329",
    x"3F59A678",
    x"3F59A9C7",
    x"3F59AD15",
    x"3F59B064",
    x"3F59B3B2",
    x"3F59B700",
    x"3F59BA4E",
    x"3F59BD9C",
    x"3F59C0EA",
    x"3F59C438",
    x"3F59C785",
    x"3F59CAD3",
    x"3F59CE20",
    x"3F59D16D",
    x"3F59D4BA",
    x"3F59D807",
    x"3F59DB54",
    x"3F59DEA1",
    x"3F59E1ED",
    x"3F59E53A",
    x"3F59E886",
    x"3F59EBD2",
    x"3F59EF1E",
    x"3F59F26A",
    x"3F59F5B6",
    x"3F59F901",
    x"3F59FC4D",
    x"3F59FF98",
    x"3F5A02E3",
    x"3F5A062E",
    x"3F5A0979",
    x"3F5A0CC4",
    x"3F5A100F",
    x"3F5A1359",
    x"3F5A16A4",
    x"3F5A19EE",
    x"3F5A1D38",
    x"3F5A2082",
    x"3F5A23CC",
    x"3F5A2716",
    x"3F5A2A60",
    x"3F5A2DA9",
    x"3F5A30F2",
    x"3F5A343C",
    x"3F5A3785",
    x"3F5A3ACE",
    x"3F5A3E17",
    x"3F5A415F",
    x"3F5A44A8",
    x"3F5A47F0",
    x"3F5A4B39",
    x"3F5A4E81",
    x"3F5A51C9",
    x"3F5A5511",
    x"3F5A5859",
    x"3F5A5BA0",
    x"3F5A5EE8",
    x"3F5A622F",
    x"3F5A6577",
    x"3F5A68BE",
    x"3F5A6C05",
    x"3F5A6F4C",
    x"3F5A7292",
    x"3F5A75D9",
    x"3F5A791F",
    x"3F5A7C66",
    x"3F5A7FAC",
    x"3F5A82F2",
    x"3F5A8638",
    x"3F5A897E",
    x"3F5A8CC3",
    x"3F5A9009",
    x"3F5A934E",
    x"3F5A9694",
    x"3F5A99D9",
    x"3F5A9D1E",
    x"3F5AA063",
    x"3F5AA3A8",
    x"3F5AA6EC",
    x"3F5AAA31",
    x"3F5AAD75",
    x"3F5AB0B9",
    x"3F5AB3FD",
    x"3F5AB741",
    x"3F5ABA85",
    x"3F5ABDC9",
    x"3F5AC10D",
    x"3F5AC450",
    x"3F5AC793",
    x"3F5ACAD6",
    x"3F5ACE1A",
    x"3F5AD15C",
    x"3F5AD49F",
    x"3F5AD7E2",
    x"3F5ADB24",
    x"3F5ADE67",
    x"3F5AE1A9",
    x"3F5AE4EB",
    x"3F5AE82D",
    x"3F5AEB6F",
    x"3F5AEEB1",
    x"3F5AF1F2",
    x"3F5AF534",
    x"3F5AF875",
    x"3F5AFBB6",
    x"3F5AFEF7",
    x"3F5B0238",
    x"3F5B0579",
    x"3F5B08BA",
    x"3F5B0BFA",
    x"3F5B0F3B",
    x"3F5B127B",
    x"3F5B15BB",
    x"3F5B18FB",
    x"3F5B1C3B",
    x"3F5B1F7B",
    x"3F5B22BB",
    x"3F5B25FA",
    x"3F5B2939",
    x"3F5B2C79",
    x"3F5B2FB8",
    x"3F5B32F7",
    x"3F5B3636",
    x"3F5B3974",
    x"3F5B3CB3",
    x"3F5B3FF1",
    x"3F5B4330",
    x"3F5B466E",
    x"3F5B49AC",
    x"3F5B4CEA",
    x"3F5B5027",
    x"3F5B5365",
    x"3F5B56A3",
    x"3F5B59E0",
    x"3F5B5D1D",
    x"3F5B605A",
    x"3F5B6397",
    x"3F5B66D4",
    x"3F5B6A11",
    x"3F5B6D4D",
    x"3F5B708A",
    x"3F5B73C6",
    x"3F5B7702",
    x"3F5B7A3E",
    x"3F5B7D7A",
    x"3F5B80B6",
    x"3F5B83F2",
    x"3F5B872D",
    x"3F5B8A69",
    x"3F5B8DA4",
    x"3F5B90DF",
    x"3F5B941A",
    x"3F5B9755",
    x"3F5B9A90",
    x"3F5B9DCA",
    x"3F5BA105",
    x"3F5BA43F",
    x"3F5BA779",
    x"3F5BAAB3",
    x"3F5BADED",
    x"3F5BB127",
    x"3F5BB461",
    x"3F5BB79A",
    x"3F5BBAD4",
    x"3F5BBE0D",
    x"3F5BC146",
    x"3F5BC47F",
    x"3F5BC7B8",
    x"3F5BCAF1",
    x"3F5BCE29",
    x"3F5BD162",
    x"3F5BD49A",
    x"3F5BD7D3",
    x"3F5BDB0B",
    x"3F5BDE43",
    x"3F5BE17A",
    x"3F5BE4B2",
    x"3F5BE7EA",
    x"3F5BEB21",
    x"3F5BEE58",
    x"3F5BF190",
    x"3F5BF4C7",
    x"3F5BF7FD",
    x"3F5BFB34",
    x"3F5BFE6B",
    x"3F5C01A1",
    x"3F5C04D8",
    x"3F5C080E",
    x"3F5C0B44",
    x"3F5C0E7A",
    x"3F5C11B0",
    x"3F5C14E6",
    x"3F5C181B",
    x"3F5C1B51",
    x"3F5C1E86",
    x"3F5C21BB",
    x"3F5C24F0",
    x"3F5C2825",
    x"3F5C2B5A",
    x"3F5C2E8E",
    x"3F5C31C3",
    x"3F5C34F7",
    x"3F5C382B",
    x"3F5C3B60",
    x"3F5C3E94",
    x"3F5C41C7",
    x"3F5C44FB",
    x"3F5C482F",
    x"3F5C4B62",
    x"3F5C4E95",
    x"3F5C51C9",
    x"3F5C54FC",
    x"3F5C582F",
    x"3F5C5B61",
    x"3F5C5E94",
    x"3F5C61C7",
    x"3F5C64F9",
    x"3F5C682B",
    x"3F5C6B5D",
    x"3F5C6E8F",
    x"3F5C71C1",
    x"3F5C74F3",
    x"3F5C7824",
    x"3F5C7B56",
    x"3F5C7E87",
    x"3F5C81B8",
    x"3F5C84EA",
    x"3F5C881A",
    x"3F5C8B4B",
    x"3F5C8E7C",
    x"3F5C91AC",
    x"3F5C94DD",
    x"3F5C980D",
    x"3F5C9B3D",
    x"3F5C9E6D",
    x"3F5CA19D",
    x"3F5CA4CD",
    x"3F5CA7FC",
    x"3F5CAB2C",
    x"3F5CAE5B",
    x"3F5CB18A",
    x"3F5CB4B9",
    x"3F5CB7E8",
    x"3F5CBB17",
    x"3F5CBE46",
    x"3F5CC174",
    x"3F5CC4A3",
    x"3F5CC7D1",
    x"3F5CCAFF",
    x"3F5CCE2D",
    x"3F5CD15B",
    x"3F5CD489",
    x"3F5CD7B6",
    x"3F5CDAE4",
    x"3F5CDE11",
    x"3F5CE13E",
    x"3F5CE46B",
    x"3F5CE798",
    x"3F5CEAC5",
    x"3F5CEDF2",
    x"3F5CF11E",
    x"3F5CF44B",
    x"3F5CF777",
    x"3F5CFAA3",
    x"3F5CFDCF",
    x"3F5D00FB",
    x"3F5D0427",
    x"3F5D0752",
    x"3F5D0A7E",
    x"3F5D0DA9",
    x"3F5D10D4",
    x"3F5D13FF",
    x"3F5D172A",
    x"3F5D1A55",
    x"3F5D1D80",
    x"3F5D20AA",
    x"3F5D23D5",
    x"3F5D26FF",
    x"3F5D2A29",
    x"3F5D2D53",
    x"3F5D307D",
    x"3F5D33A7",
    x"3F5D36D0",
    x"3F5D39FA",
    x"3F5D3D23",
    x"3F5D404C",
    x"3F5D4376",
    x"3F5D469E",
    x"3F5D49C7",
    x"3F5D4CF0",
    x"3F5D5018",
    x"3F5D5341",
    x"3F5D5669",
    x"3F5D5991",
    x"3F5D5CB9",
    x"3F5D5FE1",
    x"3F5D6309",
    x"3F5D6631",
    x"3F5D6958",
    x"3F5D6C7F",
    x"3F5D6FA7",
    x"3F5D72CE",
    x"3F5D75F5",
    x"3F5D791B",
    x"3F5D7C42",
    x"3F5D7F69",
    x"3F5D828F",
    x"3F5D85B5",
    x"3F5D88DB",
    x"3F5D8C01",
    x"3F5D8F27",
    x"3F5D924D",
    x"3F5D9573",
    x"3F5D9898",
    x"3F5D9BBD",
    x"3F5D9EE3",
    x"3F5DA208",
    x"3F5DA52D",
    x"3F5DA851",
    x"3F5DAB76",
    x"3F5DAE9B",
    x"3F5DB1BF",
    x"3F5DB4E3",
    x"3F5DB807",
    x"3F5DBB2B",
    x"3F5DBE4F",
    x"3F5DC173",
    x"3F5DC497",
    x"3F5DC7BA",
    x"3F5DCADD",
    x"3F5DCE01",
    x"3F5DD124",
    x"3F5DD447",
    x"3F5DD769",
    x"3F5DDA8C",
    x"3F5DDDAF",
    x"3F5DE0D1",
    x"3F5DE3F3",
    x"3F5DE715",
    x"3F5DEA37",
    x"3F5DED59",
    x"3F5DF07B",
    x"3F5DF39D",
    x"3F5DF6BE",
    x"3F5DF9DF",
    x"3F5DFD01",
    x"3F5E0022",
    x"3F5E0343",
    x"3F5E0663",
    x"3F5E0984",
    x"3F5E0CA5",
    x"3F5E0FC5",
    x"3F5E12E5",
    x"3F5E1605",
    x"3F5E1925",
    x"3F5E1C45",
    x"3F5E1F65",
    x"3F5E2285",
    x"3F5E25A4",
    x"3F5E28C3",
    x"3F5E2BE3",
    x"3F5E2F02",
    x"3F5E3221",
    x"3F5E353F",
    x"3F5E385E",
    x"3F5E3B7D",
    x"3F5E3E9B",
    x"3F5E41B9",
    x"3F5E44D7",
    x"3F5E47F5",
    x"3F5E4B13",
    x"3F5E4E31",
    x"3F5E514E",
    x"3F5E546C",
    x"3F5E5789",
    x"3F5E5AA6",
    x"3F5E5DC3",
    x"3F5E60E0",
    x"3F5E63FD",
    x"3F5E671A",
    x"3F5E6A36",
    x"3F5E6D53",
    x"3F5E706F",
    x"3F5E738B",
    x"3F5E76A7",
    x"3F5E79C3",
    x"3F5E7CDE",
    x"3F5E7FFA",
    x"3F5E8316",
    x"3F5E8631",
    x"3F5E894C",
    x"3F5E8C67",
    x"3F5E8F82",
    x"3F5E929D",
    x"3F5E95B7",
    x"3F5E98D2",
    x"3F5E9BEC",
    x"3F5E9F06",
    x"3F5EA221",
    x"3F5EA53A",
    x"3F5EA854",
    x"3F5EAB6E",
    x"3F5EAE88",
    x"3F5EB1A1",
    x"3F5EB4BA",
    x"3F5EB7D3",
    x"3F5EBAEC",
    x"3F5EBE05",
    x"3F5EC11E",
    x"3F5EC437",
    x"3F5EC74F",
    x"3F5ECA68",
    x"3F5ECD80",
    x"3F5ED098",
    x"3F5ED3B0",
    x"3F5ED6C8",
    x"3F5ED9DF",
    x"3F5EDCF7",
    x"3F5EE00E",
    x"3F5EE326",
    x"3F5EE63D",
    x"3F5EE954",
    x"3F5EEC6B",
    x"3F5EEF81",
    x"3F5EF298",
    x"3F5EF5AE",
    x"3F5EF8C5",
    x"3F5EFBDB",
    x"3F5EFEF1",
    x"3F5F0207",
    x"3F5F051D",
    x"3F5F0833",
    x"3F5F0B48",
    x"3F5F0E5D",
    x"3F5F1173",
    x"3F5F1488",
    x"3F5F179D",
    x"3F5F1AB2",
    x"3F5F1DC6",
    x"3F5F20DB",
    x"3F5F23EF",
    x"3F5F2704",
    x"3F5F2A18",
    x"3F5F2D2C",
    x"3F5F3040",
    x"3F5F3354",
    x"3F5F3667",
    x"3F5F397B",
    x"3F5F3C8E",
    x"3F5F3FA2",
    x"3F5F42B5",
    x"3F5F45C8",
    x"3F5F48DB",
    x"3F5F4BED",
    x"3F5F4F00",
    x"3F5F5212",
    x"3F5F5525",
    x"3F5F5837",
    x"3F5F5B49",
    x"3F5F5E5B",
    x"3F5F616C",
    x"3F5F647E",
    x"3F5F6790",
    x"3F5F6AA1",
    x"3F5F6DB2",
    x"3F5F70C3",
    x"3F5F73D4",
    x"3F5F76E5",
    x"3F5F79F6",
    x"3F5F7D06",
    x"3F5F8017",
    x"3F5F8327",
    x"3F5F8637",
    x"3F5F8947",
    x"3F5F8C57",
    x"3F5F8F67",
    x"3F5F9276",
    x"3F5F9586",
    x"3F5F9895",
    x"3F5F9BA5",
    x"3F5F9EB4",
    x"3F5FA1C3",
    x"3F5FA4D1",
    x"3F5FA7E0",
    x"3F5FAAEF",
    x"3F5FADFD",
    x"3F5FB10B",
    x"3F5FB419",
    x"3F5FB727",
    x"3F5FBA35",
    x"3F5FBD43",
    x"3F5FC051",
    x"3F5FC35E",
    x"3F5FC66B",
    x"3F5FC979",
    x"3F5FCC86",
    x"3F5FCF93",
    x"3F5FD29F",
    x"3F5FD5AC",
    x"3F5FD8B8",
    x"3F5FDBC5",
    x"3F5FDED1",
    x"3F5FE1DD",
    x"3F5FE4E9",
    x"3F5FE7F5",
    x"3F5FEB01",
    x"3F5FEE0C",
    x"3F5FF118",
    x"3F5FF423",
    x"3F5FF72E",
    x"3F5FFA39",
    x"3F5FFD44",
    x"3F60004F",
    x"3F60035A",
    x"3F600664",
    x"3F60096E",
    x"3F600C79",
    x"3F600F83",
    x"3F60128D",
    x"3F601596",
    x"3F6018A0",
    x"3F601BAA",
    x"3F601EB3",
    x"3F6021BC",
    x"3F6024C6",
    x"3F6027CF",
    x"3F602AD7",
    x"3F602DE0",
    x"3F6030E9",
    x"3F6033F1",
    x"3F6036FA",
    x"3F603A02",
    x"3F603D0A",
    x"3F604012",
    x"3F60431A",
    x"3F604621",
    x"3F604929",
    x"3F604C30",
    x"3F604F37",
    x"3F60523E",
    x"3F605545",
    x"3F60584C",
    x"3F605B53",
    x"3F605E5A",
    x"3F606160",
    x"3F606466",
    x"3F60676D",
    x"3F606A73",
    x"3F606D78",
    x"3F60707E",
    x"3F607384",
    x"3F607689",
    x"3F60798F",
    x"3F607C94",
    x"3F607F99",
    x"3F60829E",
    x"3F6085A3",
    x"3F6088A7",
    x"3F608BAC",
    x"3F608EB0",
    x"3F6091B5",
    x"3F6094B9",
    x"3F6097BD",
    x"3F609AC1",
    x"3F609DC4",
    x"3F60A0C8",
    x"3F60A3CC",
    x"3F60A6CF",
    x"3F60A9D2",
    x"3F60ACD5",
    x"3F60AFD8",
    x"3F60B2DB",
    x"3F60B5DE",
    x"3F60B8E0",
    x"3F60BBE2",
    x"3F60BEE5",
    x"3F60C1E7",
    x"3F60C4E9",
    x"3F60C7EB",
    x"3F60CAEC",
    x"3F60CDEE",
    x"3F60D0EF",
    x"3F60D3F1",
    x"3F60D6F2",
    x"3F60D9F3",
    x"3F60DCF4",
    x"3F60DFF4",
    x"3F60E2F5",
    x"3F60E5F6",
    x"3F60E8F6",
    x"3F60EBF6",
    x"3F60EEF6",
    x"3F60F1F6",
    x"3F60F4F6",
    x"3F60F7F6",
    x"3F60FAF5",
    x"3F60FDF5",
    x"3F6100F4",
    x"3F6103F3",
    x"3F6106F2",
    x"3F6109F1",
    x"3F610CF0",
    x"3F610FEE",
    x"3F6112ED",
    x"3F6115EB",
    x"3F6118E9",
    x"3F611BE7",
    x"3F611EE5",
    x"3F6121E3",
    x"3F6124E1",
    x"3F6127DE",
    x"3F612ADB",
    x"3F612DD9",
    x"3F6130D6",
    x"3F6133D3",
    x"3F6136D0",
    x"3F6139CC",
    x"3F613CC9",
    x"3F613FC5",
    x"3F6142C1",
    x"3F6145BE",
    x"3F6148BA",
    x"3F614BB5",
    x"3F614EB1",
    x"3F6151AD",
    x"3F6154A8",
    x"3F6157A4",
    x"3F615A9F",
    x"3F615D9A",
    x"3F616095",
    x"3F616390",
    x"3F61668A",
    x"3F616985",
    x"3F616C7F",
    x"3F616F79",
    x"3F617274",
    x"3F61756E",
    x"3F617867",
    x"3F617B61",
    x"3F617E5B",
    x"3F618154",
    x"3F61844D",
    x"3F618747",
    x"3F618A40",
    x"3F618D38",
    x"3F619031",
    x"3F61932A",
    x"3F619622",
    x"3F61991B",
    x"3F619C13",
    x"3F619F0B",
    x"3F61A203",
    x"3F61A4FB",
    x"3F61A7F2",
    x"3F61AAEA",
    x"3F61ADE1",
    x"3F61B0D9",
    x"3F61B3D0",
    x"3F61B6C7",
    x"3F61B9BE",
    x"3F61BCB4",
    x"3F61BFAB",
    x"3F61C2A1",
    x"3F61C598",
    x"3F61C88E",
    x"3F61CB84",
    x"3F61CE7A",
    x"3F61D16F",
    x"3F61D465",
    x"3F61D75B",
    x"3F61DA50",
    x"3F61DD45",
    x"3F61E03A",
    x"3F61E32F",
    x"3F61E624",
    x"3F61E919",
    x"3F61EC0D",
    x"3F61EF02",
    x"3F61F1F6",
    x"3F61F4EA",
    x"3F61F7DE",
    x"3F61FAD2",
    x"3F61FDC6",
    x"3F6200B9",
    x"3F6203AD",
    x"3F6206A0",
    x"3F620993",
    x"3F620C86",
    x"3F620F79",
    x"3F62126C",
    x"3F62155E",
    x"3F621851",
    x"3F621B43",
    x"3F621E35",
    x"3F622128",
    x"3F62241A",
    x"3F62270B",
    x"3F6229FD",
    x"3F622CEF",
    x"3F622FE0",
    x"3F6232D1",
    x"3F6235C2",
    x"3F6238B3",
    x"3F623BA4",
    x"3F623E95",
    x"3F624186",
    x"3F624476",
    x"3F624766",
    x"3F624A57",
    x"3F624D47",
    x"3F625036",
    x"3F625326",
    x"3F625616",
    x"3F625905",
    x"3F625BF5",
    x"3F625EE4",
    x"3F6261D3",
    x"3F6264C2",
    x"3F6267B1",
    x"3F626AA0",
    x"3F626D8E",
    x"3F62707C",
    x"3F62736B",
    x"3F627659",
    x"3F627947",
    x"3F627C35",
    x"3F627F22",
    x"3F628210",
    x"3F6284FD",
    x"3F6287EB",
    x"3F628AD8",
    x"3F628DC5",
    x"3F6290B2",
    x"3F62939F",
    x"3F62968B",
    x"3F629978",
    x"3F629C64",
    x"3F629F50",
    x"3F62A23D",
    x"3F62A528",
    x"3F62A814",
    x"3F62AB00",
    x"3F62ADEB",
    x"3F62B0D7",
    x"3F62B3C2",
    x"3F62B6AD",
    x"3F62B998",
    x"3F62BC83",
    x"3F62BF6E",
    x"3F62C258",
    x"3F62C543",
    x"3F62C82D",
    x"3F62CB17",
    x"3F62CE01",
    x"3F62D0EB",
    x"3F62D3D5",
    x"3F62D6BF",
    x"3F62D9A8",
    x"3F62DC92",
    x"3F62DF7B",
    x"3F62E264",
    x"3F62E54D",
    x"3F62E836",
    x"3F62EB1E",
    x"3F62EE07",
    x"3F62F0EF",
    x"3F62F3D8",
    x"3F62F6C0",
    x"3F62F9A8",
    x"3F62FC8F",
    x"3F62FF77",
    x"3F63025F",
    x"3F630546",
    x"3F63082E",
    x"3F630B15",
    x"3F630DFC",
    x"3F6310E3",
    x"3F6313C9",
    x"3F6316B0",
    x"3F631996",
    x"3F631C7D",
    x"3F631F63",
    x"3F632249",
    x"3F63252F",
    x"3F632815",
    x"3F632AFB",
    x"3F632DE0",
    x"3F6330C5",
    x"3F6333AB",
    x"3F633690",
    x"3F633975",
    x"3F633C5A",
    x"3F633F3E",
    x"3F634223",
    x"3F634507",
    x"3F6347EC",
    x"3F634AD0",
    x"3F634DB4",
    x"3F635098",
    x"3F63537B",
    x"3F63565F",
    x"3F635943",
    x"3F635C26",
    x"3F635F09",
    x"3F6361EC",
    x"3F6364CF",
    x"3F6367B2",
    x"3F636A95",
    x"3F636D77",
    x"3F637059",
    x"3F63733C",
    x"3F63761E",
    x"3F637900",
    x"3F637BE2",
    x"3F637EC3",
    x"3F6381A5",
    x"3F638486",
    x"3F638767",
    x"3F638A49",
    x"3F638D2A",
    x"3F63900B",
    x"3F6392EB",
    x"3F6395CC",
    x"3F6398AC",
    x"3F639B8D",
    x"3F639E6D",
    x"3F63A14D",
    x"3F63A42D",
    x"3F63A70D",
    x"3F63A9EC",
    x"3F63ACCC",
    x"3F63AFAB",
    x"3F63B28A",
    x"3F63B569",
    x"3F63B848",
    x"3F63BB27",
    x"3F63BE06",
    x"3F63C0E4",
    x"3F63C3C3",
    x"3F63C6A1",
    x"3F63C97F",
    x"3F63CC5D",
    x"3F63CF3B",
    x"3F63D219",
    x"3F63D4F6",
    x"3F63D7D4",
    x"3F63DAB1",
    x"3F63DD8E",
    x"3F63E06B",
    x"3F63E348",
    x"3F63E625",
    x"3F63E901",
    x"3F63EBDE",
    x"3F63EEBA",
    x"3F63F196",
    x"3F63F473",
    x"3F63F74E",
    x"3F63FA2A",
    x"3F63FD06",
    x"3F63FFE1",
    x"3F6402BD",
    x"3F640598",
    x"3F640873",
    x"3F640B4E",
    x"3F640E29",
    x"3F641104",
    x"3F6413DE",
    x"3F6416B9",
    x"3F641993",
    x"3F641C6D",
    x"3F641F47",
    x"3F642221",
    x"3F6424FB",
    x"3F6427D4",
    x"3F642AAE",
    x"3F642D87",
    x"3F643060",
    x"3F643339",
    x"3F643612",
    x"3F6438EB",
    x"3F643BC4",
    x"3F643E9C",
    x"3F644174",
    x"3F64444D",
    x"3F644725",
    x"3F6449FD",
    x"3F644CD5",
    x"3F644FAC",
    x"3F645284",
    x"3F64555B",
    x"3F645832",
    x"3F645B0A",
    x"3F645DE1",
    x"3F6460B7",
    x"3F64638E",
    x"3F646665",
    x"3F64693B",
    x"3F646C11",
    x"3F646EE8",
    x"3F6471BE",
    x"3F647493",
    x"3F647769",
    x"3F647A3F",
    x"3F647D14",
    x"3F647FEA",
    x"3F6482BF",
    x"3F648594",
    x"3F648869",
    x"3F648B3E",
    x"3F648E12",
    x"3F6490E7",
    x"3F6493BB",
    x"3F64968F",
    x"3F649963",
    x"3F649C37",
    x"3F649F0B",
    x"3F64A1DF",
    x"3F64A4B2",
    x"3F64A786",
    x"3F64AA59",
    x"3F64AD2C",
    x"3F64AFFF",
    x"3F64B2D2",
    x"3F64B5A5",
    x"3F64B877",
    x"3F64BB4A",
    x"3F64BE1C",
    x"3F64C0EE",
    x"3F64C3C0",
    x"3F64C692",
    x"3F64C964",
    x"3F64CC35",
    x"3F64CF07",
    x"3F64D1D8",
    x"3F64D4AA",
    x"3F64D77B",
    x"3F64DA4B",
    x"3F64DD1C",
    x"3F64DFED",
    x"3F64E2BD",
    x"3F64E58E",
    x"3F64E85E",
    x"3F64EB2E",
    x"3F64EDFE",
    x"3F64F0CE",
    x"3F64F39E",
    x"3F64F66D",
    x"3F64F93D",
    x"3F64FC0C",
    x"3F64FEDB",
    x"3F6501AA",
    x"3F650479",
    x"3F650748",
    x"3F650A16",
    x"3F650CE5",
    x"3F650FB3",
    x"3F651281",
    x"3F65154F",
    x"3F65181D",
    x"3F651AEB",
    x"3F651DB8",
    x"3F652086",
    x"3F652353",
    x"3F652620",
    x"3F6528ED",
    x"3F652BBA",
    x"3F652E87",
    x"3F653154",
    x"3F653420",
    x"3F6536ED",
    x"3F6539B9",
    x"3F653C85",
    x"3F653F51",
    x"3F65421D",
    x"3F6544E8",
    x"3F6547B4",
    x"3F654A7F",
    x"3F654D4B",
    x"3F655016",
    x"3F6552E1",
    x"3F6555AC",
    x"3F655876",
    x"3F655B41",
    x"3F655E0B",
    x"3F6560D6",
    x"3F6563A0",
    x"3F65666A",
    x"3F656934",
    x"3F656BFD",
    x"3F656EC7",
    x"3F657190",
    x"3F65745A",
    x"3F657723",
    x"3F6579EC",
    x"3F657CB5",
    x"3F657F7E",
    x"3F658246",
    x"3F65850F",
    x"3F6587D7",
    x"3F658AA0",
    x"3F658D68",
    x"3F659030",
    x"3F6592F7",
    x"3F6595BF",
    x"3F659887",
    x"3F659B4E",
    x"3F659E15",
    x"3F65A0DC",
    x"3F65A3A3",
    x"3F65A66A",
    x"3F65A931",
    x"3F65ABF7",
    x"3F65AEBE",
    x"3F65B184",
    x"3F65B44A",
    x"3F65B710",
    x"3F65B9D6",
    x"3F65BC9C",
    x"3F65BF62",
    x"3F65C227",
    x"3F65C4EC",
    x"3F65C7B1",
    x"3F65CA77",
    x"3F65CD3B",
    x"3F65D000",
    x"3F65D2C5",
    x"3F65D589",
    x"3F65D84E",
    x"3F65DB12",
    x"3F65DDD6",
    x"3F65E09A",
    x"3F65E35E",
    x"3F65E621",
    x"3F65E8E5",
    x"3F65EBA8",
    x"3F65EE6C",
    x"3F65F12F",
    x"3F65F3F2",
    x"3F65F6B4",
    x"3F65F977",
    x"3F65FC3A",
    x"3F65FEFC",
    x"3F6601BE",
    x"3F660480",
    x"3F660742",
    x"3F660A04",
    x"3F660CC6",
    x"3F660F88",
    x"3F661249",
    x"3F66150A",
    x"3F6617CC",
    x"3F661A8D",
    x"3F661D4D",
    x"3F66200E",
    x"3F6622CF",
    x"3F66258F",
    x"3F662850",
    x"3F662B10",
    x"3F662DD0",
    x"3F663090",
    x"3F663350",
    x"3F66360F",
    x"3F6638CF",
    x"3F663B8E",
    x"3F663E4D",
    x"3F66410C",
    x"3F6643CB",
    x"3F66468A",
    x"3F664949",
    x"3F664C07",
    x"3F664EC6",
    x"3F665184",
    x"3F665442",
    x"3F665700",
    x"3F6659BE",
    x"3F665C7C",
    x"3F665F39",
    x"3F6661F7",
    x"3F6664B4",
    x"3F666771",
    x"3F666A2E",
    x"3F666CEB",
    x"3F666FA8",
    x"3F667264",
    x"3F667521",
    x"3F6677DD",
    x"3F667A99",
    x"3F667D55",
    x"3F668011",
    x"3F6682CD",
    x"3F668588",
    x"3F668844",
    x"3F668AFF",
    x"3F668DBA",
    x"3F669076",
    x"3F669330",
    x"3F6695EB",
    x"3F6698A6",
    x"3F669B60",
    x"3F669E1B",
    x"3F66A0D5",
    x"3F66A38F",
    x"3F66A649",
    x"3F66A903",
    x"3F66ABBC",
    x"3F66AE76",
    x"3F66B12F",
    x"3F66B3E9",
    x"3F66B6A2",
    x"3F66B95B",
    x"3F66BC14",
    x"3F66BECC",
    x"3F66C185",
    x"3F66C43D",
    x"3F66C6F6",
    x"3F66C9AE",
    x"3F66CC66",
    x"3F66CF1E",
    x"3F66D1D5",
    x"3F66D48D",
    x"3F66D744",
    x"3F66D9FC",
    x"3F66DCB3",
    x"3F66DF6A",
    x"3F66E221",
    x"3F66E4D7",
    x"3F66E78E",
    x"3F66EA45",
    x"3F66ECFB",
    x"3F66EFB1",
    x"3F66F267",
    x"3F66F51D",
    x"3F66F7D3",
    x"3F66FA88",
    x"3F66FD3E",
    x"3F66FFF3",
    x"3F6702A9",
    x"3F67055E",
    x"3F670813",
    x"3F670AC7",
    x"3F670D7C",
    x"3F671031",
    x"3F6712E5",
    x"3F671599",
    x"3F67184D",
    x"3F671B01",
    x"3F671DB5",
    x"3F672069",
    x"3F67231C",
    x"3F6725D0",
    x"3F672883",
    x"3F672B36",
    x"3F672DE9",
    x"3F67309C",
    x"3F67334F",
    x"3F673601",
    x"3F6738B4",
    x"3F673B66",
    x"3F673E18",
    x"3F6740CA",
    x"3F67437C",
    x"3F67462E",
    x"3F6748DF",
    x"3F674B91",
    x"3F674E42",
    x"3F6750F3",
    x"3F6753A5",
    x"3F675655",
    x"3F675906",
    x"3F675BB7",
    x"3F675E67",
    x"3F676118",
    x"3F6763C8",
    x"3F676678",
    x"3F676928",
    x"3F676BD8",
    x"3F676E87",
    x"3F677137",
    x"3F6773E6",
    x"3F677695",
    x"3F677944",
    x"3F677BF3",
    x"3F677EA2",
    x"3F678151",
    x"3F6783FF",
    x"3F6786AE",
    x"3F67895C",
    x"3F678C0A",
    x"3F678EB8",
    x"3F679166",
    x"3F679414",
    x"3F6796C1",
    x"3F67996F",
    x"3F679C1C",
    x"3F679EC9",
    x"3F67A176",
    x"3F67A423",
    x"3F67A6D0",
    x"3F67A97C",
    x"3F67AC29",
    x"3F67AED5",
    x"3F67B181",
    x"3F67B42D",
    x"3F67B6D9",
    x"3F67B985",
    x"3F67BC30",
    x"3F67BEDC",
    x"3F67C187",
    x"3F67C432",
    x"3F67C6DE",
    x"3F67C988",
    x"3F67CC33",
    x"3F67CEDE",
    x"3F67D188",
    x"3F67D433",
    x"3F67D6DD",
    x"3F67D987",
    x"3F67DC31",
    x"3F67DEDB",
    x"3F67E184",
    x"3F67E42E",
    x"3F67E6D7",
    x"3F67E980",
    x"3F67EC29",
    x"3F67EED2",
    x"3F67F17B",
    x"3F67F424",
    x"3F67F6CC",
    x"3F67F975",
    x"3F67FC1D",
    x"3F67FEC5",
    x"3F68016D",
    x"3F680415",
    x"3F6806BD",
    x"3F680964",
    x"3F680C0C",
    x"3F680EB3",
    x"3F68115A",
    x"3F681401",
    x"3F6816A8",
    x"3F68194F",
    x"3F681BF5",
    x"3F681E9C",
    x"3F682142",
    x"3F6823E8",
    x"3F68268E",
    x"3F682934",
    x"3F682BDA",
    x"3F682E7F",
    x"3F683125",
    x"3F6833CA",
    x"3F68366F",
    x"3F683914",
    x"3F683BB9",
    x"3F683E5E",
    x"3F684103",
    x"3F6843A7",
    x"3F68464B",
    x"3F6848F0",
    x"3F684B94",
    x"3F684E38",
    x"3F6850DB",
    x"3F68537F",
    x"3F685623",
    x"3F6858C6",
    x"3F685B69",
    x"3F685E0C",
    x"3F6860AF",
    x"3F686352",
    x"3F6865F5",
    x"3F686897",
    x"3F686B39",
    x"3F686DDC",
    x"3F68707E",
    x"3F687320",
    x"3F6875C2",
    x"3F687863",
    x"3F687B05",
    x"3F687DA6",
    x"3F688047",
    x"3F6882E9",
    x"3F68858A",
    x"3F68882A",
    x"3F688ACB",
    x"3F688D6C",
    x"3F68900C",
    x"3F6892AC",
    x"3F68954C",
    x"3F6897EC",
    x"3F689A8C",
    x"3F689D2C",
    x"3F689FCC",
    x"3F68A26B",
    x"3F68A50A",
    x"3F68A7AA",
    x"3F68AA49",
    x"3F68ACE7",
    x"3F68AF86",
    x"3F68B225",
    x"3F68B4C3",
    x"3F68B762",
    x"3F68BA00",
    x"3F68BC9E",
    x"3F68BF3C",
    x"3F68C1D9",
    x"3F68C477",
    x"3F68C714",
    x"3F68C9B2",
    x"3F68CC4F",
    x"3F68CEEC",
    x"3F68D189",
    x"3F68D426",
    x"3F68D6C2",
    x"3F68D95F",
    x"3F68DBFB",
    x"3F68DE97",
    x"3F68E134",
    x"3F68E3CF",
    x"3F68E66B",
    x"3F68E907",
    x"3F68EBA2",
    x"3F68EE3E",
    x"3F68F0D9",
    x"3F68F374",
    x"3F68F60F",
    x"3F68F8AA",
    x"3F68FB45",
    x"3F68FDDF",
    x"3F690079",
    x"3F690314",
    x"3F6905AE",
    x"3F690848",
    x"3F690AE2",
    x"3F690D7B",
    x"3F691015",
    x"3F6912AE",
    x"3F691547",
    x"3F6917E1",
    x"3F691A7A",
    x"3F691D12",
    x"3F691FAB",
    x"3F692244",
    x"3F6924DC",
    x"3F692774",
    x"3F692A0D",
    x"3F692CA5",
    x"3F692F3C",
    x"3F6931D4",
    x"3F69346C",
    x"3F693703",
    x"3F69399A",
    x"3F693C32",
    x"3F693EC9",
    x"3F694160",
    x"3F6943F6",
    x"3F69468D",
    x"3F694923",
    x"3F694BBA",
    x"3F694E50",
    x"3F6950E6",
    x"3F69537C",
    x"3F695611",
    x"3F6958A7",
    x"3F695B3D",
    x"3F695DD2",
    x"3F696067",
    x"3F6962FC",
    x"3F696591",
    x"3F696826",
    x"3F696ABA",
    x"3F696D4F",
    x"3F696FE3",
    x"3F697277",
    x"3F69750C",
    x"3F69779F",
    x"3F697A33",
    x"3F697CC7",
    x"3F697F5A",
    x"3F6981EE",
    x"3F698481",
    x"3F698714",
    x"3F6989A7",
    x"3F698C3A",
    x"3F698ECC",
    x"3F69915F",
    x"3F6993F1",
    x"3F699684",
    x"3F699916",
    x"3F699BA8",
    x"3F699E39",
    x"3F69A0CB",
    x"3F69A35D",
    x"3F69A5EE",
    x"3F69A87F",
    x"3F69AB10",
    x"3F69ADA1",
    x"3F69B032",
    x"3F69B2C3",
    x"3F69B553",
    x"3F69B7E4",
    x"3F69BA74",
    x"3F69BD04",
    x"3F69BF94",
    x"3F69C224",
    x"3F69C4B4",
    x"3F69C743",
    x"3F69C9D3",
    x"3F69CC62",
    x"3F69CEF1",
    x"3F69D180",
    x"3F69D40F",
    x"3F69D69E",
    x"3F69D92C",
    x"3F69DBBB",
    x"3F69DE49",
    x"3F69E0D7",
    x"3F69E365",
    x"3F69E5F3",
    x"3F69E881",
    x"3F69EB0E",
    x"3F69ED9C",
    x"3F69F029",
    x"3F69F2B6",
    x"3F69F543",
    x"3F69F7D0",
    x"3F69FA5D",
    x"3F69FCEA",
    x"3F69FF76",
    x"3F6A0202",
    x"3F6A048F",
    x"3F6A071B",
    x"3F6A09A7",
    x"3F6A0C32",
    x"3F6A0EBE",
    x"3F6A1149",
    x"3F6A13D5",
    x"3F6A1660",
    x"3F6A18EB",
    x"3F6A1B76",
    x"3F6A1E01",
    x"3F6A208B",
    x"3F6A2316",
    x"3F6A25A0",
    x"3F6A282A",
    x"3F6A2AB4",
    x"3F6A2D3E",
    x"3F6A2FC8",
    x"3F6A3252",
    x"3F6A34DB",
    x"3F6A3765",
    x"3F6A39EE",
    x"3F6A3C77",
    x"3F6A3F00",
    x"3F6A4189",
    x"3F6A4411",
    x"3F6A469A",
    x"3F6A4922",
    x"3F6A4BAA",
    x"3F6A4E33",
    x"3F6A50BA",
    x"3F6A5342",
    x"3F6A55CA",
    x"3F6A5851",
    x"3F6A5AD9",
    x"3F6A5D60",
    x"3F6A5FE7",
    x"3F6A626E",
    x"3F6A64F5",
    x"3F6A677C",
    x"3F6A6A02",
    x"3F6A6C89",
    x"3F6A6F0F",
    x"3F6A7195",
    x"3F6A741B",
    x"3F6A76A1",
    x"3F6A7926",
    x"3F6A7BAC",
    x"3F6A7E31",
    x"3F6A80B7",
    x"3F6A833C",
    x"3F6A85C1",
    x"3F6A8846",
    x"3F6A8ACA",
    x"3F6A8D4F",
    x"3F6A8FD3",
    x"3F6A9258",
    x"3F6A94DC",
    x"3F6A9760",
    x"3F6A99E4",
    x"3F6A9C67",
    x"3F6A9EEB",
    x"3F6AA16E",
    x"3F6AA3F2",
    x"3F6AA675",
    x"3F6AA8F8",
    x"3F6AAB7B",
    x"3F6AADFD",
    x"3F6AB080",
    x"3F6AB302",
    x"3F6AB585",
    x"3F6AB807",
    x"3F6ABA89",
    x"3F6ABD0B",
    x"3F6ABF8C",
    x"3F6AC20E",
    x"3F6AC48F",
    x"3F6AC711",
    x"3F6AC992",
    x"3F6ACC13",
    x"3F6ACE94",
    x"3F6AD115",
    x"3F6AD395",
    x"3F6AD616",
    x"3F6AD896",
    x"3F6ADB16",
    x"3F6ADD96",
    x"3F6AE016",
    x"3F6AE296",
    x"3F6AE515",
    x"3F6AE795",
    x"3F6AEA14",
    x"3F6AEC93",
    x"3F6AEF12",
    x"3F6AF191",
    x"3F6AF410",
    x"3F6AF68F",
    x"3F6AF90D",
    x"3F6AFB8C",
    x"3F6AFE0A",
    x"3F6B0088",
    x"3F6B0306",
    x"3F6B0584",
    x"3F6B0801",
    x"3F6B0A7F",
    x"3F6B0CFC",
    x"3F6B0F79",
    x"3F6B11F6",
    x"3F6B1473",
    x"3F6B16F0",
    x"3F6B196D",
    x"3F6B1BE9",
    x"3F6B1E65",
    x"3F6B20E2",
    x"3F6B235E",
    x"3F6B25DA",
    x"3F6B2855",
    x"3F6B2AD1",
    x"3F6B2D4D",
    x"3F6B2FC8",
    x"3F6B3243",
    x"3F6B34BE",
    x"3F6B3739",
    x"3F6B39B4",
    x"3F6B3C2F",
    x"3F6B3EA9",
    x"3F6B4124",
    x"3F6B439E",
    x"3F6B4618",
    x"3F6B4892",
    x"3F6B4B0C",
    x"3F6B4D85",
    x"3F6B4FFF",
    x"3F6B5278",
    x"3F6B54F1",
    x"3F6B576B",
    x"3F6B59E3",
    x"3F6B5C5C",
    x"3F6B5ED5",
    x"3F6B614D",
    x"3F6B63C6",
    x"3F6B663E",
    x"3F6B68B6",
    x"3F6B6B2E",
    x"3F6B6DA6",
    x"3F6B701E",
    x"3F6B7295",
    x"3F6B750D",
    x"3F6B7784",
    x"3F6B79FB",
    x"3F6B7C72",
    x"3F6B7EE9",
    x"3F6B815F",
    x"3F6B83D6",
    x"3F6B864C",
    x"3F6B88C3",
    x"3F6B8B39",
    x"3F6B8DAF",
    x"3F6B9025",
    x"3F6B929A",
    x"3F6B9510",
    x"3F6B9785",
    x"3F6B99FB",
    x"3F6B9C70",
    x"3F6B9EE5",
    x"3F6BA159",
    x"3F6BA3CE",
    x"3F6BA643",
    x"3F6BA8B7",
    x"3F6BAB2B",
    x"3F6BADA0",
    x"3F6BB014",
    x"3F6BB287",
    x"3F6BB4FB",
    x"3F6BB76F",
    x"3F6BB9E2",
    x"3F6BBC55",
    x"3F6BBEC8",
    x"3F6BC13B",
    x"3F6BC3AE",
    x"3F6BC621",
    x"3F6BC894",
    x"3F6BCB06",
    x"3F6BCD78",
    x"3F6BCFEA",
    x"3F6BD25C",
    x"3F6BD4CE",
    x"3F6BD740",
    x"3F6BD9B2",
    x"3F6BDC23",
    x"3F6BDE94",
    x"3F6BE105",
    x"3F6BE376",
    x"3F6BE5E7",
    x"3F6BE858",
    x"3F6BEAC9",
    x"3F6BED39",
    x"3F6BEFA9",
    x"3F6BF21A",
    x"3F6BF48A",
    x"3F6BF6F9",
    x"3F6BF969",
    x"3F6BFBD9",
    x"3F6BFE48",
    x"3F6C00B7",
    x"3F6C0327",
    x"3F6C0596",
    x"3F6C0805",
    x"3F6C0A73",
    x"3F6C0CE2",
    x"3F6C0F50",
    x"3F6C11BF",
    x"3F6C142D",
    x"3F6C169B",
    x"3F6C1909",
    x"3F6C1B76",
    x"3F6C1DE4",
    x"3F6C2051",
    x"3F6C22BF",
    x"3F6C252C",
    x"3F6C2799",
    x"3F6C2A06",
    x"3F6C2C73",
    x"3F6C2EDF",
    x"3F6C314C",
    x"3F6C33B8",
    x"3F6C3624",
    x"3F6C3890",
    x"3F6C3AFC",
    x"3F6C3D68",
    x"3F6C3FD3",
    x"3F6C423F",
    x"3F6C44AA",
    x"3F6C4715",
    x"3F6C4980",
    x"3F6C4BEB",
    x"3F6C4E56",
    x"3F6C50C1",
    x"3F6C532B",
    x"3F6C5595",
    x"3F6C5800",
    x"3F6C5A6A",
    x"3F6C5CD4",
    x"3F6C5F3D",
    x"3F6C61A7",
    x"3F6C6410",
    x"3F6C667A",
    x"3F6C68E3",
    x"3F6C6B4C",
    x"3F6C6DB5",
    x"3F6C701E",
    x"3F6C7286",
    x"3F6C74EF",
    x"3F6C7757",
    x"3F6C79BF",
    x"3F6C7C27",
    x"3F6C7E8F",
    x"3F6C80F7",
    x"3F6C835E",
    x"3F6C85C6",
    x"3F6C882D",
    x"3F6C8A94",
    x"3F6C8CFC",
    x"3F6C8F62",
    x"3F6C91C9",
    x"3F6C9430",
    x"3F6C9696",
    x"3F6C98FD",
    x"3F6C9B63",
    x"3F6C9DC9",
    x"3F6CA02F",
    x"3F6CA295",
    x"3F6CA4FA",
    x"3F6CA760",
    x"3F6CA9C5",
    x"3F6CAC2A",
    x"3F6CAE8F",
    x"3F6CB0F4",
    x"3F6CB359",
    x"3F6CB5BD",
    x"3F6CB822",
    x"3F6CBA86",
    x"3F6CBCEA",
    x"3F6CBF4F",
    x"3F6CC1B2",
    x"3F6CC416",
    x"3F6CC67A",
    x"3F6CC8DD",
    x"3F6CCB41",
    x"3F6CCDA4",
    x"3F6CD007",
    x"3F6CD26A",
    x"3F6CD4CD",
    x"3F6CD72F",
    x"3F6CD992",
    x"3F6CDBF4",
    x"3F6CDE56",
    x"3F6CE0B8",
    x"3F6CE31A",
    x"3F6CE57C",
    x"3F6CE7DE",
    x"3F6CEA3F",
    x"3F6CECA0",
    x"3F6CEF02",
    x"3F6CF163",
    x"3F6CF3C4",
    x"3F6CF624",
    x"3F6CF885",
    x"3F6CFAE5",
    x"3F6CFD46",
    x"3F6CFFA6",
    x"3F6D0206",
    x"3F6D0466",
    x"3F6D06C6",
    x"3F6D0925",
    x"3F6D0B85",
    x"3F6D0DE4",
    x"3F6D1043",
    x"3F6D12A2",
    x"3F6D1501",
    x"3F6D1760",
    x"3F6D19BF",
    x"3F6D1C1D",
    x"3F6D1E7C",
    x"3F6D20DA",
    x"3F6D2338",
    x"3F6D2596",
    x"3F6D27F4",
    x"3F6D2A51",
    x"3F6D2CAF",
    x"3F6D2F0C",
    x"3F6D3169",
    x"3F6D33C6",
    x"3F6D3623",
    x"3F6D3880",
    x"3F6D3ADD",
    x"3F6D3D39",
    x"3F6D3F95",
    x"3F6D41F2",
    x"3F6D444E",
    x"3F6D46AA",
    x"3F6D4905",
    x"3F6D4B61",
    x"3F6D4DBC",
    x"3F6D5018",
    x"3F6D5273",
    x"3F6D54CE",
    x"3F6D5729",
    x"3F6D5984",
    x"3F6D5BDE",
    x"3F6D5E39",
    x"3F6D6093",
    x"3F6D62ED",
    x"3F6D6547",
    x"3F6D67A1",
    x"3F6D69FB",
    x"3F6D6C55",
    x"3F6D6EAE",
    x"3F6D7108",
    x"3F6D7361",
    x"3F6D75BA",
    x"3F6D7813",
    x"3F6D7A6C",
    x"3F6D7CC4",
    x"3F6D7F1D",
    x"3F6D8175",
    x"3F6D83CD",
    x"3F6D8625",
    x"3F6D887D",
    x"3F6D8AD5",
    x"3F6D8D2D",
    x"3F6D8F84",
    x"3F6D91DB",
    x"3F6D9433",
    x"3F6D968A",
    x"3F6D98E1",
    x"3F6D9B37",
    x"3F6D9D8E",
    x"3F6D9FE4",
    x"3F6DA23B",
    x"3F6DA491",
    x"3F6DA6E7",
    x"3F6DA93D",
    x"3F6DAB93",
    x"3F6DADE8",
    x"3F6DB03E",
    x"3F6DB293",
    x"3F6DB4E8",
    x"3F6DB73D",
    x"3F6DB992",
    x"3F6DBBE7",
    x"3F6DBE3C",
    x"3F6DC090",
    x"3F6DC2E4",
    x"3F6DC539",
    x"3F6DC78D",
    x"3F6DC9E1",
    x"3F6DCC34",
    x"3F6DCE88",
    x"3F6DD0DB",
    x"3F6DD32F",
    x"3F6DD582",
    x"3F6DD7D5",
    x"3F6DDA28",
    x"3F6DDC7B",
    x"3F6DDECD",
    x"3F6DE120",
    x"3F6DE372",
    x"3F6DE5C4",
    x"3F6DE816",
    x"3F6DEA68",
    x"3F6DECBA",
    x"3F6DEF0B",
    x"3F6DF15D",
    x"3F6DF3AE",
    x"3F6DF5FF",
    x"3F6DF850",
    x"3F6DFAA1",
    x"3F6DFCF2",
    x"3F6DFF43",
    x"3F6E0193",
    x"3F6E03E3",
    x"3F6E0634",
    x"3F6E0884",
    x"3F6E0AD4",
    x"3F6E0D23",
    x"3F6E0F73",
    x"3F6E11C2",
    x"3F6E1412",
    x"3F6E1661",
    x"3F6E18B0",
    x"3F6E1AFF",
    x"3F6E1D4E",
    x"3F6E1F9C",
    x"3F6E21EB",
    x"3F6E2439",
    x"3F6E2687",
    x"3F6E28D5",
    x"3F6E2B23",
    x"3F6E2D71",
    x"3F6E2FBE",
    x"3F6E320C",
    x"3F6E3459",
    x"3F6E36A6",
    x"3F6E38F3",
    x"3F6E3B40",
    x"3F6E3D8D",
    x"3F6E3FD9",
    x"3F6E4226",
    x"3F6E4472",
    x"3F6E46BE",
    x"3F6E490A",
    x"3F6E4B56",
    x"3F6E4DA2",
    x"3F6E4FEE",
    x"3F6E5239",
    x"3F6E5484",
    x"3F6E56CF",
    x"3F6E591A",
    x"3F6E5B65",
    x"3F6E5DB0",
    x"3F6E5FFB",
    x"3F6E6245",
    x"3F6E648F",
    x"3F6E66D9",
    x"3F6E6924",
    x"3F6E6B6D",
    x"3F6E6DB7",
    x"3F6E7001",
    x"3F6E724A",
    x"3F6E7493",
    x"3F6E76DD",
    x"3F6E7926",
    x"3F6E7B6E",
    x"3F6E7DB7",
    x"3F6E8000",
    x"3F6E8248",
    x"3F6E8490",
    x"3F6E86D8",
    x"3F6E8920",
    x"3F6E8B68",
    x"3F6E8DB0",
    x"3F6E8FF8",
    x"3F6E923F",
    x"3F6E9486",
    x"3F6E96CD",
    x"3F6E9914",
    x"3F6E9B5B",
    x"3F6E9DA2",
    x"3F6E9FE9",
    x"3F6EA22F",
    x"3F6EA475",
    x"3F6EA6BB",
    x"3F6EA901",
    x"3F6EAB47",
    x"3F6EAD8D",
    x"3F6EAFD2",
    x"3F6EB218",
    x"3F6EB45D",
    x"3F6EB6A2",
    x"3F6EB8E7",
    x"3F6EBB2C",
    x"3F6EBD71",
    x"3F6EBFB5",
    x"3F6EC1FA",
    x"3F6EC43E",
    x"3F6EC682",
    x"3F6EC8C6",
    x"3F6ECB0A",
    x"3F6ECD4D",
    x"3F6ECF91",
    x"3F6ED1D4",
    x"3F6ED418",
    x"3F6ED65B",
    x"3F6ED89E",
    x"3F6EDAE1",
    x"3F6EDD23",
    x"3F6EDF66",
    x"3F6EE1A8",
    x"3F6EE3EA",
    x"3F6EE62C",
    x"3F6EE86E",
    x"3F6EEAB0",
    x"3F6EECF2",
    x"3F6EEF33",
    x"3F6EF175",
    x"3F6EF3B6",
    x"3F6EF5F7",
    x"3F6EF838",
    x"3F6EFA79",
    x"3F6EFCBA",
    x"3F6EFEFA",
    x"3F6F013A",
    x"3F6F037B",
    x"3F6F05BB",
    x"3F6F07FB",
    x"3F6F0A3A",
    x"3F6F0C7A",
    x"3F6F0EBA",
    x"3F6F10F9",
    x"3F6F1338",
    x"3F6F1577",
    x"3F6F17B6",
    x"3F6F19F5",
    x"3F6F1C34",
    x"3F6F1E72",
    x"3F6F20B0",
    x"3F6F22EF",
    x"3F6F252D",
    x"3F6F276B",
    x"3F6F29A8",
    x"3F6F2BE6",
    x"3F6F2E24",
    x"3F6F3061",
    x"3F6F329E",
    x"3F6F34DB",
    x"3F6F3718",
    x"3F6F3955",
    x"3F6F3B92",
    x"3F6F3DCE",
    x"3F6F400A",
    x"3F6F4247",
    x"3F6F4483",
    x"3F6F46BE",
    x"3F6F48FA",
    x"3F6F4B36",
    x"3F6F4D71",
    x"3F6F4FAD",
    x"3F6F51E8",
    x"3F6F5423",
    x"3F6F565E",
    x"3F6F5899",
    x"3F6F5AD3",
    x"3F6F5D0E",
    x"3F6F5F48",
    x"3F6F6182",
    x"3F6F63BC",
    x"3F6F65F6",
    x"3F6F6830",
    x"3F6F6A69",
    x"3F6F6CA3",
    x"3F6F6EDC",
    x"3F6F7115",
    x"3F6F734E",
    x"3F6F7587",
    x"3F6F77C0",
    x"3F6F79F8",
    x"3F6F7C31",
    x"3F6F7E69",
    x"3F6F80A1",
    x"3F6F82D9",
    x"3F6F8511",
    x"3F6F8749",
    x"3F6F8981",
    x"3F6F8BB8",
    x"3F6F8DEF",
    x"3F6F9026",
    x"3F6F925D",
    x"3F6F9494",
    x"3F6F96CB",
    x"3F6F9902",
    x"3F6F9B38",
    x"3F6F9D6E",
    x"3F6F9FA4",
    x"3F6FA1DA",
    x"3F6FA410",
    x"3F6FA646",
    x"3F6FA87C",
    x"3F6FAAB1",
    x"3F6FACE6",
    x"3F6FAF1B",
    x"3F6FB150",
    x"3F6FB385",
    x"3F6FB5BA",
    x"3F6FB7EE",
    x"3F6FBA23",
    x"3F6FBC57",
    x"3F6FBE8B",
    x"3F6FC0BF",
    x"3F6FC2F3",
    x"3F6FC527",
    x"3F6FC75A",
    x"3F6FC98E",
    x"3F6FCBC1",
    x"3F6FCDF4",
    x"3F6FD027",
    x"3F6FD25A",
    x"3F6FD48C",
    x"3F6FD6BF",
    x"3F6FD8F1",
    x"3F6FDB24",
    x"3F6FDD56",
    x"3F6FDF88",
    x"3F6FE1B9",
    x"3F6FE3EB",
    x"3F6FE61D",
    x"3F6FE84E",
    x"3F6FEA7F",
    x"3F6FECB0",
    x"3F6FEEE1",
    x"3F6FF112",
    x"3F6FF343",
    x"3F6FF573",
    x"3F6FF7A3",
    x"3F6FF9D4",
    x"3F6FFC04",
    x"3F6FFE34",
    x"3F700063",
    x"3F700293",
    x"3F7004C3",
    x"3F7006F2",
    x"3F700921",
    x"3F700B50",
    x"3F700D7F",
    x"3F700FAE",
    x"3F7011DC",
    x"3F70140B",
    x"3F701639",
    x"3F701867",
    x"3F701A95",
    x"3F701CC3",
    x"3F701EF1",
    x"3F70211F",
    x"3F70234C",
    x"3F70257A",
    x"3F7027A7",
    x"3F7029D4",
    x"3F702C01",
    x"3F702E2D",
    x"3F70305A",
    x"3F703286",
    x"3F7034B3",
    x"3F7036DF",
    x"3F70390B",
    x"3F703B37",
    x"3F703D63",
    x"3F703F8E",
    x"3F7041BA",
    x"3F7043E5",
    x"3F704610",
    x"3F70483B",
    x"3F704A66",
    x"3F704C91",
    x"3F704EBB",
    x"3F7050E6",
    x"3F705310",
    x"3F70553A",
    x"3F705764",
    x"3F70598E",
    x"3F705BB8",
    x"3F705DE1",
    x"3F70600A",
    x"3F706234",
    x"3F70645D",
    x"3F706686",
    x"3F7068AF",
    x"3F706AD7",
    x"3F706D00",
    x"3F706F28",
    x"3F707151",
    x"3F707379",
    x"3F7075A1",
    x"3F7077C8",
    x"3F7079F0",
    x"3F707C18",
    x"3F707E3F",
    x"3F708066",
    x"3F70828D",
    x"3F7084B4",
    x"3F7086DB",
    x"3F708902",
    x"3F708B28",
    x"3F708D4F",
    x"3F708F75",
    x"3F70919B",
    x"3F7093C1",
    x"3F7095E7",
    x"3F70980C",
    x"3F709A32",
    x"3F709C57",
    x"3F709E7C",
    x"3F70A0A2",
    x"3F70A2C6",
    x"3F70A4EB",
    x"3F70A710",
    x"3F70A934",
    x"3F70AB59",
    x"3F70AD7D",
    x"3F70AFA1",
    x"3F70B1C5",
    x"3F70B3E9",
    x"3F70B60C",
    x"3F70B830",
    x"3F70BA53",
    x"3F70BC76",
    x"3F70BE99",
    x"3F70C0BC",
    x"3F70C2DF",
    x"3F70C501",
    x"3F70C724",
    x"3F70C946",
    x"3F70CB68",
    x"3F70CD8A",
    x"3F70CFAC",
    x"3F70D1CE",
    x"3F70D3F0",
    x"3F70D611",
    x"3F70D832",
    x"3F70DA54",
    x"3F70DC75",
    x"3F70DE95",
    x"3F70E0B6",
    x"3F70E2D7",
    x"3F70E4F7",
    x"3F70E717",
    x"3F70E938",
    x"3F70EB58",
    x"3F70ED77",
    x"3F70EF97",
    x"3F70F1B7",
    x"3F70F3D6",
    x"3F70F5F5",
    x"3F70F814",
    x"3F70FA33",
    x"3F70FC52",
    x"3F70FE71",
    x"3F71008F",
    x"3F7102AE",
    x"3F7104CC",
    x"3F7106EA",
    x"3F710908",
    x"3F710B26",
    x"3F710D44",
    x"3F710F61",
    x"3F71117F",
    x"3F71139C",
    x"3F7115B9",
    x"3F7117D6",
    x"3F7119F3",
    x"3F711C0F",
    x"3F711E2C",
    x"3F712048",
    x"3F712264",
    x"3F712480",
    x"3F71269C",
    x"3F7128B8",
    x"3F712AD4",
    x"3F712CEF",
    x"3F712F0B",
    x"3F713126",
    x"3F713341",
    x"3F71355C",
    x"3F713776",
    x"3F713991",
    x"3F713BAC",
    x"3F713DC6",
    x"3F713FE0",
    x"3F7141FA",
    x"3F714414",
    x"3F71462E",
    x"3F714847",
    x"3F714A61",
    x"3F714C7A",
    x"3F714E93",
    x"3F7150AC",
    x"3F7152C5",
    x"3F7154DE",
    x"3F7156F6",
    x"3F71590F",
    x"3F715B27",
    x"3F715D3F",
    x"3F715F57",
    x"3F71616F",
    x"3F716387",
    x"3F71659F",
    x"3F7167B6",
    x"3F7169CD",
    x"3F716BE4",
    x"3F716DFB",
    x"3F717012",
    x"3F717229",
    x"3F71743F",
    x"3F717656",
    x"3F71786C",
    x"3F717A82",
    x"3F717C98",
    x"3F717EAE",
    x"3F7180C4",
    x"3F7182D9",
    x"3F7184EF",
    x"3F718704",
    x"3F718919",
    x"3F718B2E",
    x"3F718D43",
    x"3F718F57",
    x"3F71916C",
    x"3F719380",
    x"3F719594",
    x"3F7197A8",
    x"3F7199BC",
    x"3F719BD0",
    x"3F719DE4",
    x"3F719FF7",
    x"3F71A20B",
    x"3F71A41E",
    x"3F71A631",
    x"3F71A844",
    x"3F71AA57",
    x"3F71AC69",
    x"3F71AE7C",
    x"3F71B08E",
    x"3F71B2A0",
    x"3F71B4B2",
    x"3F71B6C4",
    x"3F71B8D6",
    x"3F71BAE7",
    x"3F71BCF9",
    x"3F71BF0A",
    x"3F71C11B",
    x"3F71C32C",
    x"3F71C53D",
    x"3F71C74E",
    x"3F71C95F",
    x"3F71CB6F",
    x"3F71CD7F",
    x"3F71CF8F",
    x"3F71D19F",
    x"3F71D3AF",
    x"3F71D5BF",
    x"3F71D7CF",
    x"3F71D9DE",
    x"3F71DBED",
    x"3F71DDFC",
    x"3F71E00B",
    x"3F71E21A",
    x"3F71E429",
    x"3F71E637",
    x"3F71E846",
    x"3F71EA54",
    x"3F71EC62",
    x"3F71EE70",
    x"3F71F07E",
    x"3F71F28C",
    x"3F71F499",
    x"3F71F6A6",
    x"3F71F8B4",
    x"3F71FAC1",
    x"3F71FCCE",
    x"3F71FEDA",
    x"3F7200E7",
    x"3F7202F4",
    x"3F720500",
    x"3F72070C",
    x"3F720918",
    x"3F720B24",
    x"3F720D30",
    x"3F720F3C",
    x"3F721147",
    x"3F721352",
    x"3F72155E",
    x"3F721769",
    x"3F721973",
    x"3F721B7E",
    x"3F721D89",
    x"3F721F93",
    x"3F72219E",
    x"3F7223A8",
    x"3F7225B2",
    x"3F7227BC",
    x"3F7229C5",
    x"3F722BCF",
    x"3F722DD8",
    x"3F722FE2",
    x"3F7231EB",
    x"3F7233F4",
    x"3F7235FD",
    x"3F723805",
    x"3F723A0E",
    x"3F723C16",
    x"3F723E1F",
    x"3F724027",
    x"3F72422F",
    x"3F724437",
    x"3F72463E",
    x"3F724846",
    x"3F724A4D",
    x"3F724C54",
    x"3F724E5C",
    x"3F725063",
    x"3F725269",
    x"3F725470",
    x"3F725677",
    x"3F72587D",
    x"3F725A83",
    x"3F725C89",
    x"3F725E8F",
    x"3F726095",
    x"3F72629B",
    x"3F7264A0",
    x"3F7266A5",
    x"3F7268AB",
    x"3F726AB0",
    x"3F726CB5",
    x"3F726EB9",
    x"3F7270BE",
    x"3F7272C2",
    x"3F7274C7",
    x"3F7276CB",
    x"3F7278CF",
    x"3F727AD3",
    x"3F727CD7",
    x"3F727EDA",
    x"3F7280DE",
    x"3F7282E1",
    x"3F7284E4",
    x"3F7286E7",
    x"3F7288EA",
    x"3F728AED",
    x"3F728CEF",
    x"3F728EF2",
    x"3F7290F4",
    x"3F7292F6",
    x"3F7294F8",
    x"3F7296FA",
    x"3F7298FC",
    x"3F729AFD",
    x"3F729CFF",
    x"3F729F00",
    x"3F72A101",
    x"3F72A302",
    x"3F72A503",
    x"3F72A703",
    x"3F72A904",
    x"3F72AB04",
    x"3F72AD05",
    x"3F72AF05",
    x"3F72B105",
    x"3F72B304",
    x"3F72B504",
    x"3F72B704",
    x"3F72B903",
    x"3F72BB02",
    x"3F72BD01",
    x"3F72BF00",
    x"3F72C0FF",
    x"3F72C2FE",
    x"3F72C4FC",
    x"3F72C6FA",
    x"3F72C8F9",
    x"3F72CAF7",
    x"3F72CCF5",
    x"3F72CEF2",
    x"3F72D0F0",
    x"3F72D2ED",
    x"3F72D4EB",
    x"3F72D6E8",
    x"3F72D8E5",
    x"3F72DAE2",
    x"3F72DCDE",
    x"3F72DEDB",
    x"3F72E0D7",
    x"3F72E2D4",
    x"3F72E4D0",
    x"3F72E6CC",
    x"3F72E8C8",
    x"3F72EAC3",
    x"3F72ECBF",
    x"3F72EEBA",
    x"3F72F0B6",
    x"3F72F2B1",
    x"3F72F4AC",
    x"3F72F6A7",
    x"3F72F8A1",
    x"3F72FA9C",
    x"3F72FC96",
    x"3F72FE90",
    x"3F73008B",
    x"3F730284",
    x"3F73047E",
    x"3F730678",
    x"3F730871",
    x"3F730A6B",
    x"3F730C64",
    x"3F730E5D",
    x"3F731056",
    x"3F73124F",
    x"3F731447",
    x"3F731640",
    x"3F731838",
    x"3F731A30",
    x"3F731C28",
    x"3F731E20",
    x"3F732018",
    x"3F732210",
    x"3F732407",
    x"3F7325FE",
    x"3F7327F6",
    x"3F7329ED",
    x"3F732BE4",
    x"3F732DDA",
    x"3F732FD1",
    x"3F7331C7",
    x"3F7333BE",
    x"3F7335B4",
    x"3F7337AA",
    x"3F7339A0",
    x"3F733B95",
    x"3F733D8B",
    x"3F733F80",
    x"3F734175",
    x"3F73436B",
    x"3F734560",
    x"3F734754",
    x"3F734949",
    x"3F734B3E",
    x"3F734D32",
    x"3F734F26",
    x"3F73511A",
    x"3F73530E",
    x"3F735502",
    x"3F7356F6",
    x"3F7358E9",
    x"3F735ADC",
    x"3F735CD0",
    x"3F735EC3",
    x"3F7360B6",
    x"3F7362A8",
    x"3F73649B",
    x"3F73668E",
    x"3F736880",
    x"3F736A72",
    x"3F736C64",
    x"3F736E56",
    x"3F737048",
    x"3F737239",
    x"3F73742B",
    x"3F73761C",
    x"3F73780D",
    x"3F7379FE",
    x"3F737BEF",
    x"3F737DE0",
    x"3F737FD0",
    x"3F7381C1",
    x"3F7383B1",
    x"3F7385A1",
    x"3F738791",
    x"3F738981",
    x"3F738B71",
    x"3F738D60",
    x"3F738F50",
    x"3F73913F",
    x"3F73932E",
    x"3F73951D",
    x"3F73970C",
    x"3F7398FA",
    x"3F739AE9",
    x"3F739CD7",
    x"3F739EC5",
    x"3F73A0B4",
    x"3F73A2A1",
    x"3F73A48F",
    x"3F73A67D",
    x"3F73A86A",
    x"3F73AA58",
    x"3F73AC45",
    x"3F73AE32",
    x"3F73B01F",
    x"3F73B20C",
    x"3F73B3F8",
    x"3F73B5E5",
    x"3F73B7D1",
    x"3F73B9BD",
    x"3F73BBA9",
    x"3F73BD95",
    x"3F73BF81",
    x"3F73C16C",
    x"3F73C358",
    x"3F73C543",
    x"3F73C72E",
    x"3F73C919",
    x"3F73CB04",
    x"3F73CCEF",
    x"3F73CED9",
    x"3F73D0C4",
    x"3F73D2AE",
    x"3F73D498",
    x"3F73D682",
    x"3F73D86C",
    x"3F73DA56",
    x"3F73DC3F",
    x"3F73DE28",
    x"3F73E012",
    x"3F73E1FB",
    x"3F73E3E4",
    x"3F73E5CC",
    x"3F73E7B5",
    x"3F73E99E",
    x"3F73EB86",
    x"3F73ED6E",
    x"3F73EF56",
    x"3F73F13E",
    x"3F73F326",
    x"3F73F50D",
    x"3F73F6F5",
    x"3F73F8DC",
    x"3F73FAC3",
    x"3F73FCAA",
    x"3F73FE91",
    x"3F740078",
    x"3F74025F",
    x"3F740445",
    x"3F74062B",
    x"3F740812",
    x"3F7409F8",
    x"3F740BDD",
    x"3F740DC3",
    x"3F740FA9",
    x"3F74118E",
    x"3F741373",
    x"3F741558",
    x"3F74173D",
    x"3F741922",
    x"3F741B07",
    x"3F741CEB",
    x"3F741ED0",
    x"3F7420B4",
    x"3F742298",
    x"3F74247C",
    x"3F742660",
    x"3F742843",
    x"3F742A27",
    x"3F742C0A",
    x"3F742DED",
    x"3F742FD1",
    x"3F7431B3",
    x"3F743396",
    x"3F743579",
    x"3F74375B",
    x"3F74393E",
    x"3F743B20",
    x"3F743D02",
    x"3F743EE4",
    x"3F7440C5",
    x"3F7442A7",
    x"3F744488",
    x"3F74466A",
    x"3F74484B",
    x"3F744A2C",
    x"3F744C0D",
    x"3F744DED",
    x"3F744FCE",
    x"3F7451AE",
    x"3F74538F",
    x"3F74556F",
    x"3F74574F",
    x"3F74592F",
    x"3F745B0E",
    x"3F745CEE",
    x"3F745ECD",
    x"3F7460AC",
    x"3F74628B",
    x"3F74646A",
    x"3F746649",
    x"3F746828",
    x"3F746A06",
    x"3F746BE5",
    x"3F746DC3",
    x"3F746FA1",
    x"3F74717F",
    x"3F74735D",
    x"3F74753A",
    x"3F747718",
    x"3F7478F5",
    x"3F747AD2",
    x"3F747CAF",
    x"3F747E8C",
    x"3F748069",
    x"3F748245",
    x"3F748422",
    x"3F7485FE",
    x"3F7487DA",
    x"3F7489B6",
    x"3F748B92",
    x"3F748D6E",
    x"3F748F49",
    x"3F749125",
    x"3F749300",
    x"3F7494DB",
    x"3F7496B6",
    x"3F749891",
    x"3F749A6B",
    x"3F749C46",
    x"3F749E20",
    x"3F749FFA",
    x"3F74A1D5",
    x"3F74A3AE",
    x"3F74A588",
    x"3F74A762",
    x"3F74A93B",
    x"3F74AB15",
    x"3F74ACEE",
    x"3F74AEC7",
    x"3F74B0A0",
    x"3F74B279",
    x"3F74B451",
    x"3F74B62A",
    x"3F74B802",
    x"3F74B9DA",
    x"3F74BBB2",
    x"3F74BD8A",
    x"3F74BF62",
    x"3F74C139",
    x"3F74C311",
    x"3F74C4E8",
    x"3F74C6BF",
    x"3F74C896",
    x"3F74CA6D",
    x"3F74CC44",
    x"3F74CE1A",
    x"3F74CFF0",
    x"3F74D1C7",
    x"3F74D39D",
    x"3F74D573",
    x"3F74D749",
    x"3F74D91E",
    x"3F74DAF4",
    x"3F74DCC9",
    x"3F74DE9E",
    x"3F74E073",
    x"3F74E248",
    x"3F74E41D",
    x"3F74E5F2",
    x"3F74E7C6",
    x"3F74E99A",
    x"3F74EB6F",
    x"3F74ED43",
    x"3F74EF17",
    x"3F74F0EA",
    x"3F74F2BE",
    x"3F74F491",
    x"3F74F665",
    x"3F74F838",
    x"3F74FA0B",
    x"3F74FBDE",
    x"3F74FDB0",
    x"3F74FF83",
    x"3F750155",
    x"3F750327",
    x"3F7504FA",
    x"3F7506CC",
    x"3F75089D",
    x"3F750A6F",
    x"3F750C41",
    x"3F750E12",
    x"3F750FE3",
    x"3F7511B4",
    x"3F751385",
    x"3F751556",
    x"3F751727",
    x"3F7518F7",
    x"3F751AC7",
    x"3F751C98",
    x"3F751E68",
    x"3F752038",
    x"3F752207",
    x"3F7523D7",
    x"3F7525A6",
    x"3F752776",
    x"3F752945",
    x"3F752B14",
    x"3F752CE3",
    x"3F752EB1",
    x"3F753080",
    x"3F75324E",
    x"3F75341D",
    x"3F7535EB",
    x"3F7537B9",
    x"3F753987",
    x"3F753B54",
    x"3F753D22",
    x"3F753EEF",
    x"3F7540BC",
    x"3F754289",
    x"3F754456",
    x"3F754623",
    x"3F7547F0",
    x"3F7549BC",
    x"3F754B89",
    x"3F754D55",
    x"3F754F21",
    x"3F7550ED",
    x"3F7552B9",
    x"3F755484",
    x"3F755650",
    x"3F75581B",
    x"3F7559E6",
    x"3F755BB1",
    x"3F755D7C",
    x"3F755F47",
    x"3F756111",
    x"3F7562DC",
    x"3F7564A6",
    x"3F756670",
    x"3F75683A",
    x"3F756A04",
    x"3F756BCE",
    x"3F756D97",
    x"3F756F61",
    x"3F75712A",
    x"3F7572F3",
    x"3F7574BC",
    x"3F757685",
    x"3F75784D",
    x"3F757A16",
    x"3F757BDE",
    x"3F757DA7",
    x"3F757F6F",
    x"3F758136",
    x"3F7582FE",
    x"3F7584C6",
    x"3F75868D",
    x"3F758855",
    x"3F758A1C",
    x"3F758BE3",
    x"3F758DAA",
    x"3F758F70",
    x"3F759137",
    x"3F7592FE",
    x"3F7594C4",
    x"3F75968A",
    x"3F759850",
    x"3F759A16",
    x"3F759BDB",
    x"3F759DA1",
    x"3F759F66",
    x"3F75A12C",
    x"3F75A2F1",
    x"3F75A4B6",
    x"3F75A67B",
    x"3F75A83F",
    x"3F75AA04",
    x"3F75ABC8",
    x"3F75AD8C",
    x"3F75AF50",
    x"3F75B114",
    x"3F75B2D8",
    x"3F75B49C",
    x"3F75B65F",
    x"3F75B822",
    x"3F75B9E6",
    x"3F75BBA9",
    x"3F75BD6C",
    x"3F75BF2E",
    x"3F75C0F1",
    x"3F75C2B3",
    x"3F75C476",
    x"3F75C638",
    x"3F75C7FA",
    x"3F75C9BC",
    x"3F75CB7D",
    x"3F75CD3F",
    x"3F75CF00",
    x"3F75D0C2",
    x"3F75D283",
    x"3F75D444",
    x"3F75D604",
    x"3F75D7C5",
    x"3F75D986",
    x"3F75DB46",
    x"3F75DD06",
    x"3F75DEC6",
    x"3F75E086",
    x"3F75E246",
    x"3F75E406",
    x"3F75E5C5",
    x"3F75E784",
    x"3F75E944",
    x"3F75EB03",
    x"3F75ECC2",
    x"3F75EE80",
    x"3F75F03F",
    x"3F75F1FD",
    x"3F75F3BC",
    x"3F75F57A",
    x"3F75F738",
    x"3F75F8F6",
    x"3F75FAB3",
    x"3F75FC71",
    x"3F75FE2E",
    x"3F75FFEB",
    x"3F7601A9",
    x"3F760366",
    x"3F760522",
    x"3F7606DF",
    x"3F76089C",
    x"3F760A58",
    x"3F760C14",
    x"3F760DD0",
    x"3F760F8C",
    x"3F761148",
    x"3F761304",
    x"3F7614BF",
    x"3F76167A",
    x"3F761836",
    x"3F7619F1",
    x"3F761BAB",
    x"3F761D66",
    x"3F761F21",
    x"3F7620DB",
    x"3F762296",
    x"3F762450",
    x"3F76260A",
    x"3F7627C3",
    x"3F76297D",
    x"3F762B37",
    x"3F762CF0",
    x"3F762EA9",
    x"3F763063",
    x"3F76321B",
    x"3F7633D4",
    x"3F76358D",
    x"3F763745",
    x"3F7638FE",
    x"3F763AB6",
    x"3F763C6E",
    x"3F763E26",
    x"3F763FDE",
    x"3F764195",
    x"3F76434D",
    x"3F764504",
    x"3F7646BB",
    x"3F764872",
    x"3F764A29",
    x"3F764BE0",
    x"3F764D97",
    x"3F764F4D",
    x"3F765103",
    x"3F7652B9",
    x"3F76546F",
    x"3F765625",
    x"3F7657DB",
    x"3F765991",
    x"3F765B46",
    x"3F765CFB",
    x"3F765EB0",
    x"3F766065",
    x"3F76621A",
    x"3F7663CF",
    x"3F766583",
    x"3F766738",
    x"3F7668EC",
    x"3F766AA0",
    x"3F766C54",
    x"3F766E08",
    x"3F766FBB",
    x"3F76716F",
    x"3F767322",
    x"3F7674D5",
    x"3F767688",
    x"3F76783B",
    x"3F7679EE",
    x"3F767BA0",
    x"3F767D53",
    x"3F767F05",
    x"3F7680B7",
    x"3F768269",
    x"3F76841B",
    x"3F7685CD",
    x"3F76877E",
    x"3F768930",
    x"3F768AE1",
    x"3F768C92",
    x"3F768E43",
    x"3F768FF4",
    x"3F7691A4",
    x"3F769355",
    x"3F769505",
    x"3F7696B5",
    x"3F769865",
    x"3F769A15",
    x"3F769BC5",
    x"3F769D75",
    x"3F769F24",
    x"3F76A0D3",
    x"3F76A283",
    x"3F76A432",
    x"3F76A5E0",
    x"3F76A78F",
    x"3F76A93E",
    x"3F76AAEC",
    x"3F76AC9A",
    x"3F76AE49",
    x"3F76AFF7",
    x"3F76B1A4",
    x"3F76B352",
    x"3F76B500",
    x"3F76B6AD",
    x"3F76B85A",
    x"3F76BA07",
    x"3F76BBB4",
    x"3F76BD61",
    x"3F76BF0E",
    x"3F76C0BA",
    x"3F76C266",
    x"3F76C413",
    x"3F76C5BF",
    x"3F76C76B",
    x"3F76C916",
    x"3F76CAC2",
    x"3F76CC6D",
    x"3F76CE19",
    x"3F76CFC4",
    x"3F76D16F",
    x"3F76D31A",
    x"3F76D4C4",
    x"3F76D66F",
    x"3F76D819",
    x"3F76D9C4",
    x"3F76DB6E",
    x"3F76DD18",
    x"3F76DEC1",
    x"3F76E06B",
    x"3F76E215",
    x"3F76E3BE",
    x"3F76E567",
    x"3F76E710",
    x"3F76E8B9",
    x"3F76EA62",
    x"3F76EC0B",
    x"3F76EDB3",
    x"3F76EF5B",
    x"3F76F103",
    x"3F76F2AC",
    x"3F76F453",
    x"3F76F5FB",
    x"3F76F7A3",
    x"3F76F94A",
    x"3F76FAF1",
    x"3F76FC99",
    x"3F76FE40",
    x"3F76FFE6",
    x"3F77018D",
    x"3F770334",
    x"3F7704DA",
    x"3F770680",
    x"3F770826",
    x"3F7709CC",
    x"3F770B72",
    x"3F770D18",
    x"3F770EBD",
    x"3F771063",
    x"3F771208",
    x"3F7713AD",
    x"3F771552",
    x"3F7716F6",
    x"3F77189B",
    x"3F771A3F",
    x"3F771BE4",
    x"3F771D88",
    x"3F771F2C",
    x"3F7720D0",
    x"3F772274",
    x"3F772417",
    x"3F7725BA",
    x"3F77275E",
    x"3F772901",
    x"3F772AA4",
    x"3F772C47",
    x"3F772DE9",
    x"3F772F8C",
    x"3F77312E",
    x"3F7732D0",
    x"3F773472",
    x"3F773614",
    x"3F7737B6",
    x"3F773958",
    x"3F773AF9",
    x"3F773C9B",
    x"3F773E3C",
    x"3F773FDD",
    x"3F77417E",
    x"3F77431E",
    x"3F7744BF",
    x"3F77465F",
    x"3F774800",
    x"3F7749A0",
    x"3F774B40",
    x"3F774CE0",
    x"3F774E7F",
    x"3F77501F",
    x"3F7751BE",
    x"3F77535E",
    x"3F7754FD",
    x"3F77569C",
    x"3F77583A",
    x"3F7759D9",
    x"3F775B78",
    x"3F775D16",
    x"3F775EB4",
    x"3F776052",
    x"3F7761F0",
    x"3F77638E",
    x"3F77652B",
    x"3F7766C9",
    x"3F776866",
    x"3F776A03",
    x"3F776BA0",
    x"3F776D3D",
    x"3F776EDA",
    x"3F777076",
    x"3F777213",
    x"3F7773AF",
    x"3F77754B",
    x"3F7776E7",
    x"3F777883",
    x"3F777A1F",
    x"3F777BBA",
    x"3F777D56",
    x"3F777EF1",
    x"3F77808C",
    x"3F778227",
    x"3F7783C2",
    x"3F77855C",
    x"3F7786F7",
    x"3F778891",
    x"3F778A2B",
    x"3F778BC5",
    x"3F778D5F",
    x"3F778EF9",
    x"3F779092",
    x"3F77922C",
    x"3F7793C5",
    x"3F77955E",
    x"3F7796F7",
    x"3F779890",
    x"3F779A29",
    x"3F779BC1",
    x"3F779D5A",
    x"3F779EF2",
    x"3F77A08A",
    x"3F77A222",
    x"3F77A3BA",
    x"3F77A551",
    x"3F77A6E9",
    x"3F77A880",
    x"3F77AA17",
    x"3F77ABAE",
    x"3F77AD45",
    x"3F77AEDC",
    x"3F77B073",
    x"3F77B209",
    x"3F77B39F",
    x"3F77B535",
    x"3F77B6CB",
    x"3F77B861",
    x"3F77B9F7",
    x"3F77BB8D",
    x"3F77BD22",
    x"3F77BEB7",
    x"3F77C04C",
    x"3F77C1E1",
    x"3F77C376",
    x"3F77C50B",
    x"3F77C69F",
    x"3F77C834",
    x"3F77C9C8",
    x"3F77CB5C",
    x"3F77CCF0",
    x"3F77CE83",
    x"3F77D017",
    x"3F77D1AB",
    x"3F77D33E",
    x"3F77D4D1",
    x"3F77D664",
    x"3F77D7F7",
    x"3F77D98A",
    x"3F77DB1C",
    x"3F77DCAF",
    x"3F77DE41",
    x"3F77DFD3",
    x"3F77E165",
    x"3F77E2F7",
    x"3F77E488",
    x"3F77E61A",
    x"3F77E7AB",
    x"3F77E93D",
    x"3F77EACE",
    x"3F77EC5F",
    x"3F77EDEF",
    x"3F77EF80",
    x"3F77F110",
    x"3F77F2A1",
    x"3F77F431",
    x"3F77F5C1",
    x"3F77F751",
    x"3F77F8E1",
    x"3F77FA70",
    x"3F77FC00",
    x"3F77FD8F",
    x"3F77FF1E",
    x"3F7800AD",
    x"3F78023C",
    x"3F7803CA",
    x"3F780559",
    x"3F7806E7",
    x"3F780876",
    x"3F780A04",
    x"3F780B92",
    x"3F780D1F",
    x"3F780EAD",
    x"3F78103A",
    x"3F7811C8",
    x"3F781355",
    x"3F7814E2",
    x"3F78166F",
    x"3F7817FC",
    x"3F781988",
    x"3F781B15",
    x"3F781CA1",
    x"3F781E2D",
    x"3F781FB9",
    x"3F782145",
    x"3F7822D1",
    x"3F78245C",
    x"3F7825E8",
    x"3F782773",
    x"3F7828FE",
    x"3F782A89",
    x"3F782C14",
    x"3F782D9E",
    x"3F782F29",
    x"3F7830B3",
    x"3F78323D",
    x"3F7833C7",
    x"3F783551",
    x"3F7836DB",
    x"3F783865",
    x"3F7839EE",
    x"3F783B77",
    x"3F783D01",
    x"3F783E8A",
    x"3F784012",
    x"3F78419B",
    x"3F784324",
    x"3F7844AC",
    x"3F784634",
    x"3F7847BC",
    x"3F784944",
    x"3F784ACC",
    x"3F784C54",
    x"3F784DDB",
    x"3F784F63",
    x"3F7850EA",
    x"3F785271",
    x"3F7853F8",
    x"3F78557F",
    x"3F785705",
    x"3F78588C",
    x"3F785A12",
    x"3F785B98",
    x"3F785D1E",
    x"3F785EA4",
    x"3F78602A",
    x"3F7861AF",
    x"3F786335",
    x"3F7864BA",
    x"3F78663F",
    x"3F7867C4",
    x"3F786949",
    x"3F786ACE",
    x"3F786C52",
    x"3F786DD6",
    x"3F786F5B",
    x"3F7870DF",
    x"3F787263",
    x"3F7873E6",
    x"3F78756A",
    x"3F7876ED",
    x"3F787871",
    x"3F7879F4",
    x"3F787B77",
    x"3F787CFA",
    x"3F787E7D",
    x"3F787FFF",
    x"3F788182",
    x"3F788304",
    x"3F788486",
    x"3F788608",
    x"3F78878A",
    x"3F78890B",
    x"3F788A8D",
    x"3F788C0E",
    x"3F788D8F",
    x"3F788F11",
    x"3F789091",
    x"3F789212",
    x"3F789393",
    x"3F789513",
    x"3F789694",
    x"3F789814",
    x"3F789994",
    x"3F789B14",
    x"3F789C93",
    x"3F789E13",
    x"3F789F92",
    x"3F78A112",
    x"3F78A291",
    x"3F78A410",
    x"3F78A58F",
    x"3F78A70D",
    x"3F78A88C",
    x"3F78AA0A",
    x"3F78AB88",
    x"3F78AD06",
    x"3F78AE84",
    x"3F78B002",
    x"3F78B180",
    x"3F78B2FD",
    x"3F78B47B",
    x"3F78B5F8",
    x"3F78B775",
    x"3F78B8F2",
    x"3F78BA6E",
    x"3F78BBEB",
    x"3F78BD67",
    x"3F78BEE4",
    x"3F78C060",
    x"3F78C1DC",
    x"3F78C358",
    x"3F78C4D3",
    x"3F78C64F",
    x"3F78C7CA",
    x"3F78C945",
    x"3F78CAC1",
    x"3F78CC3B",
    x"3F78CDB6",
    x"3F78CF31",
    x"3F78D0AB",
    x"3F78D226",
    x"3F78D3A0",
    x"3F78D51A",
    x"3F78D694",
    x"3F78D80E",
    x"3F78D987",
    x"3F78DB01",
    x"3F78DC7A",
    x"3F78DDF3",
    x"3F78DF6C",
    x"3F78E0E5",
    x"3F78E25D",
    x"3F78E3D6",
    x"3F78E54E",
    x"3F78E6C7",
    x"3F78E83F",
    x"3F78E9B7",
    x"3F78EB2E",
    x"3F78ECA6",
    x"3F78EE1D",
    x"3F78EF95",
    x"3F78F10C",
    x"3F78F283",
    x"3F78F3FA",
    x"3F78F571",
    x"3F78F6E7",
    x"3F78F85E",
    x"3F78F9D4",
    x"3F78FB4A",
    x"3F78FCC0",
    x"3F78FE36",
    x"3F78FFAC",
    x"3F790121",
    x"3F790296",
    x"3F79040C",
    x"3F790581",
    x"3F7906F6",
    x"3F79086A",
    x"3F7909DF",
    x"3F790B54",
    x"3F790CC8",
    x"3F790E3C",
    x"3F790FB0",
    x"3F791124",
    x"3F791298",
    x"3F79140B",
    x"3F79157F",
    x"3F7916F2",
    x"3F791865",
    x"3F7919D8",
    x"3F791B4B",
    x"3F791CBE",
    x"3F791E30",
    x"3F791FA3",
    x"3F792115",
    x"3F792287",
    x"3F7923F9",
    x"3F79256B",
    x"3F7926DC",
    x"3F79284E",
    x"3F7929BF",
    x"3F792B30",
    x"3F792CA1",
    x"3F792E12",
    x"3F792F83",
    x"3F7930F3",
    x"3F793264",
    x"3F7933D4",
    x"3F793544",
    x"3F7936B4",
    x"3F793824",
    x"3F793994",
    x"3F793B03",
    x"3F793C73",
    x"3F793DE2",
    x"3F793F51",
    x"3F7940C0",
    x"3F79422F",
    x"3F79439D",
    x"3F79450C",
    x"3F79467A",
    x"3F7947E8",
    x"3F794956",
    x"3F794AC4",
    x"3F794C32",
    x"3F794D9F",
    x"3F794F0D",
    x"3F79507A",
    x"3F7951E7",
    x"3F795354",
    x"3F7954C1",
    x"3F79562E",
    x"3F79579A",
    x"3F795907",
    x"3F795A73",
    x"3F795BDF",
    x"3F795D4B",
    x"3F795EB7",
    x"3F796022",
    x"3F79618E",
    x"3F7962F9",
    x"3F796464",
    x"3F7965CF",
    x"3F79673A",
    x"3F7968A5",
    x"3F796A0F",
    x"3F796B7A",
    x"3F796CE4",
    x"3F796E4E",
    x"3F796FB8",
    x"3F797122",
    x"3F79728C",
    x"3F7973F5",
    x"3F79755F",
    x"3F7976C8",
    x"3F797831",
    x"3F79799A",
    x"3F797B03",
    x"3F797C6B",
    x"3F797DD4",
    x"3F797F3C",
    x"3F7980A4",
    x"3F79820C",
    x"3F798374",
    x"3F7984DC",
    x"3F798643",
    x"3F7987AB",
    x"3F798912",
    x"3F798A79",
    x"3F798BE0",
    x"3F798D47",
    x"3F798EAE",
    x"3F799014",
    x"3F79917A",
    x"3F7992E1",
    x"3F799447",
    x"3F7995AD",
    x"3F799712",
    x"3F799878",
    x"3F7999DE",
    x"3F799B43",
    x"3F799CA8",
    x"3F799E0D",
    x"3F799F72",
    x"3F79A0D7",
    x"3F79A23B",
    x"3F79A3A0",
    x"3F79A504",
    x"3F79A668",
    x"3F79A7CC",
    x"3F79A930",
    x"3F79AA93",
    x"3F79ABF7",
    x"3F79AD5A",
    x"3F79AEBD",
    x"3F79B020",
    x"3F79B183",
    x"3F79B2E6",
    x"3F79B449",
    x"3F79B5AB",
    x"3F79B70D",
    x"3F79B870",
    x"3F79B9D2",
    x"3F79BB33",
    x"3F79BC95",
    x"3F79BDF7",
    x"3F79BF58",
    x"3F79C0B9",
    x"3F79C21A",
    x"3F79C37B",
    x"3F79C4DC",
    x"3F79C63D",
    x"3F79C79D",
    x"3F79C8FE",
    x"3F79CA5E",
    x"3F79CBBE",
    x"3F79CD1E",
    x"3F79CE7E",
    x"3F79CFDD",
    x"3F79D13D",
    x"3F79D29C",
    x"3F79D3FB",
    x"3F79D55A",
    x"3F79D6B9",
    x"3F79D818",
    x"3F79D976",
    x"3F79DAD5",
    x"3F79DC33",
    x"3F79DD91",
    x"3F79DEEF",
    x"3F79E04D",
    x"3F79E1AA",
    x"3F79E308",
    x"3F79E465",
    x"3F79E5C2",
    x"3F79E71F",
    x"3F79E87C",
    x"3F79E9D9",
    x"3F79EB36",
    x"3F79EC92",
    x"3F79EDEE",
    x"3F79EF4A",
    x"3F79F0A6",
    x"3F79F202",
    x"3F79F35E",
    x"3F79F4B9",
    x"3F79F615",
    x"3F79F770",
    x"3F79F8CB",
    x"3F79FA26",
    x"3F79FB81",
    x"3F79FCDB",
    x"3F79FE36",
    x"3F79FF90",
    x"3F7A00EA",
    x"3F7A0244",
    x"3F7A039E",
    x"3F7A04F8",
    x"3F7A0652",
    x"3F7A07AB",
    x"3F7A0904",
    x"3F7A0A5D",
    x"3F7A0BB6",
    x"3F7A0D0F",
    x"3F7A0E68",
    x"3F7A0FC0",
    x"3F7A1119",
    x"3F7A1271",
    x"3F7A13C9",
    x"3F7A1521",
    x"3F7A1679",
    x"3F7A17D0",
    x"3F7A1928",
    x"3F7A1A7F",
    x"3F7A1BD6",
    x"3F7A1D2D",
    x"3F7A1E84",
    x"3F7A1FDB",
    x"3F7A2131",
    x"3F7A2288",
    x"3F7A23DE",
    x"3F7A2534",
    x"3F7A268A",
    x"3F7A27E0",
    x"3F7A2936",
    x"3F7A2A8B",
    x"3F7A2BE1",
    x"3F7A2D36",
    x"3F7A2E8B",
    x"3F7A2FE0",
    x"3F7A3134",
    x"3F7A3289",
    x"3F7A33DD",
    x"3F7A3532",
    x"3F7A3686",
    x"3F7A37DA",
    x"3F7A392E",
    x"3F7A3A81",
    x"3F7A3BD5",
    x"3F7A3D28",
    x"3F7A3E7C",
    x"3F7A3FCF",
    x"3F7A4122",
    x"3F7A4275",
    x"3F7A43C7",
    x"3F7A451A",
    x"3F7A466C",
    x"3F7A47BE",
    x"3F7A4910",
    x"3F7A4A62",
    x"3F7A4BB4",
    x"3F7A4D05",
    x"3F7A4E57",
    x"3F7A4FA8",
    x"3F7A50F9",
    x"3F7A524A",
    x"3F7A539B",
    x"3F7A54EC",
    x"3F7A563C",
    x"3F7A578D",
    x"3F7A58DD",
    x"3F7A5A2D",
    x"3F7A5B7D",
    x"3F7A5CCD",
    x"3F7A5E1C",
    x"3F7A5F6C",
    x"3F7A60BB",
    x"3F7A620A",
    x"3F7A6359",
    x"3F7A64A8",
    x"3F7A65F7",
    x"3F7A6745",
    x"3F7A6894",
    x"3F7A69E2",
    x"3F7A6B30",
    x"3F7A6C7E",
    x"3F7A6DCC",
    x"3F7A6F1A",
    x"3F7A7067",
    x"3F7A71B5",
    x"3F7A7302",
    x"3F7A744F",
    x"3F7A759C",
    x"3F7A76E9",
    x"3F7A7835",
    x"3F7A7982",
    x"3F7A7ACE",
    x"3F7A7C1A",
    x"3F7A7D66",
    x"3F7A7EB2",
    x"3F7A7FFE",
    x"3F7A8149",
    x"3F7A8295",
    x"3F7A83E0",
    x"3F7A852B",
    x"3F7A8676",
    x"3F7A87C1",
    x"3F7A890B",
    x"3F7A8A56",
    x"3F7A8BA0",
    x"3F7A8CEA",
    x"3F7A8E34",
    x"3F7A8F7E",
    x"3F7A90C8",
    x"3F7A9212",
    x"3F7A935B",
    x"3F7A94A4",
    x"3F7A95EE",
    x"3F7A9737",
    x"3F7A987F",
    x"3F7A99C8",
    x"3F7A9B11",
    x"3F7A9C59",
    x"3F7A9DA1",
    x"3F7A9EE9",
    x"3F7AA031",
    x"3F7AA179",
    x"3F7AA2C1",
    x"3F7AA408",
    x"3F7AA54F",
    x"3F7AA697",
    x"3F7AA7DE",
    x"3F7AA925",
    x"3F7AAA6B",
    x"3F7AABB2",
    x"3F7AACF8",
    x"3F7AAE3F",
    x"3F7AAF85",
    x"3F7AB0CB",
    x"3F7AB210",
    x"3F7AB356",
    x"3F7AB49C",
    x"3F7AB5E1",
    x"3F7AB726",
    x"3F7AB86B",
    x"3F7AB9B0",
    x"3F7ABAF5",
    x"3F7ABC3A",
    x"3F7ABD7E",
    x"3F7ABEC2",
    x"3F7AC006",
    x"3F7AC14A",
    x"3F7AC28E",
    x"3F7AC3D2",
    x"3F7AC516",
    x"3F7AC659",
    x"3F7AC79C",
    x"3F7AC8DF",
    x"3F7ACA22",
    x"3F7ACB65",
    x"3F7ACCA8",
    x"3F7ACDEA",
    x"3F7ACF2D",
    x"3F7AD06F",
    x"3F7AD1B1",
    x"3F7AD2F3",
    x"3F7AD434",
    x"3F7AD576",
    x"3F7AD6B7",
    x"3F7AD7F9",
    x"3F7AD93A",
    x"3F7ADA7B",
    x"3F7ADBBC",
    x"3F7ADCFC",
    x"3F7ADE3D",
    x"3F7ADF7D",
    x"3F7AE0BD",
    x"3F7AE1FE",
    x"3F7AE33D",
    x"3F7AE47D",
    x"3F7AE5BD",
    x"3F7AE6FC",
    x"3F7AE83C",
    x"3F7AE97B",
    x"3F7AEABA",
    x"3F7AEBF9",
    x"3F7AED37",
    x"3F7AEE76",
    x"3F7AEFB4",
    x"3F7AF0F3",
    x"3F7AF231",
    x"3F7AF36F",
    x"3F7AF4AD",
    x"3F7AF5EA",
    x"3F7AF728",
    x"3F7AF865",
    x"3F7AF9A2",
    x"3F7AFADF",
    x"3F7AFC1C",
    x"3F7AFD59",
    x"3F7AFE96",
    x"3F7AFFD2",
    x"3F7B010E",
    x"3F7B024A",
    x"3F7B0386",
    x"3F7B04C2",
    x"3F7B05FE",
    x"3F7B073A",
    x"3F7B0875",
    x"3F7B09B0",
    x"3F7B0AEB",
    x"3F7B0C26",
    x"3F7B0D61",
    x"3F7B0E9C",
    x"3F7B0FD6",
    x"3F7B1110",
    x"3F7B124B",
    x"3F7B1385",
    x"3F7B14BE",
    x"3F7B15F8",
    x"3F7B1732",
    x"3F7B186B",
    x"3F7B19A4",
    x"3F7B1ADE",
    x"3F7B1C17",
    x"3F7B1D4F",
    x"3F7B1E88",
    x"3F7B1FC1",
    x"3F7B20F9",
    x"3F7B2231",
    x"3F7B2369",
    x"3F7B24A1",
    x"3F7B25D9",
    x"3F7B2711",
    x"3F7B2848",
    x"3F7B297F",
    x"3F7B2AB6",
    x"3F7B2BED",
    x"3F7B2D24",
    x"3F7B2E5B",
    x"3F7B2F92",
    x"3F7B30C8",
    x"3F7B31FE",
    x"3F7B3334",
    x"3F7B346A",
    x"3F7B35A0",
    x"3F7B36D6",
    x"3F7B380B",
    x"3F7B3940",
    x"3F7B3A76",
    x"3F7B3BAB",
    x"3F7B3CE0",
    x"3F7B3E14",
    x"3F7B3F49",
    x"3F7B407D",
    x"3F7B41B2",
    x"3F7B42E6",
    x"3F7B441A",
    x"3F7B454E",
    x"3F7B4681",
    x"3F7B47B5",
    x"3F7B48E8",
    x"3F7B4A1B",
    x"3F7B4B4E",
    x"3F7B4C81",
    x"3F7B4DB4",
    x"3F7B4EE7",
    x"3F7B5019",
    x"3F7B514B",
    x"3F7B527E",
    x"3F7B53B0",
    x"3F7B54E1",
    x"3F7B5613",
    x"3F7B5745",
    x"3F7B5876",
    x"3F7B59A7",
    x"3F7B5AD9",
    x"3F7B5C09",
    x"3F7B5D3A",
    x"3F7B5E6B",
    x"3F7B5F9B",
    x"3F7B60CC",
    x"3F7B61FC",
    x"3F7B632C",
    x"3F7B645C",
    x"3F7B658C",
    x"3F7B66BB",
    x"3F7B67EB",
    x"3F7B691A",
    x"3F7B6A49",
    x"3F7B6B78",
    x"3F7B6CA7",
    x"3F7B6DD6",
    x"3F7B6F04",
    x"3F7B7032",
    x"3F7B7161",
    x"3F7B728F",
    x"3F7B73BD",
    x"3F7B74EA",
    x"3F7B7618",
    x"3F7B7745",
    x"3F7B7873",
    x"3F7B79A0",
    x"3F7B7ACD",
    x"3F7B7BFA",
    x"3F7B7D27",
    x"3F7B7E53",
    x"3F7B7F80",
    x"3F7B80AC",
    x"3F7B81D8",
    x"3F7B8304",
    x"3F7B8430",
    x"3F7B855B",
    x"3F7B8687",
    x"3F7B87B2",
    x"3F7B88DD",
    x"3F7B8A08",
    x"3F7B8B33",
    x"3F7B8C5E",
    x"3F7B8D89",
    x"3F7B8EB3",
    x"3F7B8FDD",
    x"3F7B9107",
    x"3F7B9231",
    x"3F7B935B",
    x"3F7B9485",
    x"3F7B95AE",
    x"3F7B96D8",
    x"3F7B9801",
    x"3F7B992A",
    x"3F7B9A53",
    x"3F7B9B7C",
    x"3F7B9CA4",
    x"3F7B9DCD",
    x"3F7B9EF5",
    x"3F7BA01D",
    x"3F7BA145",
    x"3F7BA26D",
    x"3F7BA395",
    x"3F7BA4BC",
    x"3F7BA5E4",
    x"3F7BA70B",
    x"3F7BA832",
    x"3F7BA959",
    x"3F7BAA80",
    x"3F7BABA7",
    x"3F7BACCD",
    x"3F7BADF3",
    x"3F7BAF1A",
    x"3F7BB040",
    x"3F7BB166",
    x"3F7BB28B",
    x"3F7BB3B1",
    x"3F7BB4D6",
    x"3F7BB5FC",
    x"3F7BB721",
    x"3F7BB846",
    x"3F7BB96B",
    x"3F7BBA8F",
    x"3F7BBBB4",
    x"3F7BBCD8",
    x"3F7BBDFC",
    x"3F7BBF20",
    x"3F7BC044",
    x"3F7BC168",
    x"3F7BC28C",
    x"3F7BC3AF",
    x"3F7BC4D2",
    x"3F7BC5F6",
    x"3F7BC719",
    x"3F7BC83B",
    x"3F7BC95E",
    x"3F7BCA81",
    x"3F7BCBA3",
    x"3F7BCCC5",
    x"3F7BCDE7",
    x"3F7BCF09",
    x"3F7BD02B",
    x"3F7BD14D",
    x"3F7BD26E",
    x"3F7BD390",
    x"3F7BD4B1",
    x"3F7BD5D2",
    x"3F7BD6F3",
    x"3F7BD814",
    x"3F7BD934",
    x"3F7BDA55",
    x"3F7BDB75",
    x"3F7BDC95",
    x"3F7BDDB5",
    x"3F7BDED5",
    x"3F7BDFF4",
    x"3F7BE114",
    x"3F7BE233",
    x"3F7BE353",
    x"3F7BE472",
    x"3F7BE590",
    x"3F7BE6AF",
    x"3F7BE7CE",
    x"3F7BE8EC",
    x"3F7BEA0B",
    x"3F7BEB29",
    x"3F7BEC47",
    x"3F7BED65",
    x"3F7BEE82",
    x"3F7BEFA0",
    x"3F7BF0BD",
    x"3F7BF1DA",
    x"3F7BF2F8",
    x"3F7BF415",
    x"3F7BF531",
    x"3F7BF64E",
    x"3F7BF76A",
    x"3F7BF887",
    x"3F7BF9A3",
    x"3F7BFABF",
    x"3F7BFBDB",
    x"3F7BFCF7",
    x"3F7BFE12",
    x"3F7BFF2E",
    x"3F7C0049",
    x"3F7C0164",
    x"3F7C027F",
    x"3F7C039A",
    x"3F7C04B4",
    x"3F7C05CF",
    x"3F7C06E9",
    x"3F7C0803",
    x"3F7C091E",
    x"3F7C0A37",
    x"3F7C0B51",
    x"3F7C0C6B",
    x"3F7C0D84",
    x"3F7C0E9D",
    x"3F7C0FB7",
    x"3F7C10D0",
    x"3F7C11E8",
    x"3F7C1301",
    x"3F7C141A",
    x"3F7C1532",
    x"3F7C164A",
    x"3F7C1762",
    x"3F7C187A",
    x"3F7C1992",
    x"3F7C1AAA",
    x"3F7C1BC1",
    x"3F7C1CD9",
    x"3F7C1DF0",
    x"3F7C1F07",
    x"3F7C201E",
    x"3F7C2134",
    x"3F7C224B",
    x"3F7C2361",
    x"3F7C2478",
    x"3F7C258E",
    x"3F7C26A4",
    x"3F7C27B9",
    x"3F7C28CF",
    x"3F7C29E5",
    x"3F7C2AFA",
    x"3F7C2C0F",
    x"3F7C2D24",
    x"3F7C2E39",
    x"3F7C2F4E",
    x"3F7C3062",
    x"3F7C3177",
    x"3F7C328B",
    x"3F7C339F",
    x"3F7C34B3",
    x"3F7C35C7",
    x"3F7C36DB",
    x"3F7C37EE",
    x"3F7C3902",
    x"3F7C3A15",
    x"3F7C3B28",
    x"3F7C3C3B",
    x"3F7C3D4E",
    x"3F7C3E60",
    x"3F7C3F73",
    x"3F7C4085",
    x"3F7C4197",
    x"3F7C42A9",
    x"3F7C43BB",
    x"3F7C44CD",
    x"3F7C45DE",
    x"3F7C46F0",
    x"3F7C4801",
    x"3F7C4912",
    x"3F7C4A23",
    x"3F7C4B34",
    x"3F7C4C44",
    x"3F7C4D55",
    x"3F7C4E65",
    x"3F7C4F75",
    x"3F7C5085",
    x"3F7C5195",
    x"3F7C52A5",
    x"3F7C53B4",
    x"3F7C54C4",
    x"3F7C55D3",
    x"3F7C56E2",
    x"3F7C57F1",
    x"3F7C5900",
    x"3F7C5A0F",
    x"3F7C5B1D",
    x"3F7C5C2C",
    x"3F7C5D3A",
    x"3F7C5E48",
    x"3F7C5F56",
    x"3F7C6063",
    x"3F7C6171",
    x"3F7C627E",
    x"3F7C638C",
    x"3F7C6499",
    x"3F7C65A6",
    x"3F7C66B3",
    x"3F7C67BF",
    x"3F7C68CC",
    x"3F7C69D8",
    x"3F7C6AE5",
    x"3F7C6BF1",
    x"3F7C6CFD",
    x"3F7C6E08",
    x"3F7C6F14",
    x"3F7C701F",
    x"3F7C712B",
    x"3F7C7236",
    x"3F7C7341",
    x"3F7C744C",
    x"3F7C7556",
    x"3F7C7661",
    x"3F7C776B",
    x"3F7C7876",
    x"3F7C7980",
    x"3F7C7A8A",
    x"3F7C7B94",
    x"3F7C7C9D",
    x"3F7C7DA7",
    x"3F7C7EB0",
    x"3F7C7FB9",
    x"3F7C80C2",
    x"3F7C81CB",
    x"3F7C82D4",
    x"3F7C83DC",
    x"3F7C84E5",
    x"3F7C85ED",
    x"3F7C86F5",
    x"3F7C87FD",
    x"3F7C8905",
    x"3F7C8A0D",
    x"3F7C8B14",
    x"3F7C8C1C",
    x"3F7C8D23",
    x"3F7C8E2A",
    x"3F7C8F31",
    x"3F7C9037",
    x"3F7C913E",
    x"3F7C9245",
    x"3F7C934B",
    x"3F7C9451",
    x"3F7C9557",
    x"3F7C965D",
    x"3F7C9762",
    x"3F7C9868",
    x"3F7C996D",
    x"3F7C9A73",
    x"3F7C9B78",
    x"3F7C9C7D",
    x"3F7C9D81",
    x"3F7C9E86",
    x"3F7C9F8A",
    x"3F7CA08F",
    x"3F7CA193",
    x"3F7CA297",
    x"3F7CA39B",
    x"3F7CA49F",
    x"3F7CA5A2",
    x"3F7CA6A6",
    x"3F7CA7A9",
    x"3F7CA8AC",
    x"3F7CA9AF",
    x"3F7CAAB2",
    x"3F7CABB4",
    x"3F7CACB7",
    x"3F7CADB9",
    x"3F7CAEBB",
    x"3F7CAFBD",
    x"3F7CB0BF",
    x"3F7CB1C1",
    x"3F7CB2C2",
    x"3F7CB3C4",
    x"3F7CB4C5",
    x"3F7CB5C6",
    x"3F7CB6C7",
    x"3F7CB7C8",
    x"3F7CB8C9",
    x"3F7CB9C9",
    x"3F7CBACA",
    x"3F7CBBCA",
    x"3F7CBCCA",
    x"3F7CBDCA",
    x"3F7CBECA",
    x"3F7CBFC9",
    x"3F7CC0C9",
    x"3F7CC1C8",
    x"3F7CC2C7",
    x"3F7CC3C6",
    x"3F7CC4C5",
    x"3F7CC5C4",
    x"3F7CC6C2",
    x"3F7CC7C0",
    x"3F7CC8BF",
    x"3F7CC9BD",
    x"3F7CCABB",
    x"3F7CCBB8",
    x"3F7CCCB6",
    x"3F7CCDB4",
    x"3F7CCEB1",
    x"3F7CCFAE",
    x"3F7CD0AB",
    x"3F7CD1A8",
    x"3F7CD2A5",
    x"3F7CD3A1",
    x"3F7CD49E",
    x"3F7CD59A",
    x"3F7CD696",
    x"3F7CD792",
    x"3F7CD88E",
    x"3F7CD989",
    x"3F7CDA85",
    x"3F7CDB80",
    x"3F7CDC7B",
    x"3F7CDD76",
    x"3F7CDE71",
    x"3F7CDF6C",
    x"3F7CE066",
    x"3F7CE161",
    x"3F7CE25B",
    x"3F7CE355",
    x"3F7CE44F",
    x"3F7CE549",
    x"3F7CE643",
    x"3F7CE73C",
    x"3F7CE836",
    x"3F7CE92F",
    x"3F7CEA28",
    x"3F7CEB21",
    x"3F7CEC19",
    x"3F7CED12",
    x"3F7CEE0B",
    x"3F7CEF03",
    x"3F7CEFFB",
    x"3F7CF0F3",
    x"3F7CF1EB",
    x"3F7CF2E2",
    x"3F7CF3DA",
    x"3F7CF4D1",
    x"3F7CF5C9",
    x"3F7CF6C0",
    x"3F7CF7B7",
    x"3F7CF8AD",
    x"3F7CF9A4",
    x"3F7CFA9A",
    x"3F7CFB91",
    x"3F7CFC87",
    x"3F7CFD7D",
    x"3F7CFE73",
    x"3F7CFF68",
    x"3F7D005E",
    x"3F7D0153",
    x"3F7D0249",
    x"3F7D033E",
    x"3F7D0433",
    x"3F7D0527",
    x"3F7D061C",
    x"3F7D0710",
    x"3F7D0805",
    x"3F7D08F9",
    x"3F7D09ED",
    x"3F7D0AE1",
    x"3F7D0BD5",
    x"3F7D0CC8",
    x"3F7D0DBC",
    x"3F7D0EAF",
    x"3F7D0FA2",
    x"3F7D1095",
    x"3F7D1188",
    x"3F7D127A",
    x"3F7D136D",
    x"3F7D145F",
    x"3F7D1551",
    x"3F7D1643",
    x"3F7D1735",
    x"3F7D1827",
    x"3F7D1919",
    x"3F7D1A0A",
    x"3F7D1AFB",
    x"3F7D1BEC",
    x"3F7D1CDD",
    x"3F7D1DCE",
    x"3F7D1EBF",
    x"3F7D1FAF",
    x"3F7D20A0",
    x"3F7D2190",
    x"3F7D2280",
    x"3F7D2370",
    x"3F7D2460",
    x"3F7D254F",
    x"3F7D263F",
    x"3F7D272E",
    x"3F7D281D",
    x"3F7D290C",
    x"3F7D29FB",
    x"3F7D2AEA",
    x"3F7D2BD8",
    x"3F7D2CC7",
    x"3F7D2DB5",
    x"3F7D2EA3",
    x"3F7D2F91",
    x"3F7D307F",
    x"3F7D316C",
    x"3F7D325A",
    x"3F7D3347",
    x"3F7D3434",
    x"3F7D3521",
    x"3F7D360E",
    x"3F7D36FB",
    x"3F7D37E7",
    x"3F7D38D4",
    x"3F7D39C0",
    x"3F7D3AAC",
    x"3F7D3B98",
    x"3F7D3C84",
    x"3F7D3D6F",
    x"3F7D3E5B",
    x"3F7D3F46",
    x"3F7D4031",
    x"3F7D411C",
    x"3F7D4207",
    x"3F7D42F2",
    x"3F7D43DC",
    x"3F7D44C7",
    x"3F7D45B1",
    x"3F7D469B",
    x"3F7D4785",
    x"3F7D486F",
    x"3F7D4959",
    x"3F7D4A42",
    x"3F7D4B2C",
    x"3F7D4C15",
    x"3F7D4CFE",
    x"3F7D4DE7",
    x"3F7D4ECF",
    x"3F7D4FB8",
    x"3F7D50A0",
    x"3F7D5189",
    x"3F7D5271",
    x"3F7D5359",
    x"3F7D5441",
    x"3F7D5528",
    x"3F7D5610",
    x"3F7D56F7",
    x"3F7D57DE",
    x"3F7D58C5",
    x"3F7D59AC",
    x"3F7D5A93",
    x"3F7D5B7A",
    x"3F7D5C60",
    x"3F7D5D46",
    x"3F7D5E2D",
    x"3F7D5F13",
    x"3F7D5FF8",
    x"3F7D60DE",
    x"3F7D61C4",
    x"3F7D62A9",
    x"3F7D638E",
    x"3F7D6473",
    x"3F7D6558",
    x"3F7D663D",
    x"3F7D6722",
    x"3F7D6806",
    x"3F7D68EA",
    x"3F7D69CE",
    x"3F7D6AB2",
    x"3F7D6B96",
    x"3F7D6C7A",
    x"3F7D6D5E",
    x"3F7D6E41",
    x"3F7D6F24",
    x"3F7D7007",
    x"3F7D70EA",
    x"3F7D71CD",
    x"3F7D72B0",
    x"3F7D7392",
    x"3F7D7474",
    x"3F7D7557",
    x"3F7D7639",
    x"3F7D771B",
    x"3F7D77FC",
    x"3F7D78DE",
    x"3F7D79BF",
    x"3F7D7AA0",
    x"3F7D7B82",
    x"3F7D7C62",
    x"3F7D7D43",
    x"3F7D7E24",
    x"3F7D7F04",
    x"3F7D7FE5",
    x"3F7D80C5",
    x"3F7D81A5",
    x"3F7D8285",
    x"3F7D8365",
    x"3F7D8444",
    x"3F7D8524",
    x"3F7D8603",
    x"3F7D86E2",
    x"3F7D87C1",
    x"3F7D88A0",
    x"3F7D897E",
    x"3F7D8A5D",
    x"3F7D8B3B",
    x"3F7D8C19",
    x"3F7D8CF8",
    x"3F7D8DD5",
    x"3F7D8EB3",
    x"3F7D8F91",
    x"3F7D906E",
    x"3F7D914B",
    x"3F7D9229",
    x"3F7D9306",
    x"3F7D93E2",
    x"3F7D94BF",
    x"3F7D959C",
    x"3F7D9678",
    x"3F7D9754",
    x"3F7D9830",
    x"3F7D990C",
    x"3F7D99E8",
    x"3F7D9AC4",
    x"3F7D9B9F",
    x"3F7D9C7A",
    x"3F7D9D55",
    x"3F7D9E30",
    x"3F7D9F0B",
    x"3F7D9FE6",
    x"3F7DA0C0",
    x"3F7DA19B",
    x"3F7DA275",
    x"3F7DA34F",
    x"3F7DA429",
    x"3F7DA503",
    x"3F7DA5DC",
    x"3F7DA6B6",
    x"3F7DA78F",
    x"3F7DA868",
    x"3F7DA941",
    x"3F7DAA1A",
    x"3F7DAAF3",
    x"3F7DABCC",
    x"3F7DACA4",
    x"3F7DAD7C",
    x"3F7DAE54",
    x"3F7DAF2C",
    x"3F7DB004",
    x"3F7DB0DC",
    x"3F7DB1B3",
    x"3F7DB28A",
    x"3F7DB362",
    x"3F7DB439",
    x"3F7DB510",
    x"3F7DB5E6",
    x"3F7DB6BD",
    x"3F7DB793",
    x"3F7DB869",
    x"3F7DB940",
    x"3F7DBA15",
    x"3F7DBAEB",
    x"3F7DBBC1",
    x"3F7DBC96",
    x"3F7DBD6C",
    x"3F7DBE41",
    x"3F7DBF16",
    x"3F7DBFEB",
    x"3F7DC0C0",
    x"3F7DC194",
    x"3F7DC269",
    x"3F7DC33D",
    x"3F7DC411",
    x"3F7DC4E5",
    x"3F7DC5B9",
    x"3F7DC68C",
    x"3F7DC760",
    x"3F7DC833",
    x"3F7DC906",
    x"3F7DC9DA",
    x"3F7DCAAC",
    x"3F7DCB7F",
    x"3F7DCC52",
    x"3F7DCD24",
    x"3F7DCDF6",
    x"3F7DCEC9",
    x"3F7DCF9B",
    x"3F7DD06C",
    x"3F7DD13E",
    x"3F7DD210",
    x"3F7DD2E1",
    x"3F7DD3B2",
    x"3F7DD483",
    x"3F7DD554",
    x"3F7DD625",
    x"3F7DD6F5",
    x"3F7DD7C6",
    x"3F7DD896",
    x"3F7DD966",
    x"3F7DDA36",
    x"3F7DDB06",
    x"3F7DDBD6",
    x"3F7DDCA5",
    x"3F7DDD75",
    x"3F7DDE44",
    x"3F7DDF13",
    x"3F7DDFE2",
    x"3F7DE0B1",
    x"3F7DE17F",
    x"3F7DE24E",
    x"3F7DE31C",
    x"3F7DE3EA",
    x"3F7DE4B8",
    x"3F7DE586",
    x"3F7DE654",
    x"3F7DE721",
    x"3F7DE7EF",
    x"3F7DE8BC",
    x"3F7DE989",
    x"3F7DEA56",
    x"3F7DEB23",
    x"3F7DEBEF",
    x"3F7DECBC",
    x"3F7DED88",
    x"3F7DEE54",
    x"3F7DEF20",
    x"3F7DEFEC",
    x"3F7DF0B8",
    x"3F7DF183",
    x"3F7DF24F",
    x"3F7DF31A",
    x"3F7DF3E5",
    x"3F7DF4B0",
    x"3F7DF57B",
    x"3F7DF646",
    x"3F7DF710",
    x"3F7DF7DA",
    x"3F7DF8A5",
    x"3F7DF96F",
    x"3F7DFA38",
    x"3F7DFB02",
    x"3F7DFBCC",
    x"3F7DFC95",
    x"3F7DFD5E",
    x"3F7DFE28",
    x"3F7DFEF0",
    x"3F7DFFB9",
    x"3F7E0082",
    x"3F7E014A",
    x"3F7E0213",
    x"3F7E02DB",
    x"3F7E03A3",
    x"3F7E046B",
    x"3F7E0533",
    x"3F7E05FA",
    x"3F7E06C2",
    x"3F7E0789",
    x"3F7E0850",
    x"3F7E0917",
    x"3F7E09DE",
    x"3F7E0AA4",
    x"3F7E0B6B",
    x"3F7E0C31",
    x"3F7E0CF7",
    x"3F7E0DBD",
    x"3F7E0E83",
    x"3F7E0F49",
    x"3F7E100F",
    x"3F7E10D4",
    x"3F7E1199",
    x"3F7E125F",
    x"3F7E1324",
    x"3F7E13E8",
    x"3F7E14AD",
    x"3F7E1572",
    x"3F7E1636",
    x"3F7E16FA",
    x"3F7E17BE",
    x"3F7E1882",
    x"3F7E1946",
    x"3F7E1A09",
    x"3F7E1ACD",
    x"3F7E1B90",
    x"3F7E1C53",
    x"3F7E1D16",
    x"3F7E1DD9",
    x"3F7E1E9C",
    x"3F7E1F5E",
    x"3F7E2021",
    x"3F7E20E3",
    x"3F7E21A5",
    x"3F7E2267",
    x"3F7E2329",
    x"3F7E23EA",
    x"3F7E24AC",
    x"3F7E256D",
    x"3F7E262E",
    x"3F7E26EF",
    x"3F7E27B0",
    x"3F7E2871",
    x"3F7E2931",
    x"3F7E29F2",
    x"3F7E2AB2",
    x"3F7E2B72",
    x"3F7E2C32",
    x"3F7E2CF2",
    x"3F7E2DB1",
    x"3F7E2E71",
    x"3F7E2F30",
    x"3F7E2FEF",
    x"3F7E30AE",
    x"3F7E316D",
    x"3F7E322C",
    x"3F7E32EA",
    x"3F7E33A9",
    x"3F7E3467",
    x"3F7E3525",
    x"3F7E35E3",
    x"3F7E36A1",
    x"3F7E375E",
    x"3F7E381C",
    x"3F7E38D9",
    x"3F7E3996",
    x"3F7E3A53",
    x"3F7E3B10",
    x"3F7E3BCD",
    x"3F7E3C89",
    x"3F7E3D46",
    x"3F7E3E02",
    x"3F7E3EBE",
    x"3F7E3F7A",
    x"3F7E4036",
    x"3F7E40F1",
    x"3F7E41AD",
    x"3F7E4268",
    x"3F7E4323",
    x"3F7E43DE",
    x"3F7E4499",
    x"3F7E4554",
    x"3F7E460F",
    x"3F7E46C9",
    x"3F7E4783",
    x"3F7E483D",
    x"3F7E48F7",
    x"3F7E49B1",
    x"3F7E4A6B",
    x"3F7E4B24",
    x"3F7E4BDE",
    x"3F7E4C97",
    x"3F7E4D50",
    x"3F7E4E09",
    x"3F7E4EC1",
    x"3F7E4F7A",
    x"3F7E5032",
    x"3F7E50EB",
    x"3F7E51A3",
    x"3F7E525B",
    x"3F7E5312",
    x"3F7E53CA",
    x"3F7E5482",
    x"3F7E5539",
    x"3F7E55F0",
    x"3F7E56A7",
    x"3F7E575E",
    x"3F7E5815",
    x"3F7E58CB",
    x"3F7E5982",
    x"3F7E5A38",
    x"3F7E5AEE",
    x"3F7E5BA4",
    x"3F7E5C5A",
    x"3F7E5D10",
    x"3F7E5DC5",
    x"3F7E5E7B",
    x"3F7E5F30",
    x"3F7E5FE5",
    x"3F7E609A",
    x"3F7E614E",
    x"3F7E6203",
    x"3F7E62B7",
    x"3F7E636C",
    x"3F7E6420",
    x"3F7E64D4",
    x"3F7E6588",
    x"3F7E663B",
    x"3F7E66EF",
    x"3F7E67A2",
    x"3F7E6855",
    x"3F7E6908",
    x"3F7E69BB",
    x"3F7E6A6E",
    x"3F7E6B21",
    x"3F7E6BD3",
    x"3F7E6C85",
    x"3F7E6D38",
    x"3F7E6DEA",
    x"3F7E6E9B",
    x"3F7E6F4D",
    x"3F7E6FFF",
    x"3F7E70B0",
    x"3F7E7161",
    x"3F7E7212",
    x"3F7E72C3",
    x"3F7E7374",
    x"3F7E7424",
    x"3F7E74D5",
    x"3F7E7585",
    x"3F7E7635",
    x"3F7E76E5",
    x"3F7E7795",
    x"3F7E7845",
    x"3F7E78F4",
    x"3F7E79A4",
    x"3F7E7A53",
    x"3F7E7B02",
    x"3F7E7BB1",
    x"3F7E7C60",
    x"3F7E7D0E",
    x"3F7E7DBD",
    x"3F7E7E6B",
    x"3F7E7F19",
    x"3F7E7FC7",
    x"3F7E8075",
    x"3F7E8123",
    x"3F7E81D0",
    x"3F7E827E",
    x"3F7E832B",
    x"3F7E83D8",
    x"3F7E8485",
    x"3F7E8532",
    x"3F7E85DE",
    x"3F7E868B",
    x"3F7E8737",
    x"3F7E87E3",
    x"3F7E888F",
    x"3F7E893B",
    x"3F7E89E7",
    x"3F7E8A92",
    x"3F7E8B3E",
    x"3F7E8BE9",
    x"3F7E8C94",
    x"3F7E8D3F",
    x"3F7E8DEA",
    x"3F7E8E94",
    x"3F7E8F3F",
    x"3F7E8FE9",
    x"3F7E9093",
    x"3F7E913D",
    x"3F7E91E7",
    x"3F7E9291",
    x"3F7E933A",
    x"3F7E93E4",
    x"3F7E948D",
    x"3F7E9536",
    x"3F7E95DF",
    x"3F7E9688",
    x"3F7E9731",
    x"3F7E97D9",
    x"3F7E9881",
    x"3F7E9929",
    x"3F7E99D2",
    x"3F7E9A79",
    x"3F7E9B21",
    x"3F7E9BC9",
    x"3F7E9C70",
    x"3F7E9D17",
    x"3F7E9DBE",
    x"3F7E9E65",
    x"3F7E9F0C",
    x"3F7E9FB3",
    x"3F7EA059",
    x"3F7EA100",
    x"3F7EA1A6",
    x"3F7EA24C",
    x"3F7EA2F2",
    x"3F7EA397",
    x"3F7EA43D",
    x"3F7EA4E2",
    x"3F7EA588",
    x"3F7EA62D",
    x"3F7EA6D2",
    x"3F7EA776",
    x"3F7EA81B",
    x"3F7EA8C0",
    x"3F7EA964",
    x"3F7EAA08",
    x"3F7EAAAC",
    x"3F7EAB50",
    x"3F7EABF4",
    x"3F7EAC97",
    x"3F7EAD3B",
    x"3F7EADDE",
    x"3F7EAE81",
    x"3F7EAF24",
    x"3F7EAFC7",
    x"3F7EB069",
    x"3F7EB10C",
    x"3F7EB1AE",
    x"3F7EB250",
    x"3F7EB2F2",
    x"3F7EB394",
    x"3F7EB436",
    x"3F7EB4D8",
    x"3F7EB579",
    x"3F7EB61A",
    x"3F7EB6BB",
    x"3F7EB75C",
    x"3F7EB7FD",
    x"3F7EB89E",
    x"3F7EB93E",
    x"3F7EB9DF",
    x"3F7EBA7F",
    x"3F7EBB1F",
    x"3F7EBBBF",
    x"3F7EBC5F",
    x"3F7EBCFE",
    x"3F7EBD9E",
    x"3F7EBE3D",
    x"3F7EBEDC",
    x"3F7EBF7B",
    x"3F7EC01A",
    x"3F7EC0B8",
    x"3F7EC157",
    x"3F7EC1F5",
    x"3F7EC293",
    x"3F7EC331",
    x"3F7EC3CF",
    x"3F7EC46D",
    x"3F7EC50B",
    x"3F7EC5A8",
    x"3F7EC645",
    x"3F7EC6E3",
    x"3F7EC780",
    x"3F7EC81C",
    x"3F7EC8B9",
    x"3F7EC955",
    x"3F7EC9F2",
    x"3F7ECA8E",
    x"3F7ECB2A",
    x"3F7ECBC6",
    x"3F7ECC62",
    x"3F7ECCFD",
    x"3F7ECD99",
    x"3F7ECE34",
    x"3F7ECECF",
    x"3F7ECF6A",
    x"3F7ED005",
    x"3F7ED0A0",
    x"3F7ED13A",
    x"3F7ED1D4",
    x"3F7ED26F",
    x"3F7ED309",
    x"3F7ED3A3",
    x"3F7ED43C",
    x"3F7ED4D6",
    x"3F7ED56F",
    x"3F7ED609",
    x"3F7ED6A2",
    x"3F7ED73B",
    x"3F7ED7D4",
    x"3F7ED86C",
    x"3F7ED905",
    x"3F7ED99D",
    x"3F7EDA35",
    x"3F7EDACD",
    x"3F7EDB65",
    x"3F7EDBFD",
    x"3F7EDC95",
    x"3F7EDD2C",
    x"3F7EDDC3",
    x"3F7EDE5B",
    x"3F7EDEF2",
    x"3F7EDF88",
    x"3F7EE01F",
    x"3F7EE0B6",
    x"3F7EE14C",
    x"3F7EE1E2",
    x"3F7EE278",
    x"3F7EE30E",
    x"3F7EE3A4",
    x"3F7EE43A",
    x"3F7EE4CF",
    x"3F7EE564",
    x"3F7EE5F9",
    x"3F7EE68E",
    x"3F7EE723",
    x"3F7EE7B8",
    x"3F7EE84C",
    x"3F7EE8E1",
    x"3F7EE975",
    x"3F7EEA09",
    x"3F7EEA9D",
    x"3F7EEB31",
    x"3F7EEBC4",
    x"3F7EEC58",
    x"3F7EECEB",
    x"3F7EED7E",
    x"3F7EEE11",
    x"3F7EEEA4",
    x"3F7EEF37",
    x"3F7EEFC9",
    x"3F7EF05C",
    x"3F7EF0EE",
    x"3F7EF180",
    x"3F7EF212",
    x"3F7EF2A4",
    x"3F7EF335",
    x"3F7EF3C7",
    x"3F7EF458",
    x"3F7EF4E9",
    x"3F7EF57A",
    x"3F7EF60B",
    x"3F7EF69C",
    x"3F7EF72C",
    x"3F7EF7BD",
    x"3F7EF84D",
    x"3F7EF8DD",
    x"3F7EF96D",
    x"3F7EF9FD",
    x"3F7EFA8C",
    x"3F7EFB1C",
    x"3F7EFBAB",
    x"3F7EFC3A",
    x"3F7EFCC9",
    x"3F7EFD58",
    x"3F7EFDE7",
    x"3F7EFE75",
    x"3F7EFF04",
    x"3F7EFF92",
    x"3F7F0020",
    x"3F7F00AE",
    x"3F7F013C",
    x"3F7F01C9",
    x"3F7F0257",
    x"3F7F02E4",
    x"3F7F0371",
    x"3F7F03FE",
    x"3F7F048B",
    x"3F7F0518",
    x"3F7F05A4",
    x"3F7F0631",
    x"3F7F06BD",
    x"3F7F0749",
    x"3F7F07D5",
    x"3F7F0861",
    x"3F7F08EC",
    x"3F7F0978",
    x"3F7F0A03",
    x"3F7F0A8E",
    x"3F7F0B19",
    x"3F7F0BA4",
    x"3F7F0C2F",
    x"3F7F0CB9",
    x"3F7F0D44",
    x"3F7F0DCE",
    x"3F7F0E58",
    x"3F7F0EE2",
    x"3F7F0F6C",
    x"3F7F0FF5",
    x"3F7F107F",
    x"3F7F1108",
    x"3F7F1191",
    x"3F7F121A",
    x"3F7F12A3",
    x"3F7F132C",
    x"3F7F13B4",
    x"3F7F143D",
    x"3F7F14C5",
    x"3F7F154D",
    x"3F7F15D5",
    x"3F7F165D",
    x"3F7F16E4",
    x"3F7F176C",
    x"3F7F17F3",
    x"3F7F187A",
    x"3F7F1901",
    x"3F7F1988",
    x"3F7F1A0F",
    x"3F7F1A95",
    x"3F7F1B1C",
    x"3F7F1BA2",
    x"3F7F1C28",
    x"3F7F1CAE",
    x"3F7F1D34",
    x"3F7F1DB9",
    x"3F7F1E3F",
    x"3F7F1EC4",
    x"3F7F1F49",
    x"3F7F1FCE",
    x"3F7F2053",
    x"3F7F20D8",
    x"3F7F215C",
    x"3F7F21E1",
    x"3F7F2265",
    x"3F7F22E9",
    x"3F7F236D",
    x"3F7F23F1",
    x"3F7F2475",
    x"3F7F24F8",
    x"3F7F257B",
    x"3F7F25FF",
    x"3F7F2682",
    x"3F7F2704",
    x"3F7F2787",
    x"3F7F280A",
    x"3F7F288C",
    x"3F7F290E",
    x"3F7F2990",
    x"3F7F2A12",
    x"3F7F2A94",
    x"3F7F2B16",
    x"3F7F2B97",
    x"3F7F2C19",
    x"3F7F2C9A",
    x"3F7F2D1B",
    x"3F7F2D9C",
    x"3F7F2E1C",
    x"3F7F2E9D",
    x"3F7F2F1D",
    x"3F7F2F9D",
    x"3F7F301E",
    x"3F7F309E",
    x"3F7F311D",
    x"3F7F319D",
    x"3F7F321C",
    x"3F7F329C",
    x"3F7F331B",
    x"3F7F339A",
    x"3F7F3419",
    x"3F7F3497",
    x"3F7F3516",
    x"3F7F3594",
    x"3F7F3613",
    x"3F7F3691",
    x"3F7F370F",
    x"3F7F378C",
    x"3F7F380A",
    x"3F7F3888",
    x"3F7F3905",
    x"3F7F3982",
    x"3F7F39FF",
    x"3F7F3A7C",
    x"3F7F3AF9",
    x"3F7F3B75",
    x"3F7F3BF2",
    x"3F7F3C6E",
    x"3F7F3CEA",
    x"3F7F3D66",
    x"3F7F3DE2",
    x"3F7F3E5D",
    x"3F7F3ED9",
    x"3F7F3F54",
    x"3F7F3FCF",
    x"3F7F404A",
    x"3F7F40C5",
    x"3F7F4140",
    x"3F7F41BA",
    x"3F7F4235",
    x"3F7F42AF",
    x"3F7F4329",
    x"3F7F43A3",
    x"3F7F441D",
    x"3F7F4497",
    x"3F7F4510",
    x"3F7F4589",
    x"3F7F4603",
    x"3F7F467C",
    x"3F7F46F4",
    x"3F7F476D",
    x"3F7F47E6",
    x"3F7F485E",
    x"3F7F48D6",
    x"3F7F494E",
    x"3F7F49C6",
    x"3F7F4A3E",
    x"3F7F4AB6",
    x"3F7F4B2D",
    x"3F7F4BA5",
    x"3F7F4C1C",
    x"3F7F4C93",
    x"3F7F4D0A",
    x"3F7F4D80",
    x"3F7F4DF7",
    x"3F7F4E6D",
    x"3F7F4EE4",
    x"3F7F4F5A",
    x"3F7F4FD0",
    x"3F7F5045",
    x"3F7F50BB",
    x"3F7F5131",
    x"3F7F51A6",
    x"3F7F521B",
    x"3F7F5290",
    x"3F7F5305",
    x"3F7F537A",
    x"3F7F53EE",
    x"3F7F5463",
    x"3F7F54D7",
    x"3F7F554B",
    x"3F7F55BF",
    x"3F7F5633",
    x"3F7F56A6",
    x"3F7F571A",
    x"3F7F578D",
    x"3F7F5800",
    x"3F7F5873",
    x"3F7F58E6",
    x"3F7F5959",
    x"3F7F59CC",
    x"3F7F5A3E",
    x"3F7F5AB0",
    x"3F7F5B22",
    x"3F7F5B94",
    x"3F7F5C06",
    x"3F7F5C78",
    x"3F7F5CE9",
    x"3F7F5D5A",
    x"3F7F5DCC",
    x"3F7F5E3D",
    x"3F7F5EAE",
    x"3F7F5F1E",
    x"3F7F5F8F",
    x"3F7F5FFF",
    x"3F7F606F",
    x"3F7F60E0",
    x"3F7F6150",
    x"3F7F61BF",
    x"3F7F622F",
    x"3F7F629E",
    x"3F7F630E",
    x"3F7F637D",
    x"3F7F63EC",
    x"3F7F645B",
    x"3F7F64CA",
    x"3F7F6538",
    x"3F7F65A7",
    x"3F7F6615",
    x"3F7F6683",
    x"3F7F66F1",
    x"3F7F675F",
    x"3F7F67CC",
    x"3F7F683A",
    x"3F7F68A7",
    x"3F7F6914",
    x"3F7F6981",
    x"3F7F69EE",
    x"3F7F6A5B",
    x"3F7F6AC7",
    x"3F7F6B34",
    x"3F7F6BA0",
    x"3F7F6C0C",
    x"3F7F6C78",
    x"3F7F6CE4",
    x"3F7F6D50",
    x"3F7F6DBB",
    x"3F7F6E26",
    x"3F7F6E92",
    x"3F7F6EFD",
    x"3F7F6F67",
    x"3F7F6FD2",
    x"3F7F703D",
    x"3F7F70A7",
    x"3F7F7111",
    x"3F7F717B",
    x"3F7F71E5",
    x"3F7F724F",
    x"3F7F72B9",
    x"3F7F7322",
    x"3F7F738C",
    x"3F7F73F5",
    x"3F7F745E",
    x"3F7F74C7",
    x"3F7F752F",
    x"3F7F7598",
    x"3F7F7600",
    x"3F7F7669",
    x"3F7F76D1",
    x"3F7F7739",
    x"3F7F77A0",
    x"3F7F7808",
    x"3F7F7870",
    x"3F7F78D7",
    x"3F7F793E",
    x"3F7F79A5",
    x"3F7F7A0C",
    x"3F7F7A73",
    x"3F7F7AD9",
    x"3F7F7B40",
    x"3F7F7BA6",
    x"3F7F7C0C",
    x"3F7F7C72",
    x"3F7F7CD8",
    x"3F7F7D3D",
    x"3F7F7DA3",
    x"3F7F7E08",
    x"3F7F7E6D",
    x"3F7F7ED2",
    x"3F7F7F37",
    x"3F7F7F9C",
    x"3F7F8000",
    x"3F7F8065",
    x"3F7F80C9",
    x"3F7F812D",
    x"3F7F8191",
    x"3F7F81F5",
    x"3F7F8259",
    x"3F7F82BC",
    x"3F7F831F",
    x"3F7F8383",
    x"3F7F83E6",
    x"3F7F8448",
    x"3F7F84AB",
    x"3F7F850E",
    x"3F7F8570",
    x"3F7F85D2",
    x"3F7F8634",
    x"3F7F8696",
    x"3F7F86F8",
    x"3F7F875A",
    x"3F7F87BB",
    x"3F7F881D",
    x"3F7F887E",
    x"3F7F88DF",
    x"3F7F8940",
    x"3F7F89A0",
    x"3F7F8A01",
    x"3F7F8A61",
    x"3F7F8AC2",
    x"3F7F8B22",
    x"3F7F8B82",
    x"3F7F8BE1",
    x"3F7F8C41",
    x"3F7F8CA1",
    x"3F7F8D00",
    x"3F7F8D5F",
    x"3F7F8DBE",
    x"3F7F8E1D",
    x"3F7F8E7C",
    x"3F7F8EDA",
    x"3F7F8F39",
    x"3F7F8F97",
    x"3F7F8FF5",
    x"3F7F9053",
    x"3F7F90B1",
    x"3F7F910E",
    x"3F7F916C",
    x"3F7F91C9",
    x"3F7F9226",
    x"3F7F9283",
    x"3F7F92E0",
    x"3F7F933D",
    x"3F7F9399",
    x"3F7F93F6",
    x"3F7F9452",
    x"3F7F94AE",
    x"3F7F950A",
    x"3F7F9566",
    x"3F7F95C1",
    x"3F7F961D",
    x"3F7F9678",
    x"3F7F96D3",
    x"3F7F972E",
    x"3F7F9789",
    x"3F7F97E4",
    x"3F7F983F",
    x"3F7F9899",
    x"3F7F98F3",
    x"3F7F994D",
    x"3F7F99A7",
    x"3F7F9A01",
    x"3F7F9A5B",
    x"3F7F9AB4",
    x"3F7F9B0D",
    x"3F7F9B67",
    x"3F7F9BC0",
    x"3F7F9C18",
    x"3F7F9C71",
    x"3F7F9CCA",
    x"3F7F9D22",
    x"3F7F9D7A",
    x"3F7F9DD2",
    x"3F7F9E2A",
    x"3F7F9E82",
    x"3F7F9EDA",
    x"3F7F9F31",
    x"3F7F9F89",
    x"3F7F9FE0",
    x"3F7FA037",
    x"3F7FA08E",
    x"3F7FA0E4",
    x"3F7FA13B",
    x"3F7FA191",
    x"3F7FA1E8",
    x"3F7FA23E",
    x"3F7FA294",
    x"3F7FA2E9",
    x"3F7FA33F",
    x"3F7FA394",
    x"3F7FA3EA",
    x"3F7FA43F",
    x"3F7FA494",
    x"3F7FA4E9",
    x"3F7FA53D",
    x"3F7FA592",
    x"3F7FA5E6",
    x"3F7FA63B",
    x"3F7FA68F",
    x"3F7FA6E3",
    x"3F7FA736",
    x"3F7FA78A",
    x"3F7FA7DE",
    x"3F7FA831",
    x"3F7FA884",
    x"3F7FA8D7",
    x"3F7FA92A",
    x"3F7FA97D",
    x"3F7FA9CF",
    x"3F7FAA21",
    x"3F7FAA74",
    x"3F7FAAC6",
    x"3F7FAB18",
    x"3F7FAB6A",
    x"3F7FABBB",
    x"3F7FAC0D",
    x"3F7FAC5E",
    x"3F7FACAF",
    x"3F7FAD00",
    x"3F7FAD51",
    x"3F7FADA2",
    x"3F7FADF2",
    x"3F7FAE43",
    x"3F7FAE93",
    x"3F7FAEE3",
    x"3F7FAF33",
    x"3F7FAF83",
    x"3F7FAFD2",
    x"3F7FB022",
    x"3F7FB071",
    x"3F7FB0C0",
    x"3F7FB10F",
    x"3F7FB15E",
    x"3F7FB1AD",
    x"3F7FB1FB",
    x"3F7FB24A",
    x"3F7FB298",
    x"3F7FB2E6",
    x"3F7FB334",
    x"3F7FB382",
    x"3F7FB3CF",
    x"3F7FB41D",
    x"3F7FB46A",
    x"3F7FB4B7",
    x"3F7FB504",
    x"3F7FB551",
    x"3F7FB59E",
    x"3F7FB5EA",
    x"3F7FB637",
    x"3F7FB683",
    x"3F7FB6CF",
    x"3F7FB71B",
    x"3F7FB767",
    x"3F7FB7B2",
    x"3F7FB7FE",
    x"3F7FB849",
    x"3F7FB894",
    x"3F7FB8DF",
    x"3F7FB92A",
    x"3F7FB975",
    x"3F7FB9BF",
    x"3F7FBA0A",
    x"3F7FBA54",
    x"3F7FBA9E",
    x"3F7FBAE8",
    x"3F7FBB32",
    x"3F7FBB7B",
    x"3F7FBBC5",
    x"3F7FBC0E",
    x"3F7FBC57",
    x"3F7FBCA0",
    x"3F7FBCE9",
    x"3F7FBD32",
    x"3F7FBD7A",
    x"3F7FBDC2",
    x"3F7FBE0B",
    x"3F7FBE53",
    x"3F7FBE9B",
    x"3F7FBEE2",
    x"3F7FBF2A",
    x"3F7FBF72",
    x"3F7FBFB9",
    x"3F7FC000",
    x"3F7FC047",
    x"3F7FC08E",
    x"3F7FC0D4",
    x"3F7FC11B",
    x"3F7FC161",
    x"3F7FC1A8",
    x"3F7FC1EE",
    x"3F7FC234",
    x"3F7FC279",
    x"3F7FC2BF",
    x"3F7FC304",
    x"3F7FC34A",
    x"3F7FC38F",
    x"3F7FC3D4",
    x"3F7FC419",
    x"3F7FC45D",
    x"3F7FC4A2",
    x"3F7FC4E6",
    x"3F7FC52A",
    x"3F7FC56F",
    x"3F7FC5B2",
    x"3F7FC5F6",
    x"3F7FC63A",
    x"3F7FC67D",
    x"3F7FC6C1",
    x"3F7FC704",
    x"3F7FC747",
    x"3F7FC789",
    x"3F7FC7CC",
    x"3F7FC80F",
    x"3F7FC851",
    x"3F7FC893",
    x"3F7FC8D5",
    x"3F7FC917",
    x"3F7FC959",
    x"3F7FC99B",
    x"3F7FC9DC",
    x"3F7FCA1D",
    x"3F7FCA5E",
    x"3F7FCA9F",
    x"3F7FCAE0",
    x"3F7FCB21",
    x"3F7FCB61",
    x"3F7FCBA2",
    x"3F7FCBE2",
    x"3F7FCC22",
    x"3F7FCC62",
    x"3F7FCCA2",
    x"3F7FCCE1",
    x"3F7FCD21",
    x"3F7FCD60",
    x"3F7FCD9F",
    x"3F7FCDDE",
    x"3F7FCE1D",
    x"3F7FCE5C",
    x"3F7FCE9A",
    x"3F7FCED9",
    x"3F7FCF17",
    x"3F7FCF55",
    x"3F7FCF93",
    x"3F7FCFD1",
    x"3F7FD00E",
    x"3F7FD04C",
    x"3F7FD089",
    x"3F7FD0C6",
    x"3F7FD103",
    x"3F7FD140",
    x"3F7FD17C",
    x"3F7FD1B9",
    x"3F7FD1F5",
    x"3F7FD232",
    x"3F7FD26E",
    x"3F7FD2A9",
    x"3F7FD2E5",
    x"3F7FD321",
    x"3F7FD35C",
    x"3F7FD397",
    x"3F7FD3D3",
    x"3F7FD40E",
    x"3F7FD448",
    x"3F7FD483",
    x"3F7FD4BE",
    x"3F7FD4F8",
    x"3F7FD532",
    x"3F7FD56C",
    x"3F7FD5A6",
    x"3F7FD5E0",
    x"3F7FD619",
    x"3F7FD653",
    x"3F7FD68C",
    x"3F7FD6C5",
    x"3F7FD6FE",
    x"3F7FD737",
    x"3F7FD770",
    x"3F7FD7A8",
    x"3F7FD7E1",
    x"3F7FD819",
    x"3F7FD851",
    x"3F7FD889",
    x"3F7FD8C0",
    x"3F7FD8F8",
    x"3F7FD92F",
    x"3F7FD967",
    x"3F7FD99E",
    x"3F7FD9D5",
    x"3F7FDA0C",
    x"3F7FDA42",
    x"3F7FDA79",
    x"3F7FDAAF",
    x"3F7FDAE5",
    x"3F7FDB1B",
    x"3F7FDB51",
    x"3F7FDB87",
    x"3F7FDBBD",
    x"3F7FDBF2",
    x"3F7FDC27",
    x"3F7FDC5C",
    x"3F7FDC91",
    x"3F7FDCC6",
    x"3F7FDCFB",
    x"3F7FDD2F",
    x"3F7FDD64",
    x"3F7FDD98",
    x"3F7FDDCC",
    x"3F7FDE00",
    x"3F7FDE33",
    x"3F7FDE67",
    x"3F7FDE9A",
    x"3F7FDECE",
    x"3F7FDF01",
    x"3F7FDF34",
    x"3F7FDF67",
    x"3F7FDF99",
    x"3F7FDFCC",
    x"3F7FDFFE",
    x"3F7FE030",
    x"3F7FE062",
    x"3F7FE094",
    x"3F7FE0C6",
    x"3F7FE0F8",
    x"3F7FE129",
    x"3F7FE15A",
    x"3F7FE18B",
    x"3F7FE1BC",
    x"3F7FE1ED",
    x"3F7FE21E",
    x"3F7FE24E",
    x"3F7FE27F",
    x"3F7FE2AF",
    x"3F7FE2DF",
    x"3F7FE30F",
    x"3F7FE33E",
    x"3F7FE36E",
    x"3F7FE39D",
    x"3F7FE3CD",
    x"3F7FE3FC",
    x"3F7FE42B",
    x"3F7FE459",
    x"3F7FE488",
    x"3F7FE4B7",
    x"3F7FE4E5",
    x"3F7FE513",
    x"3F7FE541",
    x"3F7FE56F",
    x"3F7FE59D",
    x"3F7FE5CA",
    x"3F7FE5F8",
    x"3F7FE625",
    x"3F7FE652",
    x"3F7FE67F",
    x"3F7FE6AC",
    x"3F7FE6D8",
    x"3F7FE705",
    x"3F7FE731",
    x"3F7FE75D",
    x"3F7FE789",
    x"3F7FE7B5",
    x"3F7FE7E1",
    x"3F7FE80D",
    x"3F7FE838",
    x"3F7FE863",
    x"3F7FE88E",
    x"3F7FE8B9",
    x"3F7FE8E4",
    x"3F7FE90F",
    x"3F7FE939",
    x"3F7FE964",
    x"3F7FE98E",
    x"3F7FE9B8",
    x"3F7FE9E2",
    x"3F7FEA0B",
    x"3F7FEA35",
    x"3F7FEA5E",
    x"3F7FEA87",
    x"3F7FEAB1",
    x"3F7FEADA",
    x"3F7FEB02",
    x"3F7FEB2B",
    x"3F7FEB53",
    x"3F7FEB7C",
    x"3F7FEBA4",
    x"3F7FEBCC",
    x"3F7FEBF4",
    x"3F7FEC1B",
    x"3F7FEC43",
    x"3F7FEC6A",
    x"3F7FEC92",
    x"3F7FECB9",
    x"3F7FECE0",
    x"3F7FED06",
    x"3F7FED2D",
    x"3F7FED54",
    x"3F7FED7A",
    x"3F7FEDA0",
    x"3F7FEDC6",
    x"3F7FEDEC",
    x"3F7FEE12",
    x"3F7FEE37",
    x"3F7FEE5D",
    x"3F7FEE82",
    x"3F7FEEA7",
    x"3F7FEECC",
    x"3F7FEEF1",
    x"3F7FEF15",
    x"3F7FEF3A",
    x"3F7FEF5E",
    x"3F7FEF82",
    x"3F7FEFA6",
    x"3F7FEFCA",
    x"3F7FEFEE",
    x"3F7FF011",
    x"3F7FF035",
    x"3F7FF058",
    x"3F7FF07B",
    x"3F7FF09E",
    x"3F7FF0C1",
    x"3F7FF0E3",
    x"3F7FF106",
    x"3F7FF128",
    x"3F7FF14A",
    x"3F7FF16C",
    x"3F7FF18E",
    x"3F7FF1B0",
    x"3F7FF1D1",
    x"3F7FF1F3",
    x"3F7FF214",
    x"3F7FF235",
    x"3F7FF256",
    x"3F7FF277",
    x"3F7FF297",
    x"3F7FF2B8",
    x"3F7FF2D8",
    x"3F7FF2F8",
    x"3F7FF318",
    x"3F7FF338",
    x"3F7FF358",
    x"3F7FF377",
    x"3F7FF397",
    x"3F7FF3B6",
    x"3F7FF3D5",
    x"3F7FF3F4",
    x"3F7FF413",
    x"3F7FF431",
    x"3F7FF450",
    x"3F7FF46E",
    x"3F7FF48C",
    x"3F7FF4AA",
    x"3F7FF4C8",
    x"3F7FF4E6",
    x"3F7FF503",
    x"3F7FF521",
    x"3F7FF53E",
    x"3F7FF55B",
    x"3F7FF578",
    x"3F7FF595",
    x"3F7FF5B1",
    x"3F7FF5CE",
    x"3F7FF5EA",
    x"3F7FF606",
    x"3F7FF622",
    x"3F7FF63E",
    x"3F7FF659",
    x"3F7FF675",
    x"3F7FF690",
    x"3F7FF6AC",
    x"3F7FF6C7",
    x"3F7FF6E2",
    x"3F7FF6FC",
    x"3F7FF717",
    x"3F7FF731",
    x"3F7FF74C",
    x"3F7FF766",
    x"3F7FF780",
    x"3F7FF79A",
    x"3F7FF7B3",
    x"3F7FF7CD",
    x"3F7FF7E6",
    x"3F7FF7FF",
    x"3F7FF818",
    x"3F7FF831",
    x"3F7FF84A",
    x"3F7FF863",
    x"3F7FF87B",
    x"3F7FF893",
    x"3F7FF8AC",
    x"3F7FF8C4",
    x"3F7FF8DB",
    x"3F7FF8F3",
    x"3F7FF90B",
    x"3F7FF922",
    x"3F7FF939",
    x"3F7FF950",
    x"3F7FF967",
    x"3F7FF97E",
    x"3F7FF994",
    x"3F7FF9AB",
    x"3F7FF9C1",
    x"3F7FF9D7",
    x"3F7FF9ED",
    x"3F7FFA03",
    x"3F7FFA19",
    x"3F7FFA2E",
    x"3F7FFA44",
    x"3F7FFA59",
    x"3F7FFA6E",
    x"3F7FFA83",
    x"3F7FFA97",
    x"3F7FFAAC",
    x"3F7FFAC1",
    x"3F7FFAD5",
    x"3F7FFAE9",
    x"3F7FFAFD",
    x"3F7FFB11",
    x"3F7FFB24",
    x"3F7FFB38",
    x"3F7FFB4B",
    x"3F7FFB5E",
    x"3F7FFB71",
    x"3F7FFB84",
    x"3F7FFB97",
    x"3F7FFBAA",
    x"3F7FFBBC",
    x"3F7FFBCE",
    x"3F7FFBE1",
    x"3F7FFBF2",
    x"3F7FFC04",
    x"3F7FFC16",
    x"3F7FFC27",
    x"3F7FFC39",
    x"3F7FFC4A",
    x"3F7FFC5B",
    x"3F7FFC6C",
    x"3F7FFC7D",
    x"3F7FFC8D",
    x"3F7FFC9E",
    x"3F7FFCAE",
    x"3F7FFCBE",
    x"3F7FFCCE",
    x"3F7FFCDE",
    x"3F7FFCED",
    x"3F7FFCFD",
    x"3F7FFD0C",
    x"3F7FFD1B",
    x"3F7FFD2B",
    x"3F7FFD39",
    x"3F7FFD48",
    x"3F7FFD57",
    x"3F7FFD65",
    x"3F7FFD73",
    x"3F7FFD81",
    x"3F7FFD8F",
    x"3F7FFD9D",
    x"3F7FFDAB",
    x"3F7FFDB8",
    x"3F7FFDC6",
    x"3F7FFDD3",
    x"3F7FFDE0",
    x"3F7FFDED",
    x"3F7FFDFA",
    x"3F7FFE06",
    x"3F7FFE13",
    x"3F7FFE1F",
    x"3F7FFE2B",
    x"3F7FFE37",
    x"3F7FFE43",
    x"3F7FFE4E",
    x"3F7FFE5A",
    x"3F7FFE65",
    x"3F7FFE70",
    x"3F7FFE7B",
    x"3F7FFE86",
    x"3F7FFE91",
    x"3F7FFE9B",
    x"3F7FFEA6",
    x"3F7FFEB0",
    x"3F7FFEBA",
    x"3F7FFEC4",
    x"3F7FFECE",
    x"3F7FFED8",
    x"3F7FFEE1",
    x"3F7FFEEA",
    x"3F7FFEF4",
    x"3F7FFEFD",
    x"3F7FFF05",
    x"3F7FFF0E",
    x"3F7FFF17",
    x"3F7FFF1F",
    x"3F7FFF27",
    x"3F7FFF30",
    x"3F7FFF37",
    x"3F7FFF3F",
    x"3F7FFF47",
    x"3F7FFF4E",
    x"3F7FFF56",
    x"3F7FFF5D",
    x"3F7FFF64",
    x"3F7FFF6B",
    x"3F7FFF71",
    x"3F7FFF78",
    x"3F7FFF7E",
    x"3F7FFF85",
    x"3F7FFF8B",
    x"3F7FFF91",
    x"3F7FFF96",
    x"3F7FFF9C",
    x"3F7FFFA2",
    x"3F7FFFA7",
    x"3F7FFFAC",
    x"3F7FFFB1",
    x"3F7FFFB6",
    x"3F7FFFBB",
    x"3F7FFFBF",
    x"3F7FFFC4",
    x"3F7FFFC8",
    x"3F7FFFCC",
    x"3F7FFFD0",
    x"3F7FFFD4",
    x"3F7FFFD7",
    x"3F7FFFDB",
    x"3F7FFFDE",
    x"3F7FFFE1",
    x"3F7FFFE4",
    x"3F7FFFE7",
    x"3F7FFFEA",
    x"3F7FFFEC",
    x"3F7FFFEF",
    x"3F7FFFF1",
    x"3F7FFFF3",
    x"3F7FFFF5",
    x"3F7FFFF7",
    x"3F7FFFF8",
    x"3F7FFFFA",
    x"3F7FFFFB",
    x"3F7FFFFC",
    x"3F7FFFFD",
    x"3F7FFFFE",
    x"3F7FFFFF",
    x"3F7FFFFF",
    x"3F800000",
    x"3F800000",
    x"3F800000",
    x"3F800000",
    x"3F800000",
    x"3F7FFFFF",
    x"3F7FFFFF",
    x"3F7FFFFE",
    x"3F7FFFFD",
    x"3F7FFFFC",
    x"3F7FFFFB",
    x"3F7FFFFA",
    x"3F7FFFF8",
    x"3F7FFFF7",
    x"3F7FFFF5",
    x"3F7FFFF3",
    x"3F7FFFF1",
    x"3F7FFFEF",
    x"3F7FFFEC",
    x"3F7FFFEA",
    x"3F7FFFE7",
    x"3F7FFFE4",
    x"3F7FFFE1",
    x"3F7FFFDE",
    x"3F7FFFDB",
    x"3F7FFFD7",
    x"3F7FFFD4",
    x"3F7FFFD0",
    x"3F7FFFCC",
    x"3F7FFFC8",
    x"3F7FFFC4",
    x"3F7FFFBF",
    x"3F7FFFBB",
    x"3F7FFFB6",
    x"3F7FFFB1",
    x"3F7FFFAC",
    x"3F7FFFA7",
    x"3F7FFFA2",
    x"3F7FFF9C",
    x"3F7FFF96",
    x"3F7FFF91",
    x"3F7FFF8B",
    x"3F7FFF85",
    x"3F7FFF7E",
    x"3F7FFF78",
    x"3F7FFF71",
    x"3F7FFF6B",
    x"3F7FFF64",
    x"3F7FFF5D",
    x"3F7FFF56",
    x"3F7FFF4E",
    x"3F7FFF47",
    x"3F7FFF3F",
    x"3F7FFF37",
    x"3F7FFF30",
    x"3F7FFF27",
    x"3F7FFF1F",
    x"3F7FFF17",
    x"3F7FFF0E",
    x"3F7FFF05",
    x"3F7FFEFD",
    x"3F7FFEF4",
    x"3F7FFEEA",
    x"3F7FFEE1",
    x"3F7FFED8",
    x"3F7FFECE",
    x"3F7FFEC4",
    x"3F7FFEBA",
    x"3F7FFEB0",
    x"3F7FFEA6",
    x"3F7FFE9B",
    x"3F7FFE91",
    x"3F7FFE86",
    x"3F7FFE7B",
    x"3F7FFE70",
    x"3F7FFE65",
    x"3F7FFE5A",
    x"3F7FFE4E",
    x"3F7FFE43",
    x"3F7FFE37",
    x"3F7FFE2B",
    x"3F7FFE1F",
    x"3F7FFE13",
    x"3F7FFE06",
    x"3F7FFDFA",
    x"3F7FFDED",
    x"3F7FFDE0",
    x"3F7FFDD3",
    x"3F7FFDC6",
    x"3F7FFDB8",
    x"3F7FFDAB",
    x"3F7FFD9D",
    x"3F7FFD8F",
    x"3F7FFD81",
    x"3F7FFD73",
    x"3F7FFD65",
    x"3F7FFD57",
    x"3F7FFD48",
    x"3F7FFD39",
    x"3F7FFD2B",
    x"3F7FFD1B",
    x"3F7FFD0C",
    x"3F7FFCFD",
    x"3F7FFCED",
    x"3F7FFCDE",
    x"3F7FFCCE",
    x"3F7FFCBE",
    x"3F7FFCAE",
    x"3F7FFC9E",
    x"3F7FFC8D",
    x"3F7FFC7D",
    x"3F7FFC6C",
    x"3F7FFC5B",
    x"3F7FFC4A",
    x"3F7FFC39",
    x"3F7FFC27",
    x"3F7FFC16",
    x"3F7FFC04",
    x"3F7FFBF2",
    x"3F7FFBE1",
    x"3F7FFBCE",
    x"3F7FFBBC",
    x"3F7FFBAA",
    x"3F7FFB97",
    x"3F7FFB84",
    x"3F7FFB71",
    x"3F7FFB5E",
    x"3F7FFB4B",
    x"3F7FFB38",
    x"3F7FFB24",
    x"3F7FFB11",
    x"3F7FFAFD",
    x"3F7FFAE9",
    x"3F7FFAD5",
    x"3F7FFAC1",
    x"3F7FFAAC",
    x"3F7FFA97",
    x"3F7FFA83",
    x"3F7FFA6E",
    x"3F7FFA59",
    x"3F7FFA44",
    x"3F7FFA2E",
    x"3F7FFA19",
    x"3F7FFA03",
    x"3F7FF9ED",
    x"3F7FF9D7",
    x"3F7FF9C1",
    x"3F7FF9AB",
    x"3F7FF994",
    x"3F7FF97E",
    x"3F7FF967",
    x"3F7FF950",
    x"3F7FF939",
    x"3F7FF922",
    x"3F7FF90B",
    x"3F7FF8F3",
    x"3F7FF8DB",
    x"3F7FF8C4",
    x"3F7FF8AC",
    x"3F7FF893",
    x"3F7FF87B",
    x"3F7FF863",
    x"3F7FF84A",
    x"3F7FF831",
    x"3F7FF818",
    x"3F7FF7FF",
    x"3F7FF7E6",
    x"3F7FF7CD",
    x"3F7FF7B3",
    x"3F7FF79A",
    x"3F7FF780",
    x"3F7FF766",
    x"3F7FF74C",
    x"3F7FF731",
    x"3F7FF717",
    x"3F7FF6FC",
    x"3F7FF6E2",
    x"3F7FF6C7",
    x"3F7FF6AC",
    x"3F7FF690",
    x"3F7FF675",
    x"3F7FF659",
    x"3F7FF63E",
    x"3F7FF622",
    x"3F7FF606",
    x"3F7FF5EA",
    x"3F7FF5CE",
    x"3F7FF5B1",
    x"3F7FF595",
    x"3F7FF578",
    x"3F7FF55B",
    x"3F7FF53E",
    x"3F7FF521",
    x"3F7FF503",
    x"3F7FF4E6",
    x"3F7FF4C8",
    x"3F7FF4AA",
    x"3F7FF48C",
    x"3F7FF46E",
    x"3F7FF450",
    x"3F7FF431",
    x"3F7FF413",
    x"3F7FF3F4",
    x"3F7FF3D5",
    x"3F7FF3B6",
    x"3F7FF397",
    x"3F7FF377",
    x"3F7FF358",
    x"3F7FF338",
    x"3F7FF318",
    x"3F7FF2F8",
    x"3F7FF2D8",
    x"3F7FF2B8",
    x"3F7FF297",
    x"3F7FF277",
    x"3F7FF256",
    x"3F7FF235",
    x"3F7FF214",
    x"3F7FF1F3",
    x"3F7FF1D1",
    x"3F7FF1B0",
    x"3F7FF18E",
    x"3F7FF16C",
    x"3F7FF14A",
    x"3F7FF128",
    x"3F7FF106",
    x"3F7FF0E3",
    x"3F7FF0C1",
    x"3F7FF09E",
    x"3F7FF07B",
    x"3F7FF058",
    x"3F7FF035",
    x"3F7FF011",
    x"3F7FEFEE",
    x"3F7FEFCA",
    x"3F7FEFA6",
    x"3F7FEF82",
    x"3F7FEF5E",
    x"3F7FEF3A",
    x"3F7FEF15",
    x"3F7FEEF1",
    x"3F7FEECC",
    x"3F7FEEA7",
    x"3F7FEE82",
    x"3F7FEE5D",
    x"3F7FEE37",
    x"3F7FEE12",
    x"3F7FEDEC",
    x"3F7FEDC6",
    x"3F7FEDA0",
    x"3F7FED7A",
    x"3F7FED54",
    x"3F7FED2D",
    x"3F7FED06",
    x"3F7FECE0",
    x"3F7FECB9",
    x"3F7FEC92",
    x"3F7FEC6A",
    x"3F7FEC43",
    x"3F7FEC1B",
    x"3F7FEBF4",
    x"3F7FEBCC",
    x"3F7FEBA4",
    x"3F7FEB7C",
    x"3F7FEB53",
    x"3F7FEB2B",
    x"3F7FEB02",
    x"3F7FEADA",
    x"3F7FEAB1",
    x"3F7FEA87",
    x"3F7FEA5E",
    x"3F7FEA35",
    x"3F7FEA0B",
    x"3F7FE9E2",
    x"3F7FE9B8",
    x"3F7FE98E",
    x"3F7FE964",
    x"3F7FE939",
    x"3F7FE90F",
    x"3F7FE8E4",
    x"3F7FE8B9",
    x"3F7FE88E",
    x"3F7FE863",
    x"3F7FE838",
    x"3F7FE80D",
    x"3F7FE7E1",
    x"3F7FE7B5",
    x"3F7FE789",
    x"3F7FE75D",
    x"3F7FE731",
    x"3F7FE705",
    x"3F7FE6D8",
    x"3F7FE6AC",
    x"3F7FE67F",
    x"3F7FE652",
    x"3F7FE625",
    x"3F7FE5F8",
    x"3F7FE5CA",
    x"3F7FE59D",
    x"3F7FE56F",
    x"3F7FE541",
    x"3F7FE513",
    x"3F7FE4E5",
    x"3F7FE4B7",
    x"3F7FE488",
    x"3F7FE459",
    x"3F7FE42B",
    x"3F7FE3FC",
    x"3F7FE3CD",
    x"3F7FE39D",
    x"3F7FE36E",
    x"3F7FE33E",
    x"3F7FE30F",
    x"3F7FE2DF",
    x"3F7FE2AF",
    x"3F7FE27F",
    x"3F7FE24E",
    x"3F7FE21E",
    x"3F7FE1ED",
    x"3F7FE1BC",
    x"3F7FE18B",
    x"3F7FE15A",
    x"3F7FE129",
    x"3F7FE0F8",
    x"3F7FE0C6",
    x"3F7FE094",
    x"3F7FE062",
    x"3F7FE030",
    x"3F7FDFFE",
    x"3F7FDFCC",
    x"3F7FDF99",
    x"3F7FDF67",
    x"3F7FDF34",
    x"3F7FDF01",
    x"3F7FDECE",
    x"3F7FDE9A",
    x"3F7FDE67",
    x"3F7FDE33",
    x"3F7FDE00",
    x"3F7FDDCC",
    x"3F7FDD98",
    x"3F7FDD64",
    x"3F7FDD2F",
    x"3F7FDCFB",
    x"3F7FDCC6",
    x"3F7FDC91",
    x"3F7FDC5C",
    x"3F7FDC27",
    x"3F7FDBF2",
    x"3F7FDBBD",
    x"3F7FDB87",
    x"3F7FDB51",
    x"3F7FDB1B",
    x"3F7FDAE5",
    x"3F7FDAAF",
    x"3F7FDA79",
    x"3F7FDA42",
    x"3F7FDA0C",
    x"3F7FD9D5",
    x"3F7FD99E",
    x"3F7FD967",
    x"3F7FD92F",
    x"3F7FD8F8",
    x"3F7FD8C0",
    x"3F7FD889",
    x"3F7FD851",
    x"3F7FD819",
    x"3F7FD7E1",
    x"3F7FD7A8",
    x"3F7FD770",
    x"3F7FD737",
    x"3F7FD6FE",
    x"3F7FD6C5",
    x"3F7FD68C",
    x"3F7FD653",
    x"3F7FD619",
    x"3F7FD5E0",
    x"3F7FD5A6",
    x"3F7FD56C",
    x"3F7FD532",
    x"3F7FD4F8",
    x"3F7FD4BE",
    x"3F7FD483",
    x"3F7FD448",
    x"3F7FD40E",
    x"3F7FD3D3",
    x"3F7FD397",
    x"3F7FD35C",
    x"3F7FD321",
    x"3F7FD2E5",
    x"3F7FD2A9",
    x"3F7FD26E",
    x"3F7FD232",
    x"3F7FD1F5",
    x"3F7FD1B9",
    x"3F7FD17C",
    x"3F7FD140",
    x"3F7FD103",
    x"3F7FD0C6",
    x"3F7FD089",
    x"3F7FD04C",
    x"3F7FD00E",
    x"3F7FCFD1",
    x"3F7FCF93",
    x"3F7FCF55",
    x"3F7FCF17",
    x"3F7FCED9",
    x"3F7FCE9A",
    x"3F7FCE5C",
    x"3F7FCE1D",
    x"3F7FCDDE",
    x"3F7FCD9F",
    x"3F7FCD60",
    x"3F7FCD21",
    x"3F7FCCE1",
    x"3F7FCCA2",
    x"3F7FCC62",
    x"3F7FCC22",
    x"3F7FCBE2",
    x"3F7FCBA2",
    x"3F7FCB61",
    x"3F7FCB21",
    x"3F7FCAE0",
    x"3F7FCA9F",
    x"3F7FCA5E",
    x"3F7FCA1D",
    x"3F7FC9DC",
    x"3F7FC99B",
    x"3F7FC959",
    x"3F7FC917",
    x"3F7FC8D5",
    x"3F7FC893",
    x"3F7FC851",
    x"3F7FC80F",
    x"3F7FC7CC",
    x"3F7FC789",
    x"3F7FC747",
    x"3F7FC704",
    x"3F7FC6C1",
    x"3F7FC67D",
    x"3F7FC63A",
    x"3F7FC5F6",
    x"3F7FC5B2",
    x"3F7FC56F",
    x"3F7FC52A",
    x"3F7FC4E6",
    x"3F7FC4A2",
    x"3F7FC45D",
    x"3F7FC419",
    x"3F7FC3D4",
    x"3F7FC38F",
    x"3F7FC34A",
    x"3F7FC304",
    x"3F7FC2BF",
    x"3F7FC279",
    x"3F7FC234",
    x"3F7FC1EE",
    x"3F7FC1A8",
    x"3F7FC161",
    x"3F7FC11B",
    x"3F7FC0D4",
    x"3F7FC08E",
    x"3F7FC047",
    x"3F7FC000",
    x"3F7FBFB9",
    x"3F7FBF72",
    x"3F7FBF2A",
    x"3F7FBEE2",
    x"3F7FBE9B",
    x"3F7FBE53",
    x"3F7FBE0B",
    x"3F7FBDC2",
    x"3F7FBD7A",
    x"3F7FBD32",
    x"3F7FBCE9",
    x"3F7FBCA0",
    x"3F7FBC57",
    x"3F7FBC0E",
    x"3F7FBBC5",
    x"3F7FBB7B",
    x"3F7FBB32",
    x"3F7FBAE8",
    x"3F7FBA9E",
    x"3F7FBA54",
    x"3F7FBA0A",
    x"3F7FB9BF",
    x"3F7FB975",
    x"3F7FB92A",
    x"3F7FB8DF",
    x"3F7FB894",
    x"3F7FB849",
    x"3F7FB7FE",
    x"3F7FB7B2",
    x"3F7FB767",
    x"3F7FB71B",
    x"3F7FB6CF",
    x"3F7FB683",
    x"3F7FB637",
    x"3F7FB5EA",
    x"3F7FB59E",
    x"3F7FB551",
    x"3F7FB504",
    x"3F7FB4B7",
    x"3F7FB46A",
    x"3F7FB41D",
    x"3F7FB3CF",
    x"3F7FB382",
    x"3F7FB334",
    x"3F7FB2E6",
    x"3F7FB298",
    x"3F7FB24A",
    x"3F7FB1FB",
    x"3F7FB1AD",
    x"3F7FB15E",
    x"3F7FB10F",
    x"3F7FB0C0",
    x"3F7FB071",
    x"3F7FB022",
    x"3F7FAFD2",
    x"3F7FAF83",
    x"3F7FAF33",
    x"3F7FAEE3",
    x"3F7FAE93",
    x"3F7FAE43",
    x"3F7FADF2",
    x"3F7FADA2",
    x"3F7FAD51",
    x"3F7FAD00",
    x"3F7FACAF",
    x"3F7FAC5E",
    x"3F7FAC0D",
    x"3F7FABBB",
    x"3F7FAB6A",
    x"3F7FAB18",
    x"3F7FAAC6",
    x"3F7FAA74",
    x"3F7FAA21",
    x"3F7FA9CF",
    x"3F7FA97D",
    x"3F7FA92A",
    x"3F7FA8D7",
    x"3F7FA884",
    x"3F7FA831",
    x"3F7FA7DE",
    x"3F7FA78A",
    x"3F7FA736",
    x"3F7FA6E3",
    x"3F7FA68F",
    x"3F7FA63B",
    x"3F7FA5E6",
    x"3F7FA592",
    x"3F7FA53D",
    x"3F7FA4E9",
    x"3F7FA494",
    x"3F7FA43F",
    x"3F7FA3EA",
    x"3F7FA394",
    x"3F7FA33F",
    x"3F7FA2E9",
    x"3F7FA294",
    x"3F7FA23E",
    x"3F7FA1E8",
    x"3F7FA191",
    x"3F7FA13B",
    x"3F7FA0E4",
    x"3F7FA08E",
    x"3F7FA037",
    x"3F7F9FE0",
    x"3F7F9F89",
    x"3F7F9F31",
    x"3F7F9EDA",
    x"3F7F9E82",
    x"3F7F9E2A",
    x"3F7F9DD2",
    x"3F7F9D7A",
    x"3F7F9D22",
    x"3F7F9CCA",
    x"3F7F9C71",
    x"3F7F9C18",
    x"3F7F9BC0",
    x"3F7F9B67",
    x"3F7F9B0D",
    x"3F7F9AB4",
    x"3F7F9A5B",
    x"3F7F9A01",
    x"3F7F99A7",
    x"3F7F994D",
    x"3F7F98F3",
    x"3F7F9899",
    x"3F7F983F",
    x"3F7F97E4",
    x"3F7F9789",
    x"3F7F972E",
    x"3F7F96D3",
    x"3F7F9678",
    x"3F7F961D",
    x"3F7F95C1",
    x"3F7F9566",
    x"3F7F950A",
    x"3F7F94AE",
    x"3F7F9452",
    x"3F7F93F6",
    x"3F7F9399",
    x"3F7F933D",
    x"3F7F92E0",
    x"3F7F9283",
    x"3F7F9226",
    x"3F7F91C9",
    x"3F7F916C",
    x"3F7F910E",
    x"3F7F90B1",
    x"3F7F9053",
    x"3F7F8FF5",
    x"3F7F8F97",
    x"3F7F8F39",
    x"3F7F8EDA",
    x"3F7F8E7C",
    x"3F7F8E1D",
    x"3F7F8DBE",
    x"3F7F8D5F",
    x"3F7F8D00",
    x"3F7F8CA1",
    x"3F7F8C41",
    x"3F7F8BE1",
    x"3F7F8B82",
    x"3F7F8B22",
    x"3F7F8AC2",
    x"3F7F8A61",
    x"3F7F8A01",
    x"3F7F89A0",
    x"3F7F8940",
    x"3F7F88DF",
    x"3F7F887E",
    x"3F7F881D",
    x"3F7F87BB",
    x"3F7F875A",
    x"3F7F86F8",
    x"3F7F8696",
    x"3F7F8634",
    x"3F7F85D2",
    x"3F7F8570",
    x"3F7F850E",
    x"3F7F84AB",
    x"3F7F8448",
    x"3F7F83E6",
    x"3F7F8383",
    x"3F7F831F",
    x"3F7F82BC",
    x"3F7F8259",
    x"3F7F81F5",
    x"3F7F8191",
    x"3F7F812D",
    x"3F7F80C9",
    x"3F7F8065",
    x"3F7F8000",
    x"3F7F7F9C",
    x"3F7F7F37",
    x"3F7F7ED2",
    x"3F7F7E6D",
    x"3F7F7E08",
    x"3F7F7DA3",
    x"3F7F7D3D",
    x"3F7F7CD8",
    x"3F7F7C72",
    x"3F7F7C0C",
    x"3F7F7BA6",
    x"3F7F7B40",
    x"3F7F7AD9",
    x"3F7F7A73",
    x"3F7F7A0C",
    x"3F7F79A5",
    x"3F7F793E",
    x"3F7F78D7",
    x"3F7F7870",
    x"3F7F7808",
    x"3F7F77A0",
    x"3F7F7739",
    x"3F7F76D1",
    x"3F7F7669",
    x"3F7F7600",
    x"3F7F7598",
    x"3F7F752F",
    x"3F7F74C7",
    x"3F7F745E",
    x"3F7F73F5",
    x"3F7F738C",
    x"3F7F7322",
    x"3F7F72B9",
    x"3F7F724F",
    x"3F7F71E5",
    x"3F7F717B",
    x"3F7F7111",
    x"3F7F70A7",
    x"3F7F703D",
    x"3F7F6FD2",
    x"3F7F6F67",
    x"3F7F6EFD",
    x"3F7F6E92",
    x"3F7F6E26",
    x"3F7F6DBB",
    x"3F7F6D50",
    x"3F7F6CE4",
    x"3F7F6C78",
    x"3F7F6C0C",
    x"3F7F6BA0",
    x"3F7F6B34",
    x"3F7F6AC7",
    x"3F7F6A5B",
    x"3F7F69EE",
    x"3F7F6981",
    x"3F7F6914",
    x"3F7F68A7",
    x"3F7F683A",
    x"3F7F67CC",
    x"3F7F675F",
    x"3F7F66F1",
    x"3F7F6683",
    x"3F7F6615",
    x"3F7F65A7",
    x"3F7F6538",
    x"3F7F64CA",
    x"3F7F645B",
    x"3F7F63EC",
    x"3F7F637D",
    x"3F7F630E",
    x"3F7F629E",
    x"3F7F622F",
    x"3F7F61BF",
    x"3F7F6150",
    x"3F7F60E0",
    x"3F7F606F",
    x"3F7F5FFF",
    x"3F7F5F8F",
    x"3F7F5F1E",
    x"3F7F5EAE",
    x"3F7F5E3D",
    x"3F7F5DCC",
    x"3F7F5D5A",
    x"3F7F5CE9",
    x"3F7F5C78",
    x"3F7F5C06",
    x"3F7F5B94",
    x"3F7F5B22",
    x"3F7F5AB0",
    x"3F7F5A3E",
    x"3F7F59CC",
    x"3F7F5959",
    x"3F7F58E6",
    x"3F7F5873",
    x"3F7F5800",
    x"3F7F578D",
    x"3F7F571A",
    x"3F7F56A6",
    x"3F7F5633",
    x"3F7F55BF",
    x"3F7F554B",
    x"3F7F54D7",
    x"3F7F5463",
    x"3F7F53EE",
    x"3F7F537A",
    x"3F7F5305",
    x"3F7F5290",
    x"3F7F521B",
    x"3F7F51A6",
    x"3F7F5131",
    x"3F7F50BB",
    x"3F7F5045",
    x"3F7F4FD0",
    x"3F7F4F5A",
    x"3F7F4EE4",
    x"3F7F4E6D",
    x"3F7F4DF7",
    x"3F7F4D80",
    x"3F7F4D0A",
    x"3F7F4C93",
    x"3F7F4C1C",
    x"3F7F4BA5",
    x"3F7F4B2D",
    x"3F7F4AB6",
    x"3F7F4A3E",
    x"3F7F49C6",
    x"3F7F494E",
    x"3F7F48D6",
    x"3F7F485E",
    x"3F7F47E6",
    x"3F7F476D",
    x"3F7F46F4",
    x"3F7F467C",
    x"3F7F4603",
    x"3F7F4589",
    x"3F7F4510",
    x"3F7F4497",
    x"3F7F441D",
    x"3F7F43A3",
    x"3F7F4329",
    x"3F7F42AF",
    x"3F7F4235",
    x"3F7F41BA",
    x"3F7F4140",
    x"3F7F40C5",
    x"3F7F404A",
    x"3F7F3FCF",
    x"3F7F3F54",
    x"3F7F3ED9",
    x"3F7F3E5D",
    x"3F7F3DE2",
    x"3F7F3D66",
    x"3F7F3CEA",
    x"3F7F3C6E",
    x"3F7F3BF2",
    x"3F7F3B75",
    x"3F7F3AF9",
    x"3F7F3A7C",
    x"3F7F39FF",
    x"3F7F3982",
    x"3F7F3905",
    x"3F7F3888",
    x"3F7F380A",
    x"3F7F378C",
    x"3F7F370F",
    x"3F7F3691",
    x"3F7F3613",
    x"3F7F3594",
    x"3F7F3516",
    x"3F7F3497",
    x"3F7F3419",
    x"3F7F339A",
    x"3F7F331B",
    x"3F7F329C",
    x"3F7F321C",
    x"3F7F319D",
    x"3F7F311D",
    x"3F7F309E",
    x"3F7F301E",
    x"3F7F2F9D",
    x"3F7F2F1D",
    x"3F7F2E9D",
    x"3F7F2E1C",
    x"3F7F2D9C",
    x"3F7F2D1B",
    x"3F7F2C9A",
    x"3F7F2C19",
    x"3F7F2B97",
    x"3F7F2B16",
    x"3F7F2A94",
    x"3F7F2A12",
    x"3F7F2990",
    x"3F7F290E",
    x"3F7F288C",
    x"3F7F280A",
    x"3F7F2787",
    x"3F7F2704",
    x"3F7F2682",
    x"3F7F25FF",
    x"3F7F257B",
    x"3F7F24F8",
    x"3F7F2475",
    x"3F7F23F1",
    x"3F7F236D",
    x"3F7F22E9",
    x"3F7F2265",
    x"3F7F21E1",
    x"3F7F215C",
    x"3F7F20D8",
    x"3F7F2053",
    x"3F7F1FCE",
    x"3F7F1F49",
    x"3F7F1EC4",
    x"3F7F1E3F",
    x"3F7F1DB9",
    x"3F7F1D34",
    x"3F7F1CAE",
    x"3F7F1C28",
    x"3F7F1BA2",
    x"3F7F1B1C",
    x"3F7F1A95",
    x"3F7F1A0F",
    x"3F7F1988",
    x"3F7F1901",
    x"3F7F187A",
    x"3F7F17F3",
    x"3F7F176C",
    x"3F7F16E4",
    x"3F7F165D",
    x"3F7F15D5",
    x"3F7F154D",
    x"3F7F14C5",
    x"3F7F143D",
    x"3F7F13B4",
    x"3F7F132C",
    x"3F7F12A3",
    x"3F7F121A",
    x"3F7F1191",
    x"3F7F1108",
    x"3F7F107F",
    x"3F7F0FF5",
    x"3F7F0F6C",
    x"3F7F0EE2",
    x"3F7F0E58",
    x"3F7F0DCE",
    x"3F7F0D44",
    x"3F7F0CB9",
    x"3F7F0C2F",
    x"3F7F0BA4",
    x"3F7F0B19",
    x"3F7F0A8E",
    x"3F7F0A03",
    x"3F7F0978",
    x"3F7F08EC",
    x"3F7F0861",
    x"3F7F07D5",
    x"3F7F0749",
    x"3F7F06BD",
    x"3F7F0631",
    x"3F7F05A4",
    x"3F7F0518",
    x"3F7F048B",
    x"3F7F03FE",
    x"3F7F0371",
    x"3F7F02E4",
    x"3F7F0257",
    x"3F7F01C9",
    x"3F7F013C",
    x"3F7F00AE",
    x"3F7F0020",
    x"3F7EFF92",
    x"3F7EFF04",
    x"3F7EFE75",
    x"3F7EFDE7",
    x"3F7EFD58",
    x"3F7EFCC9",
    x"3F7EFC3A",
    x"3F7EFBAB",
    x"3F7EFB1C",
    x"3F7EFA8C",
    x"3F7EF9FD",
    x"3F7EF96D",
    x"3F7EF8DD",
    x"3F7EF84D",
    x"3F7EF7BD",
    x"3F7EF72C",
    x"3F7EF69C",
    x"3F7EF60B",
    x"3F7EF57A",
    x"3F7EF4E9",
    x"3F7EF458",
    x"3F7EF3C7",
    x"3F7EF335",
    x"3F7EF2A4",
    x"3F7EF212",
    x"3F7EF180",
    x"3F7EF0EE",
    x"3F7EF05C",
    x"3F7EEFC9",
    x"3F7EEF37",
    x"3F7EEEA4",
    x"3F7EEE11",
    x"3F7EED7E",
    x"3F7EECEB",
    x"3F7EEC58",
    x"3F7EEBC4",
    x"3F7EEB31",
    x"3F7EEA9D",
    x"3F7EEA09",
    x"3F7EE975",
    x"3F7EE8E1",
    x"3F7EE84C",
    x"3F7EE7B8",
    x"3F7EE723",
    x"3F7EE68E",
    x"3F7EE5F9",
    x"3F7EE564",
    x"3F7EE4CF",
    x"3F7EE43A",
    x"3F7EE3A4",
    x"3F7EE30E",
    x"3F7EE278",
    x"3F7EE1E2",
    x"3F7EE14C",
    x"3F7EE0B6",
    x"3F7EE01F",
    x"3F7EDF88",
    x"3F7EDEF2",
    x"3F7EDE5B",
    x"3F7EDDC3",
    x"3F7EDD2C",
    x"3F7EDC95",
    x"3F7EDBFD",
    x"3F7EDB65",
    x"3F7EDACD",
    x"3F7EDA35",
    x"3F7ED99D",
    x"3F7ED905",
    x"3F7ED86C",
    x"3F7ED7D4",
    x"3F7ED73B",
    x"3F7ED6A2",
    x"3F7ED609",
    x"3F7ED56F",
    x"3F7ED4D6",
    x"3F7ED43C",
    x"3F7ED3A3",
    x"3F7ED309",
    x"3F7ED26F",
    x"3F7ED1D4",
    x"3F7ED13A",
    x"3F7ED0A0",
    x"3F7ED005",
    x"3F7ECF6A",
    x"3F7ECECF",
    x"3F7ECE34",
    x"3F7ECD99",
    x"3F7ECCFD",
    x"3F7ECC62",
    x"3F7ECBC6",
    x"3F7ECB2A",
    x"3F7ECA8E",
    x"3F7EC9F2",
    x"3F7EC955",
    x"3F7EC8B9",
    x"3F7EC81C",
    x"3F7EC780",
    x"3F7EC6E3",
    x"3F7EC645",
    x"3F7EC5A8",
    x"3F7EC50B",
    x"3F7EC46D",
    x"3F7EC3CF",
    x"3F7EC331",
    x"3F7EC293",
    x"3F7EC1F5",
    x"3F7EC157",
    x"3F7EC0B8",
    x"3F7EC01A",
    x"3F7EBF7B",
    x"3F7EBEDC",
    x"3F7EBE3D",
    x"3F7EBD9E",
    x"3F7EBCFE",
    x"3F7EBC5F",
    x"3F7EBBBF",
    x"3F7EBB1F",
    x"3F7EBA7F",
    x"3F7EB9DF",
    x"3F7EB93E",
    x"3F7EB89E",
    x"3F7EB7FD",
    x"3F7EB75C",
    x"3F7EB6BB",
    x"3F7EB61A",
    x"3F7EB579",
    x"3F7EB4D8",
    x"3F7EB436",
    x"3F7EB394",
    x"3F7EB2F2",
    x"3F7EB250",
    x"3F7EB1AE",
    x"3F7EB10C",
    x"3F7EB069",
    x"3F7EAFC7",
    x"3F7EAF24",
    x"3F7EAE81",
    x"3F7EADDE",
    x"3F7EAD3B",
    x"3F7EAC97",
    x"3F7EABF4",
    x"3F7EAB50",
    x"3F7EAAAC",
    x"3F7EAA08",
    x"3F7EA964",
    x"3F7EA8C0",
    x"3F7EA81B",
    x"3F7EA776",
    x"3F7EA6D2",
    x"3F7EA62D",
    x"3F7EA588",
    x"3F7EA4E2",
    x"3F7EA43D",
    x"3F7EA397",
    x"3F7EA2F2",
    x"3F7EA24C",
    x"3F7EA1A6",
    x"3F7EA100",
    x"3F7EA059",
    x"3F7E9FB3",
    x"3F7E9F0C",
    x"3F7E9E65",
    x"3F7E9DBE",
    x"3F7E9D17",
    x"3F7E9C70",
    x"3F7E9BC9",
    x"3F7E9B21",
    x"3F7E9A79",
    x"3F7E99D2",
    x"3F7E9929",
    x"3F7E9881",
    x"3F7E97D9",
    x"3F7E9731",
    x"3F7E9688",
    x"3F7E95DF",
    x"3F7E9536",
    x"3F7E948D",
    x"3F7E93E4",
    x"3F7E933A",
    x"3F7E9291",
    x"3F7E91E7",
    x"3F7E913D",
    x"3F7E9093",
    x"3F7E8FE9",
    x"3F7E8F3F",
    x"3F7E8E94",
    x"3F7E8DEA",
    x"3F7E8D3F",
    x"3F7E8C94",
    x"3F7E8BE9",
    x"3F7E8B3E",
    x"3F7E8A92",
    x"3F7E89E7",
    x"3F7E893B",
    x"3F7E888F",
    x"3F7E87E3",
    x"3F7E8737",
    x"3F7E868B",
    x"3F7E85DE",
    x"3F7E8532",
    x"3F7E8485",
    x"3F7E83D8",
    x"3F7E832B",
    x"3F7E827E",
    x"3F7E81D0",
    x"3F7E8123",
    x"3F7E8075",
    x"3F7E7FC7",
    x"3F7E7F19",
    x"3F7E7E6B",
    x"3F7E7DBD",
    x"3F7E7D0E",
    x"3F7E7C60",
    x"3F7E7BB1",
    x"3F7E7B02",
    x"3F7E7A53",
    x"3F7E79A4",
    x"3F7E78F4",
    x"3F7E7845",
    x"3F7E7795",
    x"3F7E76E5",
    x"3F7E7635",
    x"3F7E7585",
    x"3F7E74D5",
    x"3F7E7424",
    x"3F7E7374",
    x"3F7E72C3",
    x"3F7E7212",
    x"3F7E7161",
    x"3F7E70B0",
    x"3F7E6FFF",
    x"3F7E6F4D",
    x"3F7E6E9B",
    x"3F7E6DEA",
    x"3F7E6D38",
    x"3F7E6C85",
    x"3F7E6BD3",
    x"3F7E6B21",
    x"3F7E6A6E",
    x"3F7E69BB",
    x"3F7E6908",
    x"3F7E6855",
    x"3F7E67A2",
    x"3F7E66EF",
    x"3F7E663B",
    x"3F7E6588",
    x"3F7E64D4",
    x"3F7E6420",
    x"3F7E636C",
    x"3F7E62B7",
    x"3F7E6203",
    x"3F7E614E",
    x"3F7E609A",
    x"3F7E5FE5",
    x"3F7E5F30",
    x"3F7E5E7B",
    x"3F7E5DC5",
    x"3F7E5D10",
    x"3F7E5C5A",
    x"3F7E5BA4",
    x"3F7E5AEE",
    x"3F7E5A38",
    x"3F7E5982",
    x"3F7E58CB",
    x"3F7E5815",
    x"3F7E575E",
    x"3F7E56A7",
    x"3F7E55F0",
    x"3F7E5539",
    x"3F7E5482",
    x"3F7E53CA",
    x"3F7E5312",
    x"3F7E525B",
    x"3F7E51A3",
    x"3F7E50EB",
    x"3F7E5032",
    x"3F7E4F7A",
    x"3F7E4EC1",
    x"3F7E4E09",
    x"3F7E4D50",
    x"3F7E4C97",
    x"3F7E4BDE",
    x"3F7E4B24",
    x"3F7E4A6B",
    x"3F7E49B1",
    x"3F7E48F7",
    x"3F7E483D",
    x"3F7E4783",
    x"3F7E46C9",
    x"3F7E460F",
    x"3F7E4554",
    x"3F7E4499",
    x"3F7E43DE",
    x"3F7E4323",
    x"3F7E4268",
    x"3F7E41AD",
    x"3F7E40F1",
    x"3F7E4036",
    x"3F7E3F7A",
    x"3F7E3EBE",
    x"3F7E3E02",
    x"3F7E3D46",
    x"3F7E3C89",
    x"3F7E3BCD",
    x"3F7E3B10",
    x"3F7E3A53",
    x"3F7E3996",
    x"3F7E38D9",
    x"3F7E381C",
    x"3F7E375E",
    x"3F7E36A1",
    x"3F7E35E3",
    x"3F7E3525",
    x"3F7E3467",
    x"3F7E33A9",
    x"3F7E32EA",
    x"3F7E322C",
    x"3F7E316D",
    x"3F7E30AE",
    x"3F7E2FEF",
    x"3F7E2F30",
    x"3F7E2E71",
    x"3F7E2DB1",
    x"3F7E2CF2",
    x"3F7E2C32",
    x"3F7E2B72",
    x"3F7E2AB2",
    x"3F7E29F2",
    x"3F7E2931",
    x"3F7E2871",
    x"3F7E27B0",
    x"3F7E26EF",
    x"3F7E262E",
    x"3F7E256D",
    x"3F7E24AC",
    x"3F7E23EA",
    x"3F7E2329",
    x"3F7E2267",
    x"3F7E21A5",
    x"3F7E20E3",
    x"3F7E2021",
    x"3F7E1F5E",
    x"3F7E1E9C",
    x"3F7E1DD9",
    x"3F7E1D16",
    x"3F7E1C53",
    x"3F7E1B90",
    x"3F7E1ACD",
    x"3F7E1A09",
    x"3F7E1946",
    x"3F7E1882",
    x"3F7E17BE",
    x"3F7E16FA",
    x"3F7E1636",
    x"3F7E1572",
    x"3F7E14AD",
    x"3F7E13E8",
    x"3F7E1324",
    x"3F7E125F",
    x"3F7E1199",
    x"3F7E10D4",
    x"3F7E100F",
    x"3F7E0F49",
    x"3F7E0E83",
    x"3F7E0DBD",
    x"3F7E0CF7",
    x"3F7E0C31",
    x"3F7E0B6B",
    x"3F7E0AA4",
    x"3F7E09DE",
    x"3F7E0917",
    x"3F7E0850",
    x"3F7E0789",
    x"3F7E06C2",
    x"3F7E05FA",
    x"3F7E0533",
    x"3F7E046B",
    x"3F7E03A3",
    x"3F7E02DB",
    x"3F7E0213",
    x"3F7E014A",
    x"3F7E0082",
    x"3F7DFFB9",
    x"3F7DFEF0",
    x"3F7DFE28",
    x"3F7DFD5E",
    x"3F7DFC95",
    x"3F7DFBCC",
    x"3F7DFB02",
    x"3F7DFA38",
    x"3F7DF96F",
    x"3F7DF8A5",
    x"3F7DF7DA",
    x"3F7DF710",
    x"3F7DF646",
    x"3F7DF57B",
    x"3F7DF4B0",
    x"3F7DF3E5",
    x"3F7DF31A",
    x"3F7DF24F",
    x"3F7DF183",
    x"3F7DF0B8",
    x"3F7DEFEC",
    x"3F7DEF20",
    x"3F7DEE54",
    x"3F7DED88",
    x"3F7DECBC",
    x"3F7DEBEF",
    x"3F7DEB23",
    x"3F7DEA56",
    x"3F7DE989",
    x"3F7DE8BC",
    x"3F7DE7EF",
    x"3F7DE721",
    x"3F7DE654",
    x"3F7DE586",
    x"3F7DE4B8",
    x"3F7DE3EA",
    x"3F7DE31C",
    x"3F7DE24E",
    x"3F7DE17F",
    x"3F7DE0B1",
    x"3F7DDFE2",
    x"3F7DDF13",
    x"3F7DDE44",
    x"3F7DDD75",
    x"3F7DDCA5",
    x"3F7DDBD6",
    x"3F7DDB06",
    x"3F7DDA36",
    x"3F7DD966",
    x"3F7DD896",
    x"3F7DD7C6",
    x"3F7DD6F5",
    x"3F7DD625",
    x"3F7DD554",
    x"3F7DD483",
    x"3F7DD3B2",
    x"3F7DD2E1",
    x"3F7DD210",
    x"3F7DD13E",
    x"3F7DD06C",
    x"3F7DCF9B",
    x"3F7DCEC9",
    x"3F7DCDF6",
    x"3F7DCD24",
    x"3F7DCC52",
    x"3F7DCB7F",
    x"3F7DCAAC",
    x"3F7DC9DA",
    x"3F7DC906",
    x"3F7DC833",
    x"3F7DC760",
    x"3F7DC68C",
    x"3F7DC5B9",
    x"3F7DC4E5",
    x"3F7DC411",
    x"3F7DC33D",
    x"3F7DC269",
    x"3F7DC194",
    x"3F7DC0C0",
    x"3F7DBFEB",
    x"3F7DBF16",
    x"3F7DBE41",
    x"3F7DBD6C",
    x"3F7DBC96",
    x"3F7DBBC1",
    x"3F7DBAEB",
    x"3F7DBA15",
    x"3F7DB940",
    x"3F7DB869",
    x"3F7DB793",
    x"3F7DB6BD",
    x"3F7DB5E6",
    x"3F7DB510",
    x"3F7DB439",
    x"3F7DB362",
    x"3F7DB28A",
    x"3F7DB1B3",
    x"3F7DB0DC",
    x"3F7DB004",
    x"3F7DAF2C",
    x"3F7DAE54",
    x"3F7DAD7C",
    x"3F7DACA4",
    x"3F7DABCC",
    x"3F7DAAF3",
    x"3F7DAA1A",
    x"3F7DA941",
    x"3F7DA868",
    x"3F7DA78F",
    x"3F7DA6B6",
    x"3F7DA5DC",
    x"3F7DA503",
    x"3F7DA429",
    x"3F7DA34F",
    x"3F7DA275",
    x"3F7DA19B",
    x"3F7DA0C0",
    x"3F7D9FE6",
    x"3F7D9F0B",
    x"3F7D9E30",
    x"3F7D9D55",
    x"3F7D9C7A",
    x"3F7D9B9F",
    x"3F7D9AC4",
    x"3F7D99E8",
    x"3F7D990C",
    x"3F7D9830",
    x"3F7D9754",
    x"3F7D9678",
    x"3F7D959C",
    x"3F7D94BF",
    x"3F7D93E2",
    x"3F7D9306",
    x"3F7D9229",
    x"3F7D914B",
    x"3F7D906E",
    x"3F7D8F91",
    x"3F7D8EB3",
    x"3F7D8DD5",
    x"3F7D8CF8",
    x"3F7D8C19",
    x"3F7D8B3B",
    x"3F7D8A5D",
    x"3F7D897E",
    x"3F7D88A0",
    x"3F7D87C1",
    x"3F7D86E2",
    x"3F7D8603",
    x"3F7D8524",
    x"3F7D8444",
    x"3F7D8365",
    x"3F7D8285",
    x"3F7D81A5",
    x"3F7D80C5",
    x"3F7D7FE5",
    x"3F7D7F04",
    x"3F7D7E24",
    x"3F7D7D43",
    x"3F7D7C62",
    x"3F7D7B82",
    x"3F7D7AA0",
    x"3F7D79BF",
    x"3F7D78DE",
    x"3F7D77FC",
    x"3F7D771B",
    x"3F7D7639",
    x"3F7D7557",
    x"3F7D7474",
    x"3F7D7392",
    x"3F7D72B0",
    x"3F7D71CD",
    x"3F7D70EA",
    x"3F7D7007",
    x"3F7D6F24",
    x"3F7D6E41",
    x"3F7D6D5E",
    x"3F7D6C7A",
    x"3F7D6B96",
    x"3F7D6AB2",
    x"3F7D69CE",
    x"3F7D68EA",
    x"3F7D6806",
    x"3F7D6722",
    x"3F7D663D",
    x"3F7D6558",
    x"3F7D6473",
    x"3F7D638E",
    x"3F7D62A9",
    x"3F7D61C4",
    x"3F7D60DE",
    x"3F7D5FF8",
    x"3F7D5F13",
    x"3F7D5E2D",
    x"3F7D5D46",
    x"3F7D5C60",
    x"3F7D5B7A",
    x"3F7D5A93",
    x"3F7D59AC",
    x"3F7D58C5",
    x"3F7D57DE",
    x"3F7D56F7",
    x"3F7D5610",
    x"3F7D5528",
    x"3F7D5441",
    x"3F7D5359",
    x"3F7D5271",
    x"3F7D5189",
    x"3F7D50A0",
    x"3F7D4FB8",
    x"3F7D4ECF",
    x"3F7D4DE7",
    x"3F7D4CFE",
    x"3F7D4C15",
    x"3F7D4B2C",
    x"3F7D4A42",
    x"3F7D4959",
    x"3F7D486F",
    x"3F7D4785",
    x"3F7D469B",
    x"3F7D45B1",
    x"3F7D44C7",
    x"3F7D43DC",
    x"3F7D42F2",
    x"3F7D4207",
    x"3F7D411C",
    x"3F7D4031",
    x"3F7D3F46",
    x"3F7D3E5B",
    x"3F7D3D6F",
    x"3F7D3C84",
    x"3F7D3B98",
    x"3F7D3AAC",
    x"3F7D39C0",
    x"3F7D38D4",
    x"3F7D37E7",
    x"3F7D36FB",
    x"3F7D360E",
    x"3F7D3521",
    x"3F7D3434",
    x"3F7D3347",
    x"3F7D325A",
    x"3F7D316C",
    x"3F7D307F",
    x"3F7D2F91",
    x"3F7D2EA3",
    x"3F7D2DB5",
    x"3F7D2CC7",
    x"3F7D2BD8",
    x"3F7D2AEA",
    x"3F7D29FB",
    x"3F7D290C",
    x"3F7D281D",
    x"3F7D272E",
    x"3F7D263F",
    x"3F7D254F",
    x"3F7D2460",
    x"3F7D2370",
    x"3F7D2280",
    x"3F7D2190",
    x"3F7D20A0",
    x"3F7D1FAF",
    x"3F7D1EBF",
    x"3F7D1DCE",
    x"3F7D1CDD",
    x"3F7D1BEC",
    x"3F7D1AFB",
    x"3F7D1A0A",
    x"3F7D1919",
    x"3F7D1827",
    x"3F7D1735",
    x"3F7D1643",
    x"3F7D1551",
    x"3F7D145F",
    x"3F7D136D",
    x"3F7D127A",
    x"3F7D1188",
    x"3F7D1095",
    x"3F7D0FA2",
    x"3F7D0EAF",
    x"3F7D0DBC",
    x"3F7D0CC8",
    x"3F7D0BD5",
    x"3F7D0AE1",
    x"3F7D09ED",
    x"3F7D08F9",
    x"3F7D0805",
    x"3F7D0710",
    x"3F7D061C",
    x"3F7D0527",
    x"3F7D0433",
    x"3F7D033E",
    x"3F7D0249",
    x"3F7D0153",
    x"3F7D005E",
    x"3F7CFF68",
    x"3F7CFE73",
    x"3F7CFD7D",
    x"3F7CFC87",
    x"3F7CFB91",
    x"3F7CFA9A",
    x"3F7CF9A4",
    x"3F7CF8AD",
    x"3F7CF7B7",
    x"3F7CF6C0",
    x"3F7CF5C9",
    x"3F7CF4D1",
    x"3F7CF3DA",
    x"3F7CF2E2",
    x"3F7CF1EB",
    x"3F7CF0F3",
    x"3F7CEFFB",
    x"3F7CEF03",
    x"3F7CEE0B",
    x"3F7CED12",
    x"3F7CEC19",
    x"3F7CEB21",
    x"3F7CEA28",
    x"3F7CE92F",
    x"3F7CE836",
    x"3F7CE73C",
    x"3F7CE643",
    x"3F7CE549",
    x"3F7CE44F",
    x"3F7CE355",
    x"3F7CE25B",
    x"3F7CE161",
    x"3F7CE066",
    x"3F7CDF6C",
    x"3F7CDE71",
    x"3F7CDD76",
    x"3F7CDC7B",
    x"3F7CDB80",
    x"3F7CDA85",
    x"3F7CD989",
    x"3F7CD88E",
    x"3F7CD792",
    x"3F7CD696",
    x"3F7CD59A",
    x"3F7CD49E",
    x"3F7CD3A1",
    x"3F7CD2A5",
    x"3F7CD1A8",
    x"3F7CD0AB",
    x"3F7CCFAE",
    x"3F7CCEB1",
    x"3F7CCDB4",
    x"3F7CCCB6",
    x"3F7CCBB8",
    x"3F7CCABB",
    x"3F7CC9BD",
    x"3F7CC8BF",
    x"3F7CC7C0",
    x"3F7CC6C2",
    x"3F7CC5C4",
    x"3F7CC4C5",
    x"3F7CC3C6",
    x"3F7CC2C7",
    x"3F7CC1C8",
    x"3F7CC0C9",
    x"3F7CBFC9",
    x"3F7CBECA",
    x"3F7CBDCA",
    x"3F7CBCCA",
    x"3F7CBBCA",
    x"3F7CBACA",
    x"3F7CB9C9",
    x"3F7CB8C9",
    x"3F7CB7C8",
    x"3F7CB6C7",
    x"3F7CB5C6",
    x"3F7CB4C5",
    x"3F7CB3C4",
    x"3F7CB2C2",
    x"3F7CB1C1",
    x"3F7CB0BF",
    x"3F7CAFBD",
    x"3F7CAEBB",
    x"3F7CADB9",
    x"3F7CACB7",
    x"3F7CABB4",
    x"3F7CAAB2",
    x"3F7CA9AF",
    x"3F7CA8AC",
    x"3F7CA7A9",
    x"3F7CA6A6",
    x"3F7CA5A2",
    x"3F7CA49F",
    x"3F7CA39B",
    x"3F7CA297",
    x"3F7CA193",
    x"3F7CA08F",
    x"3F7C9F8A",
    x"3F7C9E86",
    x"3F7C9D81",
    x"3F7C9C7D",
    x"3F7C9B78",
    x"3F7C9A73",
    x"3F7C996D",
    x"3F7C9868",
    x"3F7C9762",
    x"3F7C965D",
    x"3F7C9557",
    x"3F7C9451",
    x"3F7C934B",
    x"3F7C9245",
    x"3F7C913E",
    x"3F7C9037",
    x"3F7C8F31",
    x"3F7C8E2A",
    x"3F7C8D23",
    x"3F7C8C1C",
    x"3F7C8B14",
    x"3F7C8A0D",
    x"3F7C8905",
    x"3F7C87FD",
    x"3F7C86F5",
    x"3F7C85ED",
    x"3F7C84E5",
    x"3F7C83DC",
    x"3F7C82D4",
    x"3F7C81CB",
    x"3F7C80C2",
    x"3F7C7FB9",
    x"3F7C7EB0",
    x"3F7C7DA7",
    x"3F7C7C9D",
    x"3F7C7B94",
    x"3F7C7A8A",
    x"3F7C7980",
    x"3F7C7876",
    x"3F7C776B",
    x"3F7C7661",
    x"3F7C7556",
    x"3F7C744C",
    x"3F7C7341",
    x"3F7C7236",
    x"3F7C712B",
    x"3F7C701F",
    x"3F7C6F14",
    x"3F7C6E08",
    x"3F7C6CFD",
    x"3F7C6BF1",
    x"3F7C6AE5",
    x"3F7C69D8",
    x"3F7C68CC",
    x"3F7C67BF",
    x"3F7C66B3",
    x"3F7C65A6",
    x"3F7C6499",
    x"3F7C638C",
    x"3F7C627E",
    x"3F7C6171",
    x"3F7C6063",
    x"3F7C5F56",
    x"3F7C5E48",
    x"3F7C5D3A",
    x"3F7C5C2C",
    x"3F7C5B1D",
    x"3F7C5A0F",
    x"3F7C5900",
    x"3F7C57F1",
    x"3F7C56E2",
    x"3F7C55D3",
    x"3F7C54C4",
    x"3F7C53B4",
    x"3F7C52A5",
    x"3F7C5195",
    x"3F7C5085",
    x"3F7C4F75",
    x"3F7C4E65",
    x"3F7C4D55",
    x"3F7C4C44",
    x"3F7C4B34",
    x"3F7C4A23",
    x"3F7C4912",
    x"3F7C4801",
    x"3F7C46F0",
    x"3F7C45DE",
    x"3F7C44CD",
    x"3F7C43BB",
    x"3F7C42A9",
    x"3F7C4197",
    x"3F7C4085",
    x"3F7C3F73",
    x"3F7C3E60",
    x"3F7C3D4E",
    x"3F7C3C3B",
    x"3F7C3B28",
    x"3F7C3A15",
    x"3F7C3902",
    x"3F7C37EE",
    x"3F7C36DB",
    x"3F7C35C7",
    x"3F7C34B3",
    x"3F7C339F",
    x"3F7C328B",
    x"3F7C3177",
    x"3F7C3062",
    x"3F7C2F4E",
    x"3F7C2E39",
    x"3F7C2D24",
    x"3F7C2C0F",
    x"3F7C2AFA",
    x"3F7C29E5",
    x"3F7C28CF",
    x"3F7C27B9",
    x"3F7C26A4",
    x"3F7C258E",
    x"3F7C2478",
    x"3F7C2361",
    x"3F7C224B",
    x"3F7C2134",
    x"3F7C201E",
    x"3F7C1F07",
    x"3F7C1DF0",
    x"3F7C1CD9",
    x"3F7C1BC1",
    x"3F7C1AAA",
    x"3F7C1992",
    x"3F7C187A",
    x"3F7C1762",
    x"3F7C164A",
    x"3F7C1532",
    x"3F7C141A",
    x"3F7C1301",
    x"3F7C11E8",
    x"3F7C10D0",
    x"3F7C0FB7",
    x"3F7C0E9D",
    x"3F7C0D84",
    x"3F7C0C6B",
    x"3F7C0B51",
    x"3F7C0A37",
    x"3F7C091E",
    x"3F7C0803",
    x"3F7C06E9",
    x"3F7C05CF",
    x"3F7C04B4",
    x"3F7C039A",
    x"3F7C027F",
    x"3F7C0164",
    x"3F7C0049",
    x"3F7BFF2E",
    x"3F7BFE12",
    x"3F7BFCF7",
    x"3F7BFBDB",
    x"3F7BFABF",
    x"3F7BF9A3",
    x"3F7BF887",
    x"3F7BF76A",
    x"3F7BF64E",
    x"3F7BF531",
    x"3F7BF415",
    x"3F7BF2F8",
    x"3F7BF1DA",
    x"3F7BF0BD",
    x"3F7BEFA0",
    x"3F7BEE82",
    x"3F7BED65",
    x"3F7BEC47",
    x"3F7BEB29",
    x"3F7BEA0B",
    x"3F7BE8EC",
    x"3F7BE7CE",
    x"3F7BE6AF",
    x"3F7BE590",
    x"3F7BE472",
    x"3F7BE353",
    x"3F7BE233",
    x"3F7BE114",
    x"3F7BDFF4",
    x"3F7BDED5",
    x"3F7BDDB5",
    x"3F7BDC95",
    x"3F7BDB75",
    x"3F7BDA55",
    x"3F7BD934",
    x"3F7BD814",
    x"3F7BD6F3",
    x"3F7BD5D2",
    x"3F7BD4B1",
    x"3F7BD390",
    x"3F7BD26E",
    x"3F7BD14D",
    x"3F7BD02B",
    x"3F7BCF09",
    x"3F7BCDE7",
    x"3F7BCCC5",
    x"3F7BCBA3",
    x"3F7BCA81",
    x"3F7BC95E",
    x"3F7BC83B",
    x"3F7BC719",
    x"3F7BC5F6",
    x"3F7BC4D2",
    x"3F7BC3AF",
    x"3F7BC28C",
    x"3F7BC168",
    x"3F7BC044",
    x"3F7BBF20",
    x"3F7BBDFC",
    x"3F7BBCD8",
    x"3F7BBBB4",
    x"3F7BBA8F",
    x"3F7BB96B",
    x"3F7BB846",
    x"3F7BB721",
    x"3F7BB5FC",
    x"3F7BB4D6",
    x"3F7BB3B1",
    x"3F7BB28B",
    x"3F7BB166",
    x"3F7BB040",
    x"3F7BAF1A",
    x"3F7BADF3",
    x"3F7BACCD",
    x"3F7BABA7",
    x"3F7BAA80",
    x"3F7BA959",
    x"3F7BA832",
    x"3F7BA70B",
    x"3F7BA5E4",
    x"3F7BA4BC",
    x"3F7BA395",
    x"3F7BA26D",
    x"3F7BA145",
    x"3F7BA01D",
    x"3F7B9EF5",
    x"3F7B9DCD",
    x"3F7B9CA4",
    x"3F7B9B7C",
    x"3F7B9A53",
    x"3F7B992A",
    x"3F7B9801",
    x"3F7B96D8",
    x"3F7B95AE",
    x"3F7B9485",
    x"3F7B935B",
    x"3F7B9231",
    x"3F7B9107",
    x"3F7B8FDD",
    x"3F7B8EB3",
    x"3F7B8D89",
    x"3F7B8C5E",
    x"3F7B8B33",
    x"3F7B8A08",
    x"3F7B88DD",
    x"3F7B87B2",
    x"3F7B8687",
    x"3F7B855B",
    x"3F7B8430",
    x"3F7B8304",
    x"3F7B81D8",
    x"3F7B80AC",
    x"3F7B7F80",
    x"3F7B7E53",
    x"3F7B7D27",
    x"3F7B7BFA",
    x"3F7B7ACD",
    x"3F7B79A0",
    x"3F7B7873",
    x"3F7B7745",
    x"3F7B7618",
    x"3F7B74EA",
    x"3F7B73BD",
    x"3F7B728F",
    x"3F7B7161",
    x"3F7B7032",
    x"3F7B6F04",
    x"3F7B6DD6",
    x"3F7B6CA7",
    x"3F7B6B78",
    x"3F7B6A49",
    x"3F7B691A",
    x"3F7B67EB",
    x"3F7B66BB",
    x"3F7B658C",
    x"3F7B645C",
    x"3F7B632C",
    x"3F7B61FC",
    x"3F7B60CC",
    x"3F7B5F9B",
    x"3F7B5E6B",
    x"3F7B5D3A",
    x"3F7B5C09",
    x"3F7B5AD9",
    x"3F7B59A7",
    x"3F7B5876",
    x"3F7B5745",
    x"3F7B5613",
    x"3F7B54E1",
    x"3F7B53B0",
    x"3F7B527E",
    x"3F7B514B",
    x"3F7B5019",
    x"3F7B4EE7",
    x"3F7B4DB4",
    x"3F7B4C81",
    x"3F7B4B4E",
    x"3F7B4A1B",
    x"3F7B48E8",
    x"3F7B47B5",
    x"3F7B4681",
    x"3F7B454E",
    x"3F7B441A",
    x"3F7B42E6",
    x"3F7B41B2",
    x"3F7B407D",
    x"3F7B3F49",
    x"3F7B3E14",
    x"3F7B3CE0",
    x"3F7B3BAB",
    x"3F7B3A76",
    x"3F7B3940",
    x"3F7B380B",
    x"3F7B36D6",
    x"3F7B35A0",
    x"3F7B346A",
    x"3F7B3334",
    x"3F7B31FE",
    x"3F7B30C8",
    x"3F7B2F92",
    x"3F7B2E5B",
    x"3F7B2D24",
    x"3F7B2BED",
    x"3F7B2AB6",
    x"3F7B297F",
    x"3F7B2848",
    x"3F7B2711",
    x"3F7B25D9",
    x"3F7B24A1",
    x"3F7B2369",
    x"3F7B2231",
    x"3F7B20F9",
    x"3F7B1FC1",
    x"3F7B1E88",
    x"3F7B1D4F",
    x"3F7B1C17",
    x"3F7B1ADE",
    x"3F7B19A4",
    x"3F7B186B",
    x"3F7B1732",
    x"3F7B15F8",
    x"3F7B14BE",
    x"3F7B1385",
    x"3F7B124B",
    x"3F7B1110",
    x"3F7B0FD6",
    x"3F7B0E9C",
    x"3F7B0D61",
    x"3F7B0C26",
    x"3F7B0AEB",
    x"3F7B09B0",
    x"3F7B0875",
    x"3F7B073A",
    x"3F7B05FE",
    x"3F7B04C2",
    x"3F7B0386",
    x"3F7B024A",
    x"3F7B010E",
    x"3F7AFFD2",
    x"3F7AFE96",
    x"3F7AFD59",
    x"3F7AFC1C",
    x"3F7AFADF",
    x"3F7AF9A2",
    x"3F7AF865",
    x"3F7AF728",
    x"3F7AF5EA",
    x"3F7AF4AD",
    x"3F7AF36F",
    x"3F7AF231",
    x"3F7AF0F3",
    x"3F7AEFB4",
    x"3F7AEE76",
    x"3F7AED37",
    x"3F7AEBF9",
    x"3F7AEABA",
    x"3F7AE97B",
    x"3F7AE83C",
    x"3F7AE6FC",
    x"3F7AE5BD",
    x"3F7AE47D",
    x"3F7AE33D",
    x"3F7AE1FE",
    x"3F7AE0BD",
    x"3F7ADF7D",
    x"3F7ADE3D",
    x"3F7ADCFC",
    x"3F7ADBBC",
    x"3F7ADA7B",
    x"3F7AD93A",
    x"3F7AD7F9",
    x"3F7AD6B7",
    x"3F7AD576",
    x"3F7AD434",
    x"3F7AD2F3",
    x"3F7AD1B1",
    x"3F7AD06F",
    x"3F7ACF2D",
    x"3F7ACDEA",
    x"3F7ACCA8",
    x"3F7ACB65",
    x"3F7ACA22",
    x"3F7AC8DF",
    x"3F7AC79C",
    x"3F7AC659",
    x"3F7AC516",
    x"3F7AC3D2",
    x"3F7AC28E",
    x"3F7AC14A",
    x"3F7AC006",
    x"3F7ABEC2",
    x"3F7ABD7E",
    x"3F7ABC3A",
    x"3F7ABAF5",
    x"3F7AB9B0",
    x"3F7AB86B",
    x"3F7AB726",
    x"3F7AB5E1",
    x"3F7AB49C",
    x"3F7AB356",
    x"3F7AB210",
    x"3F7AB0CB",
    x"3F7AAF85",
    x"3F7AAE3F",
    x"3F7AACF8",
    x"3F7AABB2",
    x"3F7AAA6B",
    x"3F7AA925",
    x"3F7AA7DE",
    x"3F7AA697",
    x"3F7AA54F",
    x"3F7AA408",
    x"3F7AA2C1",
    x"3F7AA179",
    x"3F7AA031",
    x"3F7A9EE9",
    x"3F7A9DA1",
    x"3F7A9C59",
    x"3F7A9B11",
    x"3F7A99C8",
    x"3F7A987F",
    x"3F7A9737",
    x"3F7A95EE",
    x"3F7A94A4",
    x"3F7A935B",
    x"3F7A9212",
    x"3F7A90C8",
    x"3F7A8F7E",
    x"3F7A8E34",
    x"3F7A8CEA",
    x"3F7A8BA0",
    x"3F7A8A56",
    x"3F7A890B",
    x"3F7A87C1",
    x"3F7A8676",
    x"3F7A852B",
    x"3F7A83E0",
    x"3F7A8295",
    x"3F7A8149",
    x"3F7A7FFE",
    x"3F7A7EB2",
    x"3F7A7D66",
    x"3F7A7C1A",
    x"3F7A7ACE",
    x"3F7A7982",
    x"3F7A7835",
    x"3F7A76E9",
    x"3F7A759C",
    x"3F7A744F",
    x"3F7A7302",
    x"3F7A71B5",
    x"3F7A7067",
    x"3F7A6F1A",
    x"3F7A6DCC",
    x"3F7A6C7E",
    x"3F7A6B30",
    x"3F7A69E2",
    x"3F7A6894",
    x"3F7A6745",
    x"3F7A65F7",
    x"3F7A64A8",
    x"3F7A6359",
    x"3F7A620A",
    x"3F7A60BB",
    x"3F7A5F6C",
    x"3F7A5E1C",
    x"3F7A5CCD",
    x"3F7A5B7D",
    x"3F7A5A2D",
    x"3F7A58DD",
    x"3F7A578D",
    x"3F7A563C",
    x"3F7A54EC",
    x"3F7A539B",
    x"3F7A524A",
    x"3F7A50F9",
    x"3F7A4FA8",
    x"3F7A4E57",
    x"3F7A4D05",
    x"3F7A4BB4",
    x"3F7A4A62",
    x"3F7A4910",
    x"3F7A47BE",
    x"3F7A466C",
    x"3F7A451A",
    x"3F7A43C7",
    x"3F7A4275",
    x"3F7A4122",
    x"3F7A3FCF",
    x"3F7A3E7C",
    x"3F7A3D28",
    x"3F7A3BD5",
    x"3F7A3A81",
    x"3F7A392E",
    x"3F7A37DA",
    x"3F7A3686",
    x"3F7A3532",
    x"3F7A33DD",
    x"3F7A3289",
    x"3F7A3134",
    x"3F7A2FE0",
    x"3F7A2E8B",
    x"3F7A2D36",
    x"3F7A2BE1",
    x"3F7A2A8B",
    x"3F7A2936",
    x"3F7A27E0",
    x"3F7A268A",
    x"3F7A2534",
    x"3F7A23DE",
    x"3F7A2288",
    x"3F7A2131",
    x"3F7A1FDB",
    x"3F7A1E84",
    x"3F7A1D2D",
    x"3F7A1BD6",
    x"3F7A1A7F",
    x"3F7A1928",
    x"3F7A17D0",
    x"3F7A1679",
    x"3F7A1521",
    x"3F7A13C9",
    x"3F7A1271",
    x"3F7A1119",
    x"3F7A0FC0",
    x"3F7A0E68",
    x"3F7A0D0F",
    x"3F7A0BB6",
    x"3F7A0A5D",
    x"3F7A0904",
    x"3F7A07AB",
    x"3F7A0652",
    x"3F7A04F8",
    x"3F7A039E",
    x"3F7A0244",
    x"3F7A00EA",
    x"3F79FF90",
    x"3F79FE36",
    x"3F79FCDB",
    x"3F79FB81",
    x"3F79FA26",
    x"3F79F8CB",
    x"3F79F770",
    x"3F79F615",
    x"3F79F4B9",
    x"3F79F35E",
    x"3F79F202",
    x"3F79F0A6",
    x"3F79EF4A",
    x"3F79EDEE",
    x"3F79EC92",
    x"3F79EB36",
    x"3F79E9D9",
    x"3F79E87C",
    x"3F79E71F",
    x"3F79E5C2",
    x"3F79E465",
    x"3F79E308",
    x"3F79E1AA",
    x"3F79E04D",
    x"3F79DEEF",
    x"3F79DD91",
    x"3F79DC33",
    x"3F79DAD5",
    x"3F79D976",
    x"3F79D818",
    x"3F79D6B9",
    x"3F79D55A",
    x"3F79D3FB",
    x"3F79D29C",
    x"3F79D13D",
    x"3F79CFDD",
    x"3F79CE7E",
    x"3F79CD1E",
    x"3F79CBBE",
    x"3F79CA5E",
    x"3F79C8FE",
    x"3F79C79D",
    x"3F79C63D",
    x"3F79C4DC",
    x"3F79C37B",
    x"3F79C21A",
    x"3F79C0B9",
    x"3F79BF58",
    x"3F79BDF7",
    x"3F79BC95",
    x"3F79BB33",
    x"3F79B9D2",
    x"3F79B870",
    x"3F79B70D",
    x"3F79B5AB",
    x"3F79B449",
    x"3F79B2E6",
    x"3F79B183",
    x"3F79B020",
    x"3F79AEBD",
    x"3F79AD5A",
    x"3F79ABF7",
    x"3F79AA93",
    x"3F79A930",
    x"3F79A7CC",
    x"3F79A668",
    x"3F79A504",
    x"3F79A3A0",
    x"3F79A23B",
    x"3F79A0D7",
    x"3F799F72",
    x"3F799E0D",
    x"3F799CA8",
    x"3F799B43",
    x"3F7999DE",
    x"3F799878",
    x"3F799712",
    x"3F7995AD",
    x"3F799447",
    x"3F7992E1",
    x"3F79917A",
    x"3F799014",
    x"3F798EAE",
    x"3F798D47",
    x"3F798BE0",
    x"3F798A79",
    x"3F798912",
    x"3F7987AB",
    x"3F798643",
    x"3F7984DC",
    x"3F798374",
    x"3F79820C",
    x"3F7980A4",
    x"3F797F3C",
    x"3F797DD4",
    x"3F797C6B",
    x"3F797B03",
    x"3F79799A",
    x"3F797831",
    x"3F7976C8",
    x"3F79755F",
    x"3F7973F5",
    x"3F79728C",
    x"3F797122",
    x"3F796FB8",
    x"3F796E4E",
    x"3F796CE4",
    x"3F796B7A",
    x"3F796A0F",
    x"3F7968A5",
    x"3F79673A",
    x"3F7965CF",
    x"3F796464",
    x"3F7962F9",
    x"3F79618E",
    x"3F796022",
    x"3F795EB7",
    x"3F795D4B",
    x"3F795BDF",
    x"3F795A73",
    x"3F795907",
    x"3F79579A",
    x"3F79562E",
    x"3F7954C1",
    x"3F795354",
    x"3F7951E7",
    x"3F79507A",
    x"3F794F0D",
    x"3F794D9F",
    x"3F794C32",
    x"3F794AC4",
    x"3F794956",
    x"3F7947E8",
    x"3F79467A",
    x"3F79450C",
    x"3F79439D",
    x"3F79422F",
    x"3F7940C0",
    x"3F793F51",
    x"3F793DE2",
    x"3F793C73",
    x"3F793B03",
    x"3F793994",
    x"3F793824",
    x"3F7936B4",
    x"3F793544",
    x"3F7933D4",
    x"3F793264",
    x"3F7930F3",
    x"3F792F83",
    x"3F792E12",
    x"3F792CA1",
    x"3F792B30",
    x"3F7929BF",
    x"3F79284E",
    x"3F7926DC",
    x"3F79256B",
    x"3F7923F9",
    x"3F792287",
    x"3F792115",
    x"3F791FA3",
    x"3F791E30",
    x"3F791CBE",
    x"3F791B4B",
    x"3F7919D8",
    x"3F791865",
    x"3F7916F2",
    x"3F79157F",
    x"3F79140B",
    x"3F791298",
    x"3F791124",
    x"3F790FB0",
    x"3F790E3C",
    x"3F790CC8",
    x"3F790B54",
    x"3F7909DF",
    x"3F79086A",
    x"3F7906F6",
    x"3F790581",
    x"3F79040C",
    x"3F790296",
    x"3F790121",
    x"3F78FFAC",
    x"3F78FE36",
    x"3F78FCC0",
    x"3F78FB4A",
    x"3F78F9D4",
    x"3F78F85E",
    x"3F78F6E7",
    x"3F78F571",
    x"3F78F3FA",
    x"3F78F283",
    x"3F78F10C",
    x"3F78EF95",
    x"3F78EE1D",
    x"3F78ECA6",
    x"3F78EB2E",
    x"3F78E9B7",
    x"3F78E83F",
    x"3F78E6C7",
    x"3F78E54E",
    x"3F78E3D6",
    x"3F78E25D",
    x"3F78E0E5",
    x"3F78DF6C",
    x"3F78DDF3",
    x"3F78DC7A",
    x"3F78DB01",
    x"3F78D987",
    x"3F78D80E",
    x"3F78D694",
    x"3F78D51A",
    x"3F78D3A0",
    x"3F78D226",
    x"3F78D0AB",
    x"3F78CF31",
    x"3F78CDB6",
    x"3F78CC3B",
    x"3F78CAC1",
    x"3F78C945",
    x"3F78C7CA",
    x"3F78C64F",
    x"3F78C4D3",
    x"3F78C358",
    x"3F78C1DC",
    x"3F78C060",
    x"3F78BEE4",
    x"3F78BD67",
    x"3F78BBEB",
    x"3F78BA6E",
    x"3F78B8F2",
    x"3F78B775",
    x"3F78B5F8",
    x"3F78B47B",
    x"3F78B2FD",
    x"3F78B180",
    x"3F78B002",
    x"3F78AE84",
    x"3F78AD06",
    x"3F78AB88",
    x"3F78AA0A",
    x"3F78A88C",
    x"3F78A70D",
    x"3F78A58F",
    x"3F78A410",
    x"3F78A291",
    x"3F78A112",
    x"3F789F92",
    x"3F789E13",
    x"3F789C93",
    x"3F789B14",
    x"3F789994",
    x"3F789814",
    x"3F789694",
    x"3F789513",
    x"3F789393",
    x"3F789212",
    x"3F789091",
    x"3F788F11",
    x"3F788D8F",
    x"3F788C0E",
    x"3F788A8D",
    x"3F78890B",
    x"3F78878A",
    x"3F788608",
    x"3F788486",
    x"3F788304",
    x"3F788182",
    x"3F787FFF",
    x"3F787E7D",
    x"3F787CFA",
    x"3F787B77",
    x"3F7879F4",
    x"3F787871",
    x"3F7876ED",
    x"3F78756A",
    x"3F7873E6",
    x"3F787263",
    x"3F7870DF",
    x"3F786F5B",
    x"3F786DD6",
    x"3F786C52",
    x"3F786ACE",
    x"3F786949",
    x"3F7867C4",
    x"3F78663F",
    x"3F7864BA",
    x"3F786335",
    x"3F7861AF",
    x"3F78602A",
    x"3F785EA4",
    x"3F785D1E",
    x"3F785B98",
    x"3F785A12",
    x"3F78588C",
    x"3F785705",
    x"3F78557F",
    x"3F7853F8",
    x"3F785271",
    x"3F7850EA",
    x"3F784F63",
    x"3F784DDB",
    x"3F784C54",
    x"3F784ACC",
    x"3F784944",
    x"3F7847BC",
    x"3F784634",
    x"3F7844AC",
    x"3F784324",
    x"3F78419B",
    x"3F784012",
    x"3F783E8A",
    x"3F783D01",
    x"3F783B77",
    x"3F7839EE",
    x"3F783865",
    x"3F7836DB",
    x"3F783551",
    x"3F7833C7",
    x"3F78323D",
    x"3F7830B3",
    x"3F782F29",
    x"3F782D9E",
    x"3F782C14",
    x"3F782A89",
    x"3F7828FE",
    x"3F782773",
    x"3F7825E8",
    x"3F78245C",
    x"3F7822D1",
    x"3F782145",
    x"3F781FB9",
    x"3F781E2D",
    x"3F781CA1",
    x"3F781B15",
    x"3F781988",
    x"3F7817FC",
    x"3F78166F",
    x"3F7814E2",
    x"3F781355",
    x"3F7811C8",
    x"3F78103A",
    x"3F780EAD",
    x"3F780D1F",
    x"3F780B92",
    x"3F780A04",
    x"3F780876",
    x"3F7806E7",
    x"3F780559",
    x"3F7803CA",
    x"3F78023C",
    x"3F7800AD",
    x"3F77FF1E",
    x"3F77FD8F",
    x"3F77FC00",
    x"3F77FA70",
    x"3F77F8E1",
    x"3F77F751",
    x"3F77F5C1",
    x"3F77F431",
    x"3F77F2A1",
    x"3F77F110",
    x"3F77EF80",
    x"3F77EDEF",
    x"3F77EC5F",
    x"3F77EACE",
    x"3F77E93D",
    x"3F77E7AB",
    x"3F77E61A",
    x"3F77E488",
    x"3F77E2F7",
    x"3F77E165",
    x"3F77DFD3",
    x"3F77DE41",
    x"3F77DCAF",
    x"3F77DB1C",
    x"3F77D98A",
    x"3F77D7F7",
    x"3F77D664",
    x"3F77D4D1",
    x"3F77D33E",
    x"3F77D1AB",
    x"3F77D017",
    x"3F77CE83",
    x"3F77CCF0",
    x"3F77CB5C",
    x"3F77C9C8",
    x"3F77C834",
    x"3F77C69F",
    x"3F77C50B",
    x"3F77C376",
    x"3F77C1E1",
    x"3F77C04C",
    x"3F77BEB7",
    x"3F77BD22",
    x"3F77BB8D",
    x"3F77B9F7",
    x"3F77B861",
    x"3F77B6CB",
    x"3F77B535",
    x"3F77B39F",
    x"3F77B209",
    x"3F77B073",
    x"3F77AEDC",
    x"3F77AD45",
    x"3F77ABAE",
    x"3F77AA17",
    x"3F77A880",
    x"3F77A6E9",
    x"3F77A551",
    x"3F77A3BA",
    x"3F77A222",
    x"3F77A08A",
    x"3F779EF2",
    x"3F779D5A",
    x"3F779BC1",
    x"3F779A29",
    x"3F779890",
    x"3F7796F7",
    x"3F77955E",
    x"3F7793C5",
    x"3F77922C",
    x"3F779092",
    x"3F778EF9",
    x"3F778D5F",
    x"3F778BC5",
    x"3F778A2B",
    x"3F778891",
    x"3F7786F7",
    x"3F77855C",
    x"3F7783C2",
    x"3F778227",
    x"3F77808C",
    x"3F777EF1",
    x"3F777D56",
    x"3F777BBA",
    x"3F777A1F",
    x"3F777883",
    x"3F7776E7",
    x"3F77754B",
    x"3F7773AF",
    x"3F777213",
    x"3F777076",
    x"3F776EDA",
    x"3F776D3D",
    x"3F776BA0",
    x"3F776A03",
    x"3F776866",
    x"3F7766C9",
    x"3F77652B",
    x"3F77638E",
    x"3F7761F0",
    x"3F776052",
    x"3F775EB4",
    x"3F775D16",
    x"3F775B78",
    x"3F7759D9",
    x"3F77583A",
    x"3F77569C",
    x"3F7754FD",
    x"3F77535E",
    x"3F7751BE",
    x"3F77501F",
    x"3F774E7F",
    x"3F774CE0",
    x"3F774B40",
    x"3F7749A0",
    x"3F774800",
    x"3F77465F",
    x"3F7744BF",
    x"3F77431E",
    x"3F77417E",
    x"3F773FDD",
    x"3F773E3C",
    x"3F773C9B",
    x"3F773AF9",
    x"3F773958",
    x"3F7737B6",
    x"3F773614",
    x"3F773472",
    x"3F7732D0",
    x"3F77312E",
    x"3F772F8C",
    x"3F772DE9",
    x"3F772C47",
    x"3F772AA4",
    x"3F772901",
    x"3F77275E",
    x"3F7725BA",
    x"3F772417",
    x"3F772274",
    x"3F7720D0",
    x"3F771F2C",
    x"3F771D88",
    x"3F771BE4",
    x"3F771A3F",
    x"3F77189B",
    x"3F7716F6",
    x"3F771552",
    x"3F7713AD",
    x"3F771208",
    x"3F771063",
    x"3F770EBD",
    x"3F770D18",
    x"3F770B72",
    x"3F7709CC",
    x"3F770826",
    x"3F770680",
    x"3F7704DA",
    x"3F770334",
    x"3F77018D",
    x"3F76FFE6",
    x"3F76FE40",
    x"3F76FC99",
    x"3F76FAF1",
    x"3F76F94A",
    x"3F76F7A3",
    x"3F76F5FB",
    x"3F76F453",
    x"3F76F2AC",
    x"3F76F103",
    x"3F76EF5B",
    x"3F76EDB3",
    x"3F76EC0B",
    x"3F76EA62",
    x"3F76E8B9",
    x"3F76E710",
    x"3F76E567",
    x"3F76E3BE",
    x"3F76E215",
    x"3F76E06B",
    x"3F76DEC1",
    x"3F76DD18",
    x"3F76DB6E",
    x"3F76D9C4",
    x"3F76D819",
    x"3F76D66F",
    x"3F76D4C4",
    x"3F76D31A",
    x"3F76D16F",
    x"3F76CFC4",
    x"3F76CE19",
    x"3F76CC6D",
    x"3F76CAC2",
    x"3F76C916",
    x"3F76C76B",
    x"3F76C5BF",
    x"3F76C413",
    x"3F76C266",
    x"3F76C0BA",
    x"3F76BF0E",
    x"3F76BD61",
    x"3F76BBB4",
    x"3F76BA07",
    x"3F76B85A",
    x"3F76B6AD",
    x"3F76B500",
    x"3F76B352",
    x"3F76B1A4",
    x"3F76AFF7",
    x"3F76AE49",
    x"3F76AC9A",
    x"3F76AAEC",
    x"3F76A93E",
    x"3F76A78F",
    x"3F76A5E0",
    x"3F76A432",
    x"3F76A283",
    x"3F76A0D3",
    x"3F769F24",
    x"3F769D75",
    x"3F769BC5",
    x"3F769A15",
    x"3F769865",
    x"3F7696B5",
    x"3F769505",
    x"3F769355",
    x"3F7691A4",
    x"3F768FF4",
    x"3F768E43",
    x"3F768C92",
    x"3F768AE1",
    x"3F768930",
    x"3F76877E",
    x"3F7685CD",
    x"3F76841B",
    x"3F768269",
    x"3F7680B7",
    x"3F767F05",
    x"3F767D53",
    x"3F767BA0",
    x"3F7679EE",
    x"3F76783B",
    x"3F767688",
    x"3F7674D5",
    x"3F767322",
    x"3F76716F",
    x"3F766FBB",
    x"3F766E08",
    x"3F766C54",
    x"3F766AA0",
    x"3F7668EC",
    x"3F766738",
    x"3F766583",
    x"3F7663CF",
    x"3F76621A",
    x"3F766065",
    x"3F765EB0",
    x"3F765CFB",
    x"3F765B46",
    x"3F765991",
    x"3F7657DB",
    x"3F765625",
    x"3F76546F",
    x"3F7652B9",
    x"3F765103",
    x"3F764F4D",
    x"3F764D97",
    x"3F764BE0",
    x"3F764A29",
    x"3F764872",
    x"3F7646BB",
    x"3F764504",
    x"3F76434D",
    x"3F764195",
    x"3F763FDE",
    x"3F763E26",
    x"3F763C6E",
    x"3F763AB6",
    x"3F7638FE",
    x"3F763745",
    x"3F76358D",
    x"3F7633D4",
    x"3F76321B",
    x"3F763063",
    x"3F762EA9",
    x"3F762CF0",
    x"3F762B37",
    x"3F76297D",
    x"3F7627C3",
    x"3F76260A",
    x"3F762450",
    x"3F762296",
    x"3F7620DB",
    x"3F761F21",
    x"3F761D66",
    x"3F761BAB",
    x"3F7619F1",
    x"3F761836",
    x"3F76167A",
    x"3F7614BF",
    x"3F761304",
    x"3F761148",
    x"3F760F8C",
    x"3F760DD0",
    x"3F760C14",
    x"3F760A58",
    x"3F76089C",
    x"3F7606DF",
    x"3F760522",
    x"3F760366",
    x"3F7601A9",
    x"3F75FFEB",
    x"3F75FE2E",
    x"3F75FC71",
    x"3F75FAB3",
    x"3F75F8F6",
    x"3F75F738",
    x"3F75F57A",
    x"3F75F3BC",
    x"3F75F1FD",
    x"3F75F03F",
    x"3F75EE80",
    x"3F75ECC2",
    x"3F75EB03",
    x"3F75E944",
    x"3F75E784",
    x"3F75E5C5",
    x"3F75E406",
    x"3F75E246",
    x"3F75E086",
    x"3F75DEC6",
    x"3F75DD06",
    x"3F75DB46",
    x"3F75D986",
    x"3F75D7C5",
    x"3F75D604",
    x"3F75D444",
    x"3F75D283",
    x"3F75D0C2",
    x"3F75CF00",
    x"3F75CD3F",
    x"3F75CB7D",
    x"3F75C9BC",
    x"3F75C7FA",
    x"3F75C638",
    x"3F75C476",
    x"3F75C2B3",
    x"3F75C0F1",
    x"3F75BF2E",
    x"3F75BD6C",
    x"3F75BBA9",
    x"3F75B9E6",
    x"3F75B822",
    x"3F75B65F",
    x"3F75B49C",
    x"3F75B2D8",
    x"3F75B114",
    x"3F75AF50",
    x"3F75AD8C",
    x"3F75ABC8",
    x"3F75AA04",
    x"3F75A83F",
    x"3F75A67B",
    x"3F75A4B6",
    x"3F75A2F1",
    x"3F75A12C",
    x"3F759F66",
    x"3F759DA1",
    x"3F759BDB",
    x"3F759A16",
    x"3F759850",
    x"3F75968A",
    x"3F7594C4",
    x"3F7592FE",
    x"3F759137",
    x"3F758F70",
    x"3F758DAA",
    x"3F758BE3",
    x"3F758A1C",
    x"3F758855",
    x"3F75868D",
    x"3F7584C6",
    x"3F7582FE",
    x"3F758136",
    x"3F757F6F",
    x"3F757DA7",
    x"3F757BDE",
    x"3F757A16",
    x"3F75784D",
    x"3F757685",
    x"3F7574BC",
    x"3F7572F3",
    x"3F75712A",
    x"3F756F61",
    x"3F756D97",
    x"3F756BCE",
    x"3F756A04",
    x"3F75683A",
    x"3F756670",
    x"3F7564A6",
    x"3F7562DC",
    x"3F756111",
    x"3F755F47",
    x"3F755D7C",
    x"3F755BB1",
    x"3F7559E6",
    x"3F75581B",
    x"3F755650",
    x"3F755484",
    x"3F7552B9",
    x"3F7550ED",
    x"3F754F21",
    x"3F754D55",
    x"3F754B89",
    x"3F7549BC",
    x"3F7547F0",
    x"3F754623",
    x"3F754456",
    x"3F754289",
    x"3F7540BC",
    x"3F753EEF",
    x"3F753D22",
    x"3F753B54",
    x"3F753987",
    x"3F7537B9",
    x"3F7535EB",
    x"3F75341D",
    x"3F75324E",
    x"3F753080",
    x"3F752EB1",
    x"3F752CE3",
    x"3F752B14",
    x"3F752945",
    x"3F752776",
    x"3F7525A6",
    x"3F7523D7",
    x"3F752207",
    x"3F752038",
    x"3F751E68",
    x"3F751C98",
    x"3F751AC7",
    x"3F7518F7",
    x"3F751727",
    x"3F751556",
    x"3F751385",
    x"3F7511B4",
    x"3F750FE3",
    x"3F750E12",
    x"3F750C41",
    x"3F750A6F",
    x"3F75089D",
    x"3F7506CC",
    x"3F7504FA",
    x"3F750327",
    x"3F750155",
    x"3F74FF83",
    x"3F74FDB0",
    x"3F74FBDE",
    x"3F74FA0B",
    x"3F74F838",
    x"3F74F665",
    x"3F74F491",
    x"3F74F2BE",
    x"3F74F0EA",
    x"3F74EF17",
    x"3F74ED43",
    x"3F74EB6F",
    x"3F74E99A",
    x"3F74E7C6",
    x"3F74E5F2",
    x"3F74E41D",
    x"3F74E248",
    x"3F74E073",
    x"3F74DE9E",
    x"3F74DCC9",
    x"3F74DAF4",
    x"3F74D91E",
    x"3F74D749",
    x"3F74D573",
    x"3F74D39D",
    x"3F74D1C7",
    x"3F74CFF0",
    x"3F74CE1A",
    x"3F74CC44",
    x"3F74CA6D",
    x"3F74C896",
    x"3F74C6BF",
    x"3F74C4E8",
    x"3F74C311",
    x"3F74C139",
    x"3F74BF62",
    x"3F74BD8A",
    x"3F74BBB2",
    x"3F74B9DA",
    x"3F74B802",
    x"3F74B62A",
    x"3F74B451",
    x"3F74B279",
    x"3F74B0A0",
    x"3F74AEC7",
    x"3F74ACEE",
    x"3F74AB15",
    x"3F74A93B",
    x"3F74A762",
    x"3F74A588",
    x"3F74A3AE",
    x"3F74A1D5",
    x"3F749FFA",
    x"3F749E20",
    x"3F749C46",
    x"3F749A6B",
    x"3F749891",
    x"3F7496B6",
    x"3F7494DB",
    x"3F749300",
    x"3F749125",
    x"3F748F49",
    x"3F748D6E",
    x"3F748B92",
    x"3F7489B6",
    x"3F7487DA",
    x"3F7485FE",
    x"3F748422",
    x"3F748245",
    x"3F748069",
    x"3F747E8C",
    x"3F747CAF",
    x"3F747AD2",
    x"3F7478F5",
    x"3F747718",
    x"3F74753A",
    x"3F74735D",
    x"3F74717F",
    x"3F746FA1",
    x"3F746DC3",
    x"3F746BE5",
    x"3F746A06",
    x"3F746828",
    x"3F746649",
    x"3F74646A",
    x"3F74628B",
    x"3F7460AC",
    x"3F745ECD",
    x"3F745CEE",
    x"3F745B0E",
    x"3F74592F",
    x"3F74574F",
    x"3F74556F",
    x"3F74538F",
    x"3F7451AE",
    x"3F744FCE",
    x"3F744DED",
    x"3F744C0D",
    x"3F744A2C",
    x"3F74484B",
    x"3F74466A",
    x"3F744488",
    x"3F7442A7",
    x"3F7440C5",
    x"3F743EE4",
    x"3F743D02",
    x"3F743B20",
    x"3F74393E",
    x"3F74375B",
    x"3F743579",
    x"3F743396",
    x"3F7431B3",
    x"3F742FD1",
    x"3F742DED",
    x"3F742C0A",
    x"3F742A27",
    x"3F742843",
    x"3F742660",
    x"3F74247C",
    x"3F742298",
    x"3F7420B4",
    x"3F741ED0",
    x"3F741CEB",
    x"3F741B07",
    x"3F741922",
    x"3F74173D",
    x"3F741558",
    x"3F741373",
    x"3F74118E",
    x"3F740FA9",
    x"3F740DC3",
    x"3F740BDD",
    x"3F7409F8",
    x"3F740812",
    x"3F74062B",
    x"3F740445",
    x"3F74025F",
    x"3F740078",
    x"3F73FE91",
    x"3F73FCAA",
    x"3F73FAC3",
    x"3F73F8DC",
    x"3F73F6F5",
    x"3F73F50D",
    x"3F73F326",
    x"3F73F13E",
    x"3F73EF56",
    x"3F73ED6E",
    x"3F73EB86",
    x"3F73E99E",
    x"3F73E7B5",
    x"3F73E5CC",
    x"3F73E3E4",
    x"3F73E1FB",
    x"3F73E012",
    x"3F73DE28",
    x"3F73DC3F",
    x"3F73DA56",
    x"3F73D86C",
    x"3F73D682",
    x"3F73D498",
    x"3F73D2AE",
    x"3F73D0C4",
    x"3F73CED9",
    x"3F73CCEF",
    x"3F73CB04",
    x"3F73C919",
    x"3F73C72E",
    x"3F73C543",
    x"3F73C358",
    x"3F73C16C",
    x"3F73BF81",
    x"3F73BD95",
    x"3F73BBA9",
    x"3F73B9BD",
    x"3F73B7D1",
    x"3F73B5E5",
    x"3F73B3F8",
    x"3F73B20C",
    x"3F73B01F",
    x"3F73AE32",
    x"3F73AC45",
    x"3F73AA58",
    x"3F73A86A",
    x"3F73A67D",
    x"3F73A48F",
    x"3F73A2A1",
    x"3F73A0B4",
    x"3F739EC5",
    x"3F739CD7",
    x"3F739AE9",
    x"3F7398FA",
    x"3F73970C",
    x"3F73951D",
    x"3F73932E",
    x"3F73913F",
    x"3F738F50",
    x"3F738D60",
    x"3F738B71",
    x"3F738981",
    x"3F738791",
    x"3F7385A1",
    x"3F7383B1",
    x"3F7381C1",
    x"3F737FD0",
    x"3F737DE0",
    x"3F737BEF",
    x"3F7379FE",
    x"3F73780D",
    x"3F73761C",
    x"3F73742B",
    x"3F737239",
    x"3F737048",
    x"3F736E56",
    x"3F736C64",
    x"3F736A72",
    x"3F736880",
    x"3F73668E",
    x"3F73649B",
    x"3F7362A8",
    x"3F7360B6",
    x"3F735EC3",
    x"3F735CD0",
    x"3F735ADC",
    x"3F7358E9",
    x"3F7356F6",
    x"3F735502",
    x"3F73530E",
    x"3F73511A",
    x"3F734F26",
    x"3F734D32",
    x"3F734B3E",
    x"3F734949",
    x"3F734754",
    x"3F734560",
    x"3F73436B",
    x"3F734175",
    x"3F733F80",
    x"3F733D8B",
    x"3F733B95",
    x"3F7339A0",
    x"3F7337AA",
    x"3F7335B4",
    x"3F7333BE",
    x"3F7331C7",
    x"3F732FD1",
    x"3F732DDA",
    x"3F732BE4",
    x"3F7329ED",
    x"3F7327F6",
    x"3F7325FE",
    x"3F732407",
    x"3F732210",
    x"3F732018",
    x"3F731E20",
    x"3F731C28",
    x"3F731A30",
    x"3F731838",
    x"3F731640",
    x"3F731447",
    x"3F73124F",
    x"3F731056",
    x"3F730E5D",
    x"3F730C64",
    x"3F730A6B",
    x"3F730871",
    x"3F730678",
    x"3F73047E",
    x"3F730284",
    x"3F73008B",
    x"3F72FE90",
    x"3F72FC96",
    x"3F72FA9C",
    x"3F72F8A1",
    x"3F72F6A7",
    x"3F72F4AC",
    x"3F72F2B1",
    x"3F72F0B6",
    x"3F72EEBA",
    x"3F72ECBF",
    x"3F72EAC3",
    x"3F72E8C8",
    x"3F72E6CC",
    x"3F72E4D0",
    x"3F72E2D4",
    x"3F72E0D7",
    x"3F72DEDB",
    x"3F72DCDE",
    x"3F72DAE2",
    x"3F72D8E5",
    x"3F72D6E8",
    x"3F72D4EB",
    x"3F72D2ED",
    x"3F72D0F0",
    x"3F72CEF2",
    x"3F72CCF5",
    x"3F72CAF7",
    x"3F72C8F9",
    x"3F72C6FA",
    x"3F72C4FC",
    x"3F72C2FE",
    x"3F72C0FF",
    x"3F72BF00",
    x"3F72BD01",
    x"3F72BB02",
    x"3F72B903",
    x"3F72B704",
    x"3F72B504",
    x"3F72B304",
    x"3F72B105",
    x"3F72AF05",
    x"3F72AD05",
    x"3F72AB04",
    x"3F72A904",
    x"3F72A703",
    x"3F72A503",
    x"3F72A302",
    x"3F72A101",
    x"3F729F00",
    x"3F729CFF",
    x"3F729AFD",
    x"3F7298FC",
    x"3F7296FA",
    x"3F7294F8",
    x"3F7292F6",
    x"3F7290F4",
    x"3F728EF2",
    x"3F728CEF",
    x"3F728AED",
    x"3F7288EA",
    x"3F7286E7",
    x"3F7284E4",
    x"3F7282E1",
    x"3F7280DE",
    x"3F727EDA",
    x"3F727CD7",
    x"3F727AD3",
    x"3F7278CF",
    x"3F7276CB",
    x"3F7274C7",
    x"3F7272C2",
    x"3F7270BE",
    x"3F726EB9",
    x"3F726CB5",
    x"3F726AB0",
    x"3F7268AB",
    x"3F7266A5",
    x"3F7264A0",
    x"3F72629B",
    x"3F726095",
    x"3F725E8F",
    x"3F725C89",
    x"3F725A83",
    x"3F72587D",
    x"3F725677",
    x"3F725470",
    x"3F725269",
    x"3F725063",
    x"3F724E5C",
    x"3F724C54",
    x"3F724A4D",
    x"3F724846",
    x"3F72463E",
    x"3F724437",
    x"3F72422F",
    x"3F724027",
    x"3F723E1F",
    x"3F723C16",
    x"3F723A0E",
    x"3F723805",
    x"3F7235FD",
    x"3F7233F4",
    x"3F7231EB",
    x"3F722FE2",
    x"3F722DD8",
    x"3F722BCF",
    x"3F7229C5",
    x"3F7227BC",
    x"3F7225B2",
    x"3F7223A8",
    x"3F72219E",
    x"3F721F93",
    x"3F721D89",
    x"3F721B7E",
    x"3F721973",
    x"3F721769",
    x"3F72155E",
    x"3F721352",
    x"3F721147",
    x"3F720F3C",
    x"3F720D30",
    x"3F720B24",
    x"3F720918",
    x"3F72070C",
    x"3F720500",
    x"3F7202F4",
    x"3F7200E7",
    x"3F71FEDA",
    x"3F71FCCE",
    x"3F71FAC1",
    x"3F71F8B4",
    x"3F71F6A6",
    x"3F71F499",
    x"3F71F28C",
    x"3F71F07E",
    x"3F71EE70",
    x"3F71EC62",
    x"3F71EA54",
    x"3F71E846",
    x"3F71E637",
    x"3F71E429",
    x"3F71E21A",
    x"3F71E00B",
    x"3F71DDFC",
    x"3F71DBED",
    x"3F71D9DE",
    x"3F71D7CF",
    x"3F71D5BF",
    x"3F71D3AF",
    x"3F71D19F",
    x"3F71CF8F",
    x"3F71CD7F",
    x"3F71CB6F",
    x"3F71C95F",
    x"3F71C74E",
    x"3F71C53D",
    x"3F71C32C",
    x"3F71C11B",
    x"3F71BF0A",
    x"3F71BCF9",
    x"3F71BAE7",
    x"3F71B8D6",
    x"3F71B6C4",
    x"3F71B4B2",
    x"3F71B2A0",
    x"3F71B08E",
    x"3F71AE7C",
    x"3F71AC69",
    x"3F71AA57",
    x"3F71A844",
    x"3F71A631",
    x"3F71A41E",
    x"3F71A20B",
    x"3F719FF7",
    x"3F719DE4",
    x"3F719BD0",
    x"3F7199BC",
    x"3F7197A8",
    x"3F719594",
    x"3F719380",
    x"3F71916C",
    x"3F718F57",
    x"3F718D43",
    x"3F718B2E",
    x"3F718919",
    x"3F718704",
    x"3F7184EF",
    x"3F7182D9",
    x"3F7180C4",
    x"3F717EAE",
    x"3F717C98",
    x"3F717A82",
    x"3F71786C",
    x"3F717656",
    x"3F71743F",
    x"3F717229",
    x"3F717012",
    x"3F716DFB",
    x"3F716BE4",
    x"3F7169CD",
    x"3F7167B6",
    x"3F71659F",
    x"3F716387",
    x"3F71616F",
    x"3F715F57",
    x"3F715D3F",
    x"3F715B27",
    x"3F71590F",
    x"3F7156F6",
    x"3F7154DE",
    x"3F7152C5",
    x"3F7150AC",
    x"3F714E93",
    x"3F714C7A",
    x"3F714A61",
    x"3F714847",
    x"3F71462E",
    x"3F714414",
    x"3F7141FA",
    x"3F713FE0",
    x"3F713DC6",
    x"3F713BAC",
    x"3F713991",
    x"3F713776",
    x"3F71355C",
    x"3F713341",
    x"3F713126",
    x"3F712F0B",
    x"3F712CEF",
    x"3F712AD4",
    x"3F7128B8",
    x"3F71269C",
    x"3F712480",
    x"3F712264",
    x"3F712048",
    x"3F711E2C",
    x"3F711C0F",
    x"3F7119F3",
    x"3F7117D6",
    x"3F7115B9",
    x"3F71139C",
    x"3F71117F",
    x"3F710F61",
    x"3F710D44",
    x"3F710B26",
    x"3F710908",
    x"3F7106EA",
    x"3F7104CC",
    x"3F7102AE",
    x"3F71008F",
    x"3F70FE71",
    x"3F70FC52",
    x"3F70FA33",
    x"3F70F814",
    x"3F70F5F5",
    x"3F70F3D6",
    x"3F70F1B7",
    x"3F70EF97",
    x"3F70ED77",
    x"3F70EB58",
    x"3F70E938",
    x"3F70E717",
    x"3F70E4F7",
    x"3F70E2D7",
    x"3F70E0B6",
    x"3F70DE95",
    x"3F70DC75",
    x"3F70DA54",
    x"3F70D832",
    x"3F70D611",
    x"3F70D3F0",
    x"3F70D1CE",
    x"3F70CFAC",
    x"3F70CD8A",
    x"3F70CB68",
    x"3F70C946",
    x"3F70C724",
    x"3F70C501",
    x"3F70C2DF",
    x"3F70C0BC",
    x"3F70BE99",
    x"3F70BC76",
    x"3F70BA53",
    x"3F70B830",
    x"3F70B60C",
    x"3F70B3E9",
    x"3F70B1C5",
    x"3F70AFA1",
    x"3F70AD7D",
    x"3F70AB59",
    x"3F70A934",
    x"3F70A710",
    x"3F70A4EB",
    x"3F70A2C6",
    x"3F70A0A2",
    x"3F709E7C",
    x"3F709C57",
    x"3F709A32",
    x"3F70980C",
    x"3F7095E7",
    x"3F7093C1",
    x"3F70919B",
    x"3F708F75",
    x"3F708D4F",
    x"3F708B28",
    x"3F708902",
    x"3F7086DB",
    x"3F7084B4",
    x"3F70828D",
    x"3F708066",
    x"3F707E3F",
    x"3F707C18",
    x"3F7079F0",
    x"3F7077C8",
    x"3F7075A1",
    x"3F707379",
    x"3F707151",
    x"3F706F28",
    x"3F706D00",
    x"3F706AD7",
    x"3F7068AF",
    x"3F706686",
    x"3F70645D",
    x"3F706234",
    x"3F70600A",
    x"3F705DE1",
    x"3F705BB8",
    x"3F70598E",
    x"3F705764",
    x"3F70553A",
    x"3F705310",
    x"3F7050E6",
    x"3F704EBB",
    x"3F704C91",
    x"3F704A66",
    x"3F70483B",
    x"3F704610",
    x"3F7043E5",
    x"3F7041BA",
    x"3F703F8E",
    x"3F703D63",
    x"3F703B37",
    x"3F70390B",
    x"3F7036DF",
    x"3F7034B3",
    x"3F703286",
    x"3F70305A",
    x"3F702E2D",
    x"3F702C01",
    x"3F7029D4",
    x"3F7027A7",
    x"3F70257A",
    x"3F70234C",
    x"3F70211F",
    x"3F701EF1",
    x"3F701CC3",
    x"3F701A95",
    x"3F701867",
    x"3F701639",
    x"3F70140B",
    x"3F7011DC",
    x"3F700FAE",
    x"3F700D7F",
    x"3F700B50",
    x"3F700921",
    x"3F7006F2",
    x"3F7004C3",
    x"3F700293",
    x"3F700063",
    x"3F6FFE34",
    x"3F6FFC04",
    x"3F6FF9D4",
    x"3F6FF7A3",
    x"3F6FF573",
    x"3F6FF343",
    x"3F6FF112",
    x"3F6FEEE1",
    x"3F6FECB0",
    x"3F6FEA7F",
    x"3F6FE84E",
    x"3F6FE61D",
    x"3F6FE3EB",
    x"3F6FE1B9",
    x"3F6FDF88",
    x"3F6FDD56",
    x"3F6FDB24",
    x"3F6FD8F1",
    x"3F6FD6BF",
    x"3F6FD48C",
    x"3F6FD25A",
    x"3F6FD027",
    x"3F6FCDF4",
    x"3F6FCBC1",
    x"3F6FC98E",
    x"3F6FC75A",
    x"3F6FC527",
    x"3F6FC2F3",
    x"3F6FC0BF",
    x"3F6FBE8B",
    x"3F6FBC57",
    x"3F6FBA23",
    x"3F6FB7EE",
    x"3F6FB5BA",
    x"3F6FB385",
    x"3F6FB150",
    x"3F6FAF1B",
    x"3F6FACE6",
    x"3F6FAAB1",
    x"3F6FA87C",
    x"3F6FA646",
    x"3F6FA410",
    x"3F6FA1DA",
    x"3F6F9FA4",
    x"3F6F9D6E",
    x"3F6F9B38",
    x"3F6F9902",
    x"3F6F96CB",
    x"3F6F9494",
    x"3F6F925D",
    x"3F6F9026",
    x"3F6F8DEF",
    x"3F6F8BB8",
    x"3F6F8981",
    x"3F6F8749",
    x"3F6F8511",
    x"3F6F82D9",
    x"3F6F80A1",
    x"3F6F7E69",
    x"3F6F7C31",
    x"3F6F79F8",
    x"3F6F77C0",
    x"3F6F7587",
    x"3F6F734E",
    x"3F6F7115",
    x"3F6F6EDC",
    x"3F6F6CA3",
    x"3F6F6A69",
    x"3F6F6830",
    x"3F6F65F6",
    x"3F6F63BC",
    x"3F6F6182",
    x"3F6F5F48",
    x"3F6F5D0E",
    x"3F6F5AD3",
    x"3F6F5899",
    x"3F6F565E",
    x"3F6F5423",
    x"3F6F51E8",
    x"3F6F4FAD",
    x"3F6F4D71",
    x"3F6F4B36",
    x"3F6F48FA",
    x"3F6F46BE",
    x"3F6F4483",
    x"3F6F4247",
    x"3F6F400A",
    x"3F6F3DCE",
    x"3F6F3B92",
    x"3F6F3955",
    x"3F6F3718",
    x"3F6F34DB",
    x"3F6F329E",
    x"3F6F3061",
    x"3F6F2E24",
    x"3F6F2BE6",
    x"3F6F29A8",
    x"3F6F276B",
    x"3F6F252D",
    x"3F6F22EF",
    x"3F6F20B0",
    x"3F6F1E72",
    x"3F6F1C34",
    x"3F6F19F5",
    x"3F6F17B6",
    x"3F6F1577",
    x"3F6F1338",
    x"3F6F10F9",
    x"3F6F0EBA",
    x"3F6F0C7A",
    x"3F6F0A3A",
    x"3F6F07FB",
    x"3F6F05BB",
    x"3F6F037B",
    x"3F6F013A",
    x"3F6EFEFA",
    x"3F6EFCBA",
    x"3F6EFA79",
    x"3F6EF838",
    x"3F6EF5F7",
    x"3F6EF3B6",
    x"3F6EF175",
    x"3F6EEF33",
    x"3F6EECF2",
    x"3F6EEAB0",
    x"3F6EE86E",
    x"3F6EE62C",
    x"3F6EE3EA",
    x"3F6EE1A8",
    x"3F6EDF66",
    x"3F6EDD23",
    x"3F6EDAE1",
    x"3F6ED89E",
    x"3F6ED65B",
    x"3F6ED418",
    x"3F6ED1D4",
    x"3F6ECF91",
    x"3F6ECD4D",
    x"3F6ECB0A",
    x"3F6EC8C6",
    x"3F6EC682",
    x"3F6EC43E",
    x"3F6EC1FA",
    x"3F6EBFB5",
    x"3F6EBD71",
    x"3F6EBB2C",
    x"3F6EB8E7",
    x"3F6EB6A2",
    x"3F6EB45D",
    x"3F6EB218",
    x"3F6EAFD2",
    x"3F6EAD8D",
    x"3F6EAB47",
    x"3F6EA901",
    x"3F6EA6BB",
    x"3F6EA475",
    x"3F6EA22F",
    x"3F6E9FE9",
    x"3F6E9DA2",
    x"3F6E9B5B",
    x"3F6E9914",
    x"3F6E96CD",
    x"3F6E9486",
    x"3F6E923F",
    x"3F6E8FF8",
    x"3F6E8DB0",
    x"3F6E8B68",
    x"3F6E8920",
    x"3F6E86D8",
    x"3F6E8490",
    x"3F6E8248",
    x"3F6E8000",
    x"3F6E7DB7",
    x"3F6E7B6E",
    x"3F6E7926",
    x"3F6E76DD",
    x"3F6E7493",
    x"3F6E724A",
    x"3F6E7001",
    x"3F6E6DB7",
    x"3F6E6B6D",
    x"3F6E6924",
    x"3F6E66D9",
    x"3F6E648F",
    x"3F6E6245",
    x"3F6E5FFB",
    x"3F6E5DB0",
    x"3F6E5B65",
    x"3F6E591A",
    x"3F6E56CF",
    x"3F6E5484",
    x"3F6E5239",
    x"3F6E4FEE",
    x"3F6E4DA2",
    x"3F6E4B56",
    x"3F6E490A",
    x"3F6E46BE",
    x"3F6E4472",
    x"3F6E4226",
    x"3F6E3FD9",
    x"3F6E3D8D",
    x"3F6E3B40",
    x"3F6E38F3",
    x"3F6E36A6",
    x"3F6E3459",
    x"3F6E320C",
    x"3F6E2FBE",
    x"3F6E2D71",
    x"3F6E2B23",
    x"3F6E28D5",
    x"3F6E2687",
    x"3F6E2439",
    x"3F6E21EB",
    x"3F6E1F9C",
    x"3F6E1D4E",
    x"3F6E1AFF",
    x"3F6E18B0",
    x"3F6E1661",
    x"3F6E1412",
    x"3F6E11C2",
    x"3F6E0F73",
    x"3F6E0D23",
    x"3F6E0AD4",
    x"3F6E0884",
    x"3F6E0634",
    x"3F6E03E3",
    x"3F6E0193",
    x"3F6DFF43",
    x"3F6DFCF2",
    x"3F6DFAA1",
    x"3F6DF850",
    x"3F6DF5FF",
    x"3F6DF3AE",
    x"3F6DF15D",
    x"3F6DEF0B",
    x"3F6DECBA",
    x"3F6DEA68",
    x"3F6DE816",
    x"3F6DE5C4",
    x"3F6DE372",
    x"3F6DE120",
    x"3F6DDECD",
    x"3F6DDC7B",
    x"3F6DDA28",
    x"3F6DD7D5",
    x"3F6DD582",
    x"3F6DD32F",
    x"3F6DD0DB",
    x"3F6DCE88",
    x"3F6DCC34",
    x"3F6DC9E1",
    x"3F6DC78D",
    x"3F6DC539",
    x"3F6DC2E4",
    x"3F6DC090",
    x"3F6DBE3C",
    x"3F6DBBE7",
    x"3F6DB992",
    x"3F6DB73D",
    x"3F6DB4E8",
    x"3F6DB293",
    x"3F6DB03E",
    x"3F6DADE8",
    x"3F6DAB93",
    x"3F6DA93D",
    x"3F6DA6E7",
    x"3F6DA491",
    x"3F6DA23B",
    x"3F6D9FE4",
    x"3F6D9D8E",
    x"3F6D9B37",
    x"3F6D98E1",
    x"3F6D968A",
    x"3F6D9433",
    x"3F6D91DB",
    x"3F6D8F84",
    x"3F6D8D2D",
    x"3F6D8AD5",
    x"3F6D887D",
    x"3F6D8625",
    x"3F6D83CD",
    x"3F6D8175",
    x"3F6D7F1D",
    x"3F6D7CC4",
    x"3F6D7A6C",
    x"3F6D7813",
    x"3F6D75BA",
    x"3F6D7361",
    x"3F6D7108",
    x"3F6D6EAE",
    x"3F6D6C55",
    x"3F6D69FB",
    x"3F6D67A1",
    x"3F6D6547",
    x"3F6D62ED",
    x"3F6D6093",
    x"3F6D5E39",
    x"3F6D5BDE",
    x"3F6D5984",
    x"3F6D5729",
    x"3F6D54CE",
    x"3F6D5273",
    x"3F6D5018",
    x"3F6D4DBC",
    x"3F6D4B61",
    x"3F6D4905",
    x"3F6D46AA",
    x"3F6D444E",
    x"3F6D41F2",
    x"3F6D3F95",
    x"3F6D3D39",
    x"3F6D3ADD",
    x"3F6D3880",
    x"3F6D3623",
    x"3F6D33C6",
    x"3F6D3169",
    x"3F6D2F0C",
    x"3F6D2CAF",
    x"3F6D2A51",
    x"3F6D27F4",
    x"3F6D2596",
    x"3F6D2338",
    x"3F6D20DA",
    x"3F6D1E7C",
    x"3F6D1C1D",
    x"3F6D19BF",
    x"3F6D1760",
    x"3F6D1501",
    x"3F6D12A2",
    x"3F6D1043",
    x"3F6D0DE4",
    x"3F6D0B85",
    x"3F6D0925",
    x"3F6D06C6",
    x"3F6D0466",
    x"3F6D0206",
    x"3F6CFFA6",
    x"3F6CFD46",
    x"3F6CFAE5",
    x"3F6CF885",
    x"3F6CF624",
    x"3F6CF3C4",
    x"3F6CF163",
    x"3F6CEF02",
    x"3F6CECA0",
    x"3F6CEA3F",
    x"3F6CE7DE",
    x"3F6CE57C",
    x"3F6CE31A",
    x"3F6CE0B8",
    x"3F6CDE56",
    x"3F6CDBF4",
    x"3F6CD992",
    x"3F6CD72F",
    x"3F6CD4CD",
    x"3F6CD26A",
    x"3F6CD007",
    x"3F6CCDA4",
    x"3F6CCB41",
    x"3F6CC8DD",
    x"3F6CC67A",
    x"3F6CC416",
    x"3F6CC1B2",
    x"3F6CBF4F",
    x"3F6CBCEA",
    x"3F6CBA86",
    x"3F6CB822",
    x"3F6CB5BD",
    x"3F6CB359",
    x"3F6CB0F4",
    x"3F6CAE8F",
    x"3F6CAC2A",
    x"3F6CA9C5",
    x"3F6CA760",
    x"3F6CA4FA",
    x"3F6CA295",
    x"3F6CA02F",
    x"3F6C9DC9",
    x"3F6C9B63",
    x"3F6C98FD",
    x"3F6C9696",
    x"3F6C9430",
    x"3F6C91C9",
    x"3F6C8F62",
    x"3F6C8CFC",
    x"3F6C8A94",
    x"3F6C882D",
    x"3F6C85C6",
    x"3F6C835E",
    x"3F6C80F7",
    x"3F6C7E8F",
    x"3F6C7C27",
    x"3F6C79BF",
    x"3F6C7757",
    x"3F6C74EF",
    x"3F6C7286",
    x"3F6C701E",
    x"3F6C6DB5",
    x"3F6C6B4C",
    x"3F6C68E3",
    x"3F6C667A",
    x"3F6C6410",
    x"3F6C61A7",
    x"3F6C5F3D",
    x"3F6C5CD4",
    x"3F6C5A6A",
    x"3F6C5800",
    x"3F6C5595",
    x"3F6C532B",
    x"3F6C50C1",
    x"3F6C4E56",
    x"3F6C4BEB",
    x"3F6C4980",
    x"3F6C4715",
    x"3F6C44AA",
    x"3F6C423F",
    x"3F6C3FD3",
    x"3F6C3D68",
    x"3F6C3AFC",
    x"3F6C3890",
    x"3F6C3624",
    x"3F6C33B8",
    x"3F6C314C",
    x"3F6C2EDF",
    x"3F6C2C73",
    x"3F6C2A06",
    x"3F6C2799",
    x"3F6C252C",
    x"3F6C22BF",
    x"3F6C2051",
    x"3F6C1DE4",
    x"3F6C1B76",
    x"3F6C1909",
    x"3F6C169B",
    x"3F6C142D",
    x"3F6C11BF",
    x"3F6C0F50",
    x"3F6C0CE2",
    x"3F6C0A73",
    x"3F6C0805",
    x"3F6C0596",
    x"3F6C0327",
    x"3F6C00B7",
    x"3F6BFE48",
    x"3F6BFBD9",
    x"3F6BF969",
    x"3F6BF6F9",
    x"3F6BF48A",
    x"3F6BF21A",
    x"3F6BEFA9",
    x"3F6BED39",
    x"3F6BEAC9",
    x"3F6BE858",
    x"3F6BE5E7",
    x"3F6BE376",
    x"3F6BE105",
    x"3F6BDE94",
    x"3F6BDC23",
    x"3F6BD9B2",
    x"3F6BD740",
    x"3F6BD4CE",
    x"3F6BD25C",
    x"3F6BCFEA",
    x"3F6BCD78",
    x"3F6BCB06",
    x"3F6BC894",
    x"3F6BC621",
    x"3F6BC3AE",
    x"3F6BC13B",
    x"3F6BBEC8",
    x"3F6BBC55",
    x"3F6BB9E2",
    x"3F6BB76F",
    x"3F6BB4FB",
    x"3F6BB287",
    x"3F6BB014",
    x"3F6BADA0",
    x"3F6BAB2B",
    x"3F6BA8B7",
    x"3F6BA643",
    x"3F6BA3CE",
    x"3F6BA159",
    x"3F6B9EE5",
    x"3F6B9C70",
    x"3F6B99FB",
    x"3F6B9785",
    x"3F6B9510",
    x"3F6B929A",
    x"3F6B9025",
    x"3F6B8DAF",
    x"3F6B8B39",
    x"3F6B88C3",
    x"3F6B864C",
    x"3F6B83D6",
    x"3F6B815F",
    x"3F6B7EE9",
    x"3F6B7C72",
    x"3F6B79FB",
    x"3F6B7784",
    x"3F6B750D",
    x"3F6B7295",
    x"3F6B701E",
    x"3F6B6DA6",
    x"3F6B6B2E",
    x"3F6B68B6",
    x"3F6B663E",
    x"3F6B63C6",
    x"3F6B614D",
    x"3F6B5ED5",
    x"3F6B5C5C",
    x"3F6B59E3",
    x"3F6B576B",
    x"3F6B54F1",
    x"3F6B5278",
    x"3F6B4FFF",
    x"3F6B4D85",
    x"3F6B4B0C",
    x"3F6B4892",
    x"3F6B4618",
    x"3F6B439E",
    x"3F6B4124",
    x"3F6B3EA9",
    x"3F6B3C2F",
    x"3F6B39B4",
    x"3F6B3739",
    x"3F6B34BE",
    x"3F6B3243",
    x"3F6B2FC8",
    x"3F6B2D4D",
    x"3F6B2AD1",
    x"3F6B2855",
    x"3F6B25DA",
    x"3F6B235E",
    x"3F6B20E2",
    x"3F6B1E65",
    x"3F6B1BE9",
    x"3F6B196D",
    x"3F6B16F0",
    x"3F6B1473",
    x"3F6B11F6",
    x"3F6B0F79",
    x"3F6B0CFC",
    x"3F6B0A7F",
    x"3F6B0801",
    x"3F6B0584",
    x"3F6B0306",
    x"3F6B0088",
    x"3F6AFE0A",
    x"3F6AFB8C",
    x"3F6AF90D",
    x"3F6AF68F",
    x"3F6AF410",
    x"3F6AF191",
    x"3F6AEF12",
    x"3F6AEC93",
    x"3F6AEA14",
    x"3F6AE795",
    x"3F6AE515",
    x"3F6AE296",
    x"3F6AE016",
    x"3F6ADD96",
    x"3F6ADB16",
    x"3F6AD896",
    x"3F6AD616",
    x"3F6AD395",
    x"3F6AD115",
    x"3F6ACE94",
    x"3F6ACC13",
    x"3F6AC992",
    x"3F6AC711",
    x"3F6AC48F",
    x"3F6AC20E",
    x"3F6ABF8C",
    x"3F6ABD0B",
    x"3F6ABA89",
    x"3F6AB807",
    x"3F6AB585",
    x"3F6AB302",
    x"3F6AB080",
    x"3F6AADFD",
    x"3F6AAB7B",
    x"3F6AA8F8",
    x"3F6AA675",
    x"3F6AA3F2",
    x"3F6AA16E",
    x"3F6A9EEB",
    x"3F6A9C67",
    x"3F6A99E4",
    x"3F6A9760",
    x"3F6A94DC",
    x"3F6A9258",
    x"3F6A8FD3",
    x"3F6A8D4F",
    x"3F6A8ACA",
    x"3F6A8846",
    x"3F6A85C1",
    x"3F6A833C",
    x"3F6A80B7",
    x"3F6A7E31",
    x"3F6A7BAC",
    x"3F6A7926",
    x"3F6A76A1",
    x"3F6A741B",
    x"3F6A7195",
    x"3F6A6F0F",
    x"3F6A6C89",
    x"3F6A6A02",
    x"3F6A677C",
    x"3F6A64F5",
    x"3F6A626E",
    x"3F6A5FE7",
    x"3F6A5D60",
    x"3F6A5AD9",
    x"3F6A5851",
    x"3F6A55CA",
    x"3F6A5342",
    x"3F6A50BA",
    x"3F6A4E33",
    x"3F6A4BAA",
    x"3F6A4922",
    x"3F6A469A",
    x"3F6A4411",
    x"3F6A4189",
    x"3F6A3F00",
    x"3F6A3C77",
    x"3F6A39EE",
    x"3F6A3765",
    x"3F6A34DB",
    x"3F6A3252",
    x"3F6A2FC8",
    x"3F6A2D3E",
    x"3F6A2AB4",
    x"3F6A282A",
    x"3F6A25A0",
    x"3F6A2316",
    x"3F6A208B",
    x"3F6A1E01",
    x"3F6A1B76",
    x"3F6A18EB",
    x"3F6A1660",
    x"3F6A13D5",
    x"3F6A1149",
    x"3F6A0EBE",
    x"3F6A0C32",
    x"3F6A09A7",
    x"3F6A071B",
    x"3F6A048F",
    x"3F6A0202",
    x"3F69FF76",
    x"3F69FCEA",
    x"3F69FA5D",
    x"3F69F7D0",
    x"3F69F543",
    x"3F69F2B6",
    x"3F69F029",
    x"3F69ED9C",
    x"3F69EB0E",
    x"3F69E881",
    x"3F69E5F3",
    x"3F69E365",
    x"3F69E0D7",
    x"3F69DE49",
    x"3F69DBBB",
    x"3F69D92C",
    x"3F69D69E",
    x"3F69D40F",
    x"3F69D180",
    x"3F69CEF1",
    x"3F69CC62",
    x"3F69C9D3",
    x"3F69C743",
    x"3F69C4B4",
    x"3F69C224",
    x"3F69BF94",
    x"3F69BD04",
    x"3F69BA74",
    x"3F69B7E4",
    x"3F69B553",
    x"3F69B2C3",
    x"3F69B032",
    x"3F69ADA1",
    x"3F69AB10",
    x"3F69A87F",
    x"3F69A5EE",
    x"3F69A35D",
    x"3F69A0CB",
    x"3F699E39",
    x"3F699BA8",
    x"3F699916",
    x"3F699684",
    x"3F6993F1",
    x"3F69915F",
    x"3F698ECC",
    x"3F698C3A",
    x"3F6989A7",
    x"3F698714",
    x"3F698481",
    x"3F6981EE",
    x"3F697F5A",
    x"3F697CC7",
    x"3F697A33",
    x"3F69779F",
    x"3F69750C",
    x"3F697277",
    x"3F696FE3",
    x"3F696D4F",
    x"3F696ABA",
    x"3F696826",
    x"3F696591",
    x"3F6962FC",
    x"3F696067",
    x"3F695DD2",
    x"3F695B3D",
    x"3F6958A7",
    x"3F695611",
    x"3F69537C",
    x"3F6950E6",
    x"3F694E50",
    x"3F694BBA",
    x"3F694923",
    x"3F69468D",
    x"3F6943F6",
    x"3F694160",
    x"3F693EC9",
    x"3F693C32",
    x"3F69399A",
    x"3F693703",
    x"3F69346C",
    x"3F6931D4",
    x"3F692F3C",
    x"3F692CA5",
    x"3F692A0D",
    x"3F692774",
    x"3F6924DC",
    x"3F692244",
    x"3F691FAB",
    x"3F691D12",
    x"3F691A7A",
    x"3F6917E1",
    x"3F691547",
    x"3F6912AE",
    x"3F691015",
    x"3F690D7B",
    x"3F690AE2",
    x"3F690848",
    x"3F6905AE",
    x"3F690314",
    x"3F690079",
    x"3F68FDDF",
    x"3F68FB45",
    x"3F68F8AA",
    x"3F68F60F",
    x"3F68F374",
    x"3F68F0D9",
    x"3F68EE3E",
    x"3F68EBA2",
    x"3F68E907",
    x"3F68E66B",
    x"3F68E3CF",
    x"3F68E134",
    x"3F68DE97",
    x"3F68DBFB",
    x"3F68D95F",
    x"3F68D6C2",
    x"3F68D426",
    x"3F68D189",
    x"3F68CEEC",
    x"3F68CC4F",
    x"3F68C9B2",
    x"3F68C714",
    x"3F68C477",
    x"3F68C1D9",
    x"3F68BF3C",
    x"3F68BC9E",
    x"3F68BA00",
    x"3F68B762",
    x"3F68B4C3",
    x"3F68B225",
    x"3F68AF86",
    x"3F68ACE7",
    x"3F68AA49",
    x"3F68A7AA",
    x"3F68A50A",
    x"3F68A26B",
    x"3F689FCC",
    x"3F689D2C",
    x"3F689A8C",
    x"3F6897EC",
    x"3F68954C",
    x"3F6892AC",
    x"3F68900C",
    x"3F688D6C",
    x"3F688ACB",
    x"3F68882A",
    x"3F68858A",
    x"3F6882E9",
    x"3F688047",
    x"3F687DA6",
    x"3F687B05",
    x"3F687863",
    x"3F6875C2",
    x"3F687320",
    x"3F68707E",
    x"3F686DDC",
    x"3F686B39",
    x"3F686897",
    x"3F6865F5",
    x"3F686352",
    x"3F6860AF",
    x"3F685E0C",
    x"3F685B69",
    x"3F6858C6",
    x"3F685623",
    x"3F68537F",
    x"3F6850DB",
    x"3F684E38",
    x"3F684B94",
    x"3F6848F0",
    x"3F68464B",
    x"3F6843A7",
    x"3F684103",
    x"3F683E5E",
    x"3F683BB9",
    x"3F683914",
    x"3F68366F",
    x"3F6833CA",
    x"3F683125",
    x"3F682E7F",
    x"3F682BDA",
    x"3F682934",
    x"3F68268E",
    x"3F6823E8",
    x"3F682142",
    x"3F681E9C",
    x"3F681BF5",
    x"3F68194F",
    x"3F6816A8",
    x"3F681401",
    x"3F68115A",
    x"3F680EB3",
    x"3F680C0C",
    x"3F680964",
    x"3F6806BD",
    x"3F680415",
    x"3F68016D",
    x"3F67FEC5",
    x"3F67FC1D",
    x"3F67F975",
    x"3F67F6CC",
    x"3F67F424",
    x"3F67F17B",
    x"3F67EED2",
    x"3F67EC29",
    x"3F67E980",
    x"3F67E6D7",
    x"3F67E42E",
    x"3F67E184",
    x"3F67DEDB",
    x"3F67DC31",
    x"3F67D987",
    x"3F67D6DD",
    x"3F67D433",
    x"3F67D188",
    x"3F67CEDE",
    x"3F67CC33",
    x"3F67C988",
    x"3F67C6DE",
    x"3F67C432",
    x"3F67C187",
    x"3F67BEDC",
    x"3F67BC30",
    x"3F67B985",
    x"3F67B6D9",
    x"3F67B42D",
    x"3F67B181",
    x"3F67AED5",
    x"3F67AC29",
    x"3F67A97C",
    x"3F67A6D0",
    x"3F67A423",
    x"3F67A176",
    x"3F679EC9",
    x"3F679C1C",
    x"3F67996F",
    x"3F6796C1",
    x"3F679414",
    x"3F679166",
    x"3F678EB8",
    x"3F678C0A",
    x"3F67895C",
    x"3F6786AE",
    x"3F6783FF",
    x"3F678151",
    x"3F677EA2",
    x"3F677BF3",
    x"3F677944",
    x"3F677695",
    x"3F6773E6",
    x"3F677137",
    x"3F676E87",
    x"3F676BD8",
    x"3F676928",
    x"3F676678",
    x"3F6763C8",
    x"3F676118",
    x"3F675E67",
    x"3F675BB7",
    x"3F675906",
    x"3F675655",
    x"3F6753A5",
    x"3F6750F3",
    x"3F674E42",
    x"3F674B91",
    x"3F6748DF",
    x"3F67462E",
    x"3F67437C",
    x"3F6740CA",
    x"3F673E18",
    x"3F673B66",
    x"3F6738B4",
    x"3F673601",
    x"3F67334F",
    x"3F67309C",
    x"3F672DE9",
    x"3F672B36",
    x"3F672883",
    x"3F6725D0",
    x"3F67231C",
    x"3F672069",
    x"3F671DB5",
    x"3F671B01",
    x"3F67184D",
    x"3F671599",
    x"3F6712E5",
    x"3F671031",
    x"3F670D7C",
    x"3F670AC7",
    x"3F670813",
    x"3F67055E",
    x"3F6702A9",
    x"3F66FFF3",
    x"3F66FD3E",
    x"3F66FA88",
    x"3F66F7D3",
    x"3F66F51D",
    x"3F66F267",
    x"3F66EFB1",
    x"3F66ECFB",
    x"3F66EA45",
    x"3F66E78E",
    x"3F66E4D7",
    x"3F66E221",
    x"3F66DF6A",
    x"3F66DCB3",
    x"3F66D9FC",
    x"3F66D744",
    x"3F66D48D",
    x"3F66D1D5",
    x"3F66CF1E",
    x"3F66CC66",
    x"3F66C9AE",
    x"3F66C6F6",
    x"3F66C43D",
    x"3F66C185",
    x"3F66BECC",
    x"3F66BC14",
    x"3F66B95B",
    x"3F66B6A2",
    x"3F66B3E9",
    x"3F66B12F",
    x"3F66AE76",
    x"3F66ABBC",
    x"3F66A903",
    x"3F66A649",
    x"3F66A38F",
    x"3F66A0D5",
    x"3F669E1B",
    x"3F669B60",
    x"3F6698A6",
    x"3F6695EB",
    x"3F669330",
    x"3F669076",
    x"3F668DBA",
    x"3F668AFF",
    x"3F668844",
    x"3F668588",
    x"3F6682CD",
    x"3F668011",
    x"3F667D55",
    x"3F667A99",
    x"3F6677DD",
    x"3F667521",
    x"3F667264",
    x"3F666FA8",
    x"3F666CEB",
    x"3F666A2E",
    x"3F666771",
    x"3F6664B4",
    x"3F6661F7",
    x"3F665F39",
    x"3F665C7C",
    x"3F6659BE",
    x"3F665700",
    x"3F665442",
    x"3F665184",
    x"3F664EC6",
    x"3F664C07",
    x"3F664949",
    x"3F66468A",
    x"3F6643CB",
    x"3F66410C",
    x"3F663E4D",
    x"3F663B8E",
    x"3F6638CF",
    x"3F66360F",
    x"3F663350",
    x"3F663090",
    x"3F662DD0",
    x"3F662B10",
    x"3F662850",
    x"3F66258F",
    x"3F6622CF",
    x"3F66200E",
    x"3F661D4D",
    x"3F661A8D",
    x"3F6617CC",
    x"3F66150A",
    x"3F661249",
    x"3F660F88",
    x"3F660CC6",
    x"3F660A04",
    x"3F660742",
    x"3F660480",
    x"3F6601BE",
    x"3F65FEFC",
    x"3F65FC3A",
    x"3F65F977",
    x"3F65F6B4",
    x"3F65F3F2",
    x"3F65F12F",
    x"3F65EE6C",
    x"3F65EBA8",
    x"3F65E8E5",
    x"3F65E621",
    x"3F65E35E",
    x"3F65E09A",
    x"3F65DDD6",
    x"3F65DB12",
    x"3F65D84E",
    x"3F65D589",
    x"3F65D2C5",
    x"3F65D000",
    x"3F65CD3B",
    x"3F65CA77",
    x"3F65C7B1",
    x"3F65C4EC",
    x"3F65C227",
    x"3F65BF62",
    x"3F65BC9C",
    x"3F65B9D6",
    x"3F65B710",
    x"3F65B44A",
    x"3F65B184",
    x"3F65AEBE",
    x"3F65ABF7",
    x"3F65A931",
    x"3F65A66A",
    x"3F65A3A3",
    x"3F65A0DC",
    x"3F659E15",
    x"3F659B4E",
    x"3F659887",
    x"3F6595BF",
    x"3F6592F7",
    x"3F659030",
    x"3F658D68",
    x"3F658AA0",
    x"3F6587D7",
    x"3F65850F",
    x"3F658246",
    x"3F657F7E",
    x"3F657CB5",
    x"3F6579EC",
    x"3F657723",
    x"3F65745A",
    x"3F657190",
    x"3F656EC7",
    x"3F656BFD",
    x"3F656934",
    x"3F65666A",
    x"3F6563A0",
    x"3F6560D6",
    x"3F655E0B",
    x"3F655B41",
    x"3F655876",
    x"3F6555AC",
    x"3F6552E1",
    x"3F655016",
    x"3F654D4B",
    x"3F654A7F",
    x"3F6547B4",
    x"3F6544E8",
    x"3F65421D",
    x"3F653F51",
    x"3F653C85",
    x"3F6539B9",
    x"3F6536ED",
    x"3F653420",
    x"3F653154",
    x"3F652E87",
    x"3F652BBA",
    x"3F6528ED",
    x"3F652620",
    x"3F652353",
    x"3F652086",
    x"3F651DB8",
    x"3F651AEB",
    x"3F65181D",
    x"3F65154F",
    x"3F651281",
    x"3F650FB3",
    x"3F650CE5",
    x"3F650A16",
    x"3F650748",
    x"3F650479",
    x"3F6501AA",
    x"3F64FEDB",
    x"3F64FC0C",
    x"3F64F93D",
    x"3F64F66D",
    x"3F64F39E",
    x"3F64F0CE",
    x"3F64EDFE",
    x"3F64EB2E",
    x"3F64E85E",
    x"3F64E58E",
    x"3F64E2BD",
    x"3F64DFED",
    x"3F64DD1C",
    x"3F64DA4B",
    x"3F64D77B",
    x"3F64D4AA",
    x"3F64D1D8",
    x"3F64CF07",
    x"3F64CC35",
    x"3F64C964",
    x"3F64C692",
    x"3F64C3C0",
    x"3F64C0EE",
    x"3F64BE1C",
    x"3F64BB4A",
    x"3F64B877",
    x"3F64B5A5",
    x"3F64B2D2",
    x"3F64AFFF",
    x"3F64AD2C",
    x"3F64AA59",
    x"3F64A786",
    x"3F64A4B2",
    x"3F64A1DF",
    x"3F649F0B",
    x"3F649C37",
    x"3F649963",
    x"3F64968F",
    x"3F6493BB",
    x"3F6490E7",
    x"3F648E12",
    x"3F648B3E",
    x"3F648869",
    x"3F648594",
    x"3F6482BF",
    x"3F647FEA",
    x"3F647D14",
    x"3F647A3F",
    x"3F647769",
    x"3F647493",
    x"3F6471BE",
    x"3F646EE8",
    x"3F646C11",
    x"3F64693B",
    x"3F646665",
    x"3F64638E",
    x"3F6460B7",
    x"3F645DE1",
    x"3F645B0A",
    x"3F645832",
    x"3F64555B",
    x"3F645284",
    x"3F644FAC",
    x"3F644CD5",
    x"3F6449FD",
    x"3F644725",
    x"3F64444D",
    x"3F644174",
    x"3F643E9C",
    x"3F643BC4",
    x"3F6438EB",
    x"3F643612",
    x"3F643339",
    x"3F643060",
    x"3F642D87",
    x"3F642AAE",
    x"3F6427D4",
    x"3F6424FB",
    x"3F642221",
    x"3F641F47",
    x"3F641C6D",
    x"3F641993",
    x"3F6416B9",
    x"3F6413DE",
    x"3F641104",
    x"3F640E29",
    x"3F640B4E",
    x"3F640873",
    x"3F640598",
    x"3F6402BD",
    x"3F63FFE1",
    x"3F63FD06",
    x"3F63FA2A",
    x"3F63F74E",
    x"3F63F473",
    x"3F63F196",
    x"3F63EEBA",
    x"3F63EBDE",
    x"3F63E901",
    x"3F63E625",
    x"3F63E348",
    x"3F63E06B",
    x"3F63DD8E",
    x"3F63DAB1",
    x"3F63D7D4",
    x"3F63D4F6",
    x"3F63D219",
    x"3F63CF3B",
    x"3F63CC5D",
    x"3F63C97F",
    x"3F63C6A1",
    x"3F63C3C3",
    x"3F63C0E4",
    x"3F63BE06",
    x"3F63BB27",
    x"3F63B848",
    x"3F63B569",
    x"3F63B28A",
    x"3F63AFAB",
    x"3F63ACCC",
    x"3F63A9EC",
    x"3F63A70D",
    x"3F63A42D",
    x"3F63A14D",
    x"3F639E6D",
    x"3F639B8D",
    x"3F6398AC",
    x"3F6395CC",
    x"3F6392EB",
    x"3F63900B",
    x"3F638D2A",
    x"3F638A49",
    x"3F638767",
    x"3F638486",
    x"3F6381A5",
    x"3F637EC3",
    x"3F637BE2",
    x"3F637900",
    x"3F63761E",
    x"3F63733C",
    x"3F637059",
    x"3F636D77",
    x"3F636A95",
    x"3F6367B2",
    x"3F6364CF",
    x"3F6361EC",
    x"3F635F09",
    x"3F635C26",
    x"3F635943",
    x"3F63565F",
    x"3F63537B",
    x"3F635098",
    x"3F634DB4",
    x"3F634AD0",
    x"3F6347EC",
    x"3F634507",
    x"3F634223",
    x"3F633F3E",
    x"3F633C5A",
    x"3F633975",
    x"3F633690",
    x"3F6333AB",
    x"3F6330C5",
    x"3F632DE0",
    x"3F632AFB",
    x"3F632815",
    x"3F63252F",
    x"3F632249",
    x"3F631F63",
    x"3F631C7D",
    x"3F631996",
    x"3F6316B0",
    x"3F6313C9",
    x"3F6310E3",
    x"3F630DFC",
    x"3F630B15",
    x"3F63082E",
    x"3F630546",
    x"3F63025F",
    x"3F62FF77",
    x"3F62FC8F",
    x"3F62F9A8",
    x"3F62F6C0",
    x"3F62F3D8",
    x"3F62F0EF",
    x"3F62EE07",
    x"3F62EB1E",
    x"3F62E836",
    x"3F62E54D",
    x"3F62E264",
    x"3F62DF7B",
    x"3F62DC92",
    x"3F62D9A8",
    x"3F62D6BF",
    x"3F62D3D5",
    x"3F62D0EB",
    x"3F62CE01",
    x"3F62CB17",
    x"3F62C82D",
    x"3F62C543",
    x"3F62C258",
    x"3F62BF6E",
    x"3F62BC83",
    x"3F62B998",
    x"3F62B6AD",
    x"3F62B3C2",
    x"3F62B0D7",
    x"3F62ADEB",
    x"3F62AB00",
    x"3F62A814",
    x"3F62A528",
    x"3F62A23D",
    x"3F629F50",
    x"3F629C64",
    x"3F629978",
    x"3F62968B",
    x"3F62939F",
    x"3F6290B2",
    x"3F628DC5",
    x"3F628AD8",
    x"3F6287EB",
    x"3F6284FD",
    x"3F628210",
    x"3F627F22",
    x"3F627C35",
    x"3F627947",
    x"3F627659",
    x"3F62736B",
    x"3F62707C",
    x"3F626D8E",
    x"3F626AA0",
    x"3F6267B1",
    x"3F6264C2",
    x"3F6261D3",
    x"3F625EE4",
    x"3F625BF5",
    x"3F625905",
    x"3F625616",
    x"3F625326",
    x"3F625036",
    x"3F624D47",
    x"3F624A57",
    x"3F624766",
    x"3F624476",
    x"3F624186",
    x"3F623E95",
    x"3F623BA4",
    x"3F6238B3",
    x"3F6235C2",
    x"3F6232D1",
    x"3F622FE0",
    x"3F622CEF",
    x"3F6229FD",
    x"3F62270B",
    x"3F62241A",
    x"3F622128",
    x"3F621E35",
    x"3F621B43",
    x"3F621851",
    x"3F62155E",
    x"3F62126C",
    x"3F620F79",
    x"3F620C86",
    x"3F620993",
    x"3F6206A0",
    x"3F6203AD",
    x"3F6200B9",
    x"3F61FDC6",
    x"3F61FAD2",
    x"3F61F7DE",
    x"3F61F4EA",
    x"3F61F1F6",
    x"3F61EF02",
    x"3F61EC0D",
    x"3F61E919",
    x"3F61E624",
    x"3F61E32F",
    x"3F61E03A",
    x"3F61DD45",
    x"3F61DA50",
    x"3F61D75B",
    x"3F61D465",
    x"3F61D16F",
    x"3F61CE7A",
    x"3F61CB84",
    x"3F61C88E",
    x"3F61C598",
    x"3F61C2A1",
    x"3F61BFAB",
    x"3F61BCB4",
    x"3F61B9BE",
    x"3F61B6C7",
    x"3F61B3D0",
    x"3F61B0D9",
    x"3F61ADE1",
    x"3F61AAEA",
    x"3F61A7F2",
    x"3F61A4FB",
    x"3F61A203",
    x"3F619F0B",
    x"3F619C13",
    x"3F61991B",
    x"3F619622",
    x"3F61932A",
    x"3F619031",
    x"3F618D38",
    x"3F618A40",
    x"3F618747",
    x"3F61844D",
    x"3F618154",
    x"3F617E5B",
    x"3F617B61",
    x"3F617867",
    x"3F61756E",
    x"3F617274",
    x"3F616F79",
    x"3F616C7F",
    x"3F616985",
    x"3F61668A",
    x"3F616390",
    x"3F616095",
    x"3F615D9A",
    x"3F615A9F",
    x"3F6157A4",
    x"3F6154A8",
    x"3F6151AD",
    x"3F614EB1",
    x"3F614BB5",
    x"3F6148BA",
    x"3F6145BE",
    x"3F6142C1",
    x"3F613FC5",
    x"3F613CC9",
    x"3F6139CC",
    x"3F6136D0",
    x"3F6133D3",
    x"3F6130D6",
    x"3F612DD9",
    x"3F612ADB",
    x"3F6127DE",
    x"3F6124E1",
    x"3F6121E3",
    x"3F611EE5",
    x"3F611BE7",
    x"3F6118E9",
    x"3F6115EB",
    x"3F6112ED",
    x"3F610FEE",
    x"3F610CF0",
    x"3F6109F1",
    x"3F6106F2",
    x"3F6103F3",
    x"3F6100F4",
    x"3F60FDF5",
    x"3F60FAF5",
    x"3F60F7F6",
    x"3F60F4F6",
    x"3F60F1F6",
    x"3F60EEF6",
    x"3F60EBF6",
    x"3F60E8F6",
    x"3F60E5F6",
    x"3F60E2F5",
    x"3F60DFF4",
    x"3F60DCF4",
    x"3F60D9F3",
    x"3F60D6F2",
    x"3F60D3F1",
    x"3F60D0EF",
    x"3F60CDEE",
    x"3F60CAEC",
    x"3F60C7EB",
    x"3F60C4E9",
    x"3F60C1E7",
    x"3F60BEE5",
    x"3F60BBE2",
    x"3F60B8E0",
    x"3F60B5DE",
    x"3F60B2DB",
    x"3F60AFD8",
    x"3F60ACD5",
    x"3F60A9D2",
    x"3F60A6CF",
    x"3F60A3CC",
    x"3F60A0C8",
    x"3F609DC4",
    x"3F609AC1",
    x"3F6097BD",
    x"3F6094B9",
    x"3F6091B5",
    x"3F608EB0",
    x"3F608BAC",
    x"3F6088A7",
    x"3F6085A3",
    x"3F60829E",
    x"3F607F99",
    x"3F607C94",
    x"3F60798F",
    x"3F607689",
    x"3F607384",
    x"3F60707E",
    x"3F606D78",
    x"3F606A73",
    x"3F60676D",
    x"3F606466",
    x"3F606160",
    x"3F605E5A",
    x"3F605B53",
    x"3F60584C",
    x"3F605545",
    x"3F60523E",
    x"3F604F37",
    x"3F604C30",
    x"3F604929",
    x"3F604621",
    x"3F60431A",
    x"3F604012",
    x"3F603D0A",
    x"3F603A02",
    x"3F6036FA",
    x"3F6033F1",
    x"3F6030E9",
    x"3F602DE0",
    x"3F602AD7",
    x"3F6027CF",
    x"3F6024C6",
    x"3F6021BC",
    x"3F601EB3",
    x"3F601BAA",
    x"3F6018A0",
    x"3F601596",
    x"3F60128D",
    x"3F600F83",
    x"3F600C79",
    x"3F60096E",
    x"3F600664",
    x"3F60035A",
    x"3F60004F",
    x"3F5FFD44",
    x"3F5FFA39",
    x"3F5FF72E",
    x"3F5FF423",
    x"3F5FF118",
    x"3F5FEE0C",
    x"3F5FEB01",
    x"3F5FE7F5",
    x"3F5FE4E9",
    x"3F5FE1DD",
    x"3F5FDED1",
    x"3F5FDBC5",
    x"3F5FD8B8",
    x"3F5FD5AC",
    x"3F5FD29F",
    x"3F5FCF93",
    x"3F5FCC86",
    x"3F5FC979",
    x"3F5FC66B",
    x"3F5FC35E",
    x"3F5FC051",
    x"3F5FBD43",
    x"3F5FBA35",
    x"3F5FB727",
    x"3F5FB419",
    x"3F5FB10B",
    x"3F5FADFD",
    x"3F5FAAEF",
    x"3F5FA7E0",
    x"3F5FA4D1",
    x"3F5FA1C3",
    x"3F5F9EB4",
    x"3F5F9BA5",
    x"3F5F9895",
    x"3F5F9586",
    x"3F5F9276",
    x"3F5F8F67",
    x"3F5F8C57",
    x"3F5F8947",
    x"3F5F8637",
    x"3F5F8327",
    x"3F5F8017",
    x"3F5F7D06",
    x"3F5F79F6",
    x"3F5F76E5",
    x"3F5F73D4",
    x"3F5F70C3",
    x"3F5F6DB2",
    x"3F5F6AA1",
    x"3F5F6790",
    x"3F5F647E",
    x"3F5F616C",
    x"3F5F5E5B",
    x"3F5F5B49",
    x"3F5F5837",
    x"3F5F5525",
    x"3F5F5212",
    x"3F5F4F00",
    x"3F5F4BED",
    x"3F5F48DB",
    x"3F5F45C8",
    x"3F5F42B5",
    x"3F5F3FA2",
    x"3F5F3C8E",
    x"3F5F397B",
    x"3F5F3667",
    x"3F5F3354",
    x"3F5F3040",
    x"3F5F2D2C",
    x"3F5F2A18",
    x"3F5F2704",
    x"3F5F23EF",
    x"3F5F20DB",
    x"3F5F1DC6",
    x"3F5F1AB2",
    x"3F5F179D",
    x"3F5F1488",
    x"3F5F1173",
    x"3F5F0E5D",
    x"3F5F0B48",
    x"3F5F0833",
    x"3F5F051D",
    x"3F5F0207",
    x"3F5EFEF1",
    x"3F5EFBDB",
    x"3F5EF8C5",
    x"3F5EF5AE",
    x"3F5EF298",
    x"3F5EEF81",
    x"3F5EEC6B",
    x"3F5EE954",
    x"3F5EE63D",
    x"3F5EE326",
    x"3F5EE00E",
    x"3F5EDCF7",
    x"3F5ED9DF",
    x"3F5ED6C8",
    x"3F5ED3B0",
    x"3F5ED098",
    x"3F5ECD80",
    x"3F5ECA68",
    x"3F5EC74F",
    x"3F5EC437",
    x"3F5EC11E",
    x"3F5EBE05",
    x"3F5EBAEC",
    x"3F5EB7D3",
    x"3F5EB4BA",
    x"3F5EB1A1",
    x"3F5EAE88",
    x"3F5EAB6E",
    x"3F5EA854",
    x"3F5EA53A",
    x"3F5EA221",
    x"3F5E9F06",
    x"3F5E9BEC",
    x"3F5E98D2",
    x"3F5E95B7",
    x"3F5E929D",
    x"3F5E8F82",
    x"3F5E8C67",
    x"3F5E894C",
    x"3F5E8631",
    x"3F5E8316",
    x"3F5E7FFA",
    x"3F5E7CDE",
    x"3F5E79C3",
    x"3F5E76A7",
    x"3F5E738B",
    x"3F5E706F",
    x"3F5E6D53",
    x"3F5E6A36",
    x"3F5E671A",
    x"3F5E63FD",
    x"3F5E60E0",
    x"3F5E5DC3",
    x"3F5E5AA6",
    x"3F5E5789",
    x"3F5E546C",
    x"3F5E514E",
    x"3F5E4E31",
    x"3F5E4B13",
    x"3F5E47F5",
    x"3F5E44D7",
    x"3F5E41B9",
    x"3F5E3E9B",
    x"3F5E3B7D",
    x"3F5E385E",
    x"3F5E353F",
    x"3F5E3221",
    x"3F5E2F02",
    x"3F5E2BE3",
    x"3F5E28C3",
    x"3F5E25A4",
    x"3F5E2285",
    x"3F5E1F65",
    x"3F5E1C45",
    x"3F5E1925",
    x"3F5E1605",
    x"3F5E12E5",
    x"3F5E0FC5",
    x"3F5E0CA5",
    x"3F5E0984",
    x"3F5E0663",
    x"3F5E0343",
    x"3F5E0022",
    x"3F5DFD01",
    x"3F5DF9DF",
    x"3F5DF6BE",
    x"3F5DF39D",
    x"3F5DF07B",
    x"3F5DED59",
    x"3F5DEA37",
    x"3F5DE715",
    x"3F5DE3F3",
    x"3F5DE0D1",
    x"3F5DDDAF",
    x"3F5DDA8C",
    x"3F5DD769",
    x"3F5DD447",
    x"3F5DD124",
    x"3F5DCE01",
    x"3F5DCADD",
    x"3F5DC7BA",
    x"3F5DC497",
    x"3F5DC173",
    x"3F5DBE4F",
    x"3F5DBB2B",
    x"3F5DB807",
    x"3F5DB4E3",
    x"3F5DB1BF",
    x"3F5DAE9B",
    x"3F5DAB76",
    x"3F5DA851",
    x"3F5DA52D",
    x"3F5DA208",
    x"3F5D9EE3",
    x"3F5D9BBD",
    x"3F5D9898",
    x"3F5D9573",
    x"3F5D924D",
    x"3F5D8F27",
    x"3F5D8C01",
    x"3F5D88DB",
    x"3F5D85B5",
    x"3F5D828F",
    x"3F5D7F69",
    x"3F5D7C42",
    x"3F5D791B",
    x"3F5D75F5",
    x"3F5D72CE",
    x"3F5D6FA7",
    x"3F5D6C7F",
    x"3F5D6958",
    x"3F5D6631",
    x"3F5D6309",
    x"3F5D5FE1",
    x"3F5D5CB9",
    x"3F5D5991",
    x"3F5D5669",
    x"3F5D5341",
    x"3F5D5018",
    x"3F5D4CF0",
    x"3F5D49C7",
    x"3F5D469E",
    x"3F5D4376",
    x"3F5D404C",
    x"3F5D3D23",
    x"3F5D39FA",
    x"3F5D36D0",
    x"3F5D33A7",
    x"3F5D307D",
    x"3F5D2D53",
    x"3F5D2A29",
    x"3F5D26FF",
    x"3F5D23D5",
    x"3F5D20AA",
    x"3F5D1D80",
    x"3F5D1A55",
    x"3F5D172A",
    x"3F5D13FF",
    x"3F5D10D4",
    x"3F5D0DA9",
    x"3F5D0A7E",
    x"3F5D0752",
    x"3F5D0427",
    x"3F5D00FB",
    x"3F5CFDCF",
    x"3F5CFAA3",
    x"3F5CF777",
    x"3F5CF44B",
    x"3F5CF11E",
    x"3F5CEDF2",
    x"3F5CEAC5",
    x"3F5CE798",
    x"3F5CE46B",
    x"3F5CE13E",
    x"3F5CDE11",
    x"3F5CDAE4",
    x"3F5CD7B6",
    x"3F5CD489",
    x"3F5CD15B",
    x"3F5CCE2D",
    x"3F5CCAFF",
    x"3F5CC7D1",
    x"3F5CC4A3",
    x"3F5CC174",
    x"3F5CBE46",
    x"3F5CBB17",
    x"3F5CB7E8",
    x"3F5CB4B9",
    x"3F5CB18A",
    x"3F5CAE5B",
    x"3F5CAB2C",
    x"3F5CA7FC",
    x"3F5CA4CD",
    x"3F5CA19D",
    x"3F5C9E6D",
    x"3F5C9B3D",
    x"3F5C980D",
    x"3F5C94DD",
    x"3F5C91AC",
    x"3F5C8E7C",
    x"3F5C8B4B",
    x"3F5C881A",
    x"3F5C84EA",
    x"3F5C81B8",
    x"3F5C7E87",
    x"3F5C7B56",
    x"3F5C7824",
    x"3F5C74F3",
    x"3F5C71C1",
    x"3F5C6E8F",
    x"3F5C6B5D",
    x"3F5C682B",
    x"3F5C64F9",
    x"3F5C61C7",
    x"3F5C5E94",
    x"3F5C5B61",
    x"3F5C582F",
    x"3F5C54FC",
    x"3F5C51C9",
    x"3F5C4E95",
    x"3F5C4B62",
    x"3F5C482F",
    x"3F5C44FB",
    x"3F5C41C7",
    x"3F5C3E94",
    x"3F5C3B60",
    x"3F5C382B",
    x"3F5C34F7",
    x"3F5C31C3",
    x"3F5C2E8E",
    x"3F5C2B5A",
    x"3F5C2825",
    x"3F5C24F0",
    x"3F5C21BB",
    x"3F5C1E86",
    x"3F5C1B51",
    x"3F5C181B",
    x"3F5C14E6",
    x"3F5C11B0",
    x"3F5C0E7A",
    x"3F5C0B44",
    x"3F5C080E",
    x"3F5C04D8",
    x"3F5C01A1",
    x"3F5BFE6B",
    x"3F5BFB34",
    x"3F5BF7FD",
    x"3F5BF4C7",
    x"3F5BF190",
    x"3F5BEE58",
    x"3F5BEB21",
    x"3F5BE7EA",
    x"3F5BE4B2",
    x"3F5BE17A",
    x"3F5BDE43",
    x"3F5BDB0B",
    x"3F5BD7D3",
    x"3F5BD49A",
    x"3F5BD162",
    x"3F5BCE29",
    x"3F5BCAF1",
    x"3F5BC7B8",
    x"3F5BC47F",
    x"3F5BC146",
    x"3F5BBE0D",
    x"3F5BBAD4",
    x"3F5BB79A",
    x"3F5BB461",
    x"3F5BB127",
    x"3F5BADED",
    x"3F5BAAB3",
    x"3F5BA779",
    x"3F5BA43F",
    x"3F5BA105",
    x"3F5B9DCA",
    x"3F5B9A90",
    x"3F5B9755",
    x"3F5B941A",
    x"3F5B90DF",
    x"3F5B8DA4",
    x"3F5B8A69",
    x"3F5B872D",
    x"3F5B83F2",
    x"3F5B80B6",
    x"3F5B7D7A",
    x"3F5B7A3E",
    x"3F5B7702",
    x"3F5B73C6",
    x"3F5B708A",
    x"3F5B6D4D",
    x"3F5B6A11",
    x"3F5B66D4",
    x"3F5B6397",
    x"3F5B605A",
    x"3F5B5D1D",
    x"3F5B59E0",
    x"3F5B56A3",
    x"3F5B5365",
    x"3F5B5027",
    x"3F5B4CEA",
    x"3F5B49AC",
    x"3F5B466E",
    x"3F5B4330",
    x"3F5B3FF1",
    x"3F5B3CB3",
    x"3F5B3974",
    x"3F5B3636",
    x"3F5B32F7",
    x"3F5B2FB8",
    x"3F5B2C79",
    x"3F5B2939",
    x"3F5B25FA",
    x"3F5B22BB",
    x"3F5B1F7B",
    x"3F5B1C3B",
    x"3F5B18FB",
    x"3F5B15BB",
    x"3F5B127B",
    x"3F5B0F3B",
    x"3F5B0BFA",
    x"3F5B08BA",
    x"3F5B0579",
    x"3F5B0238",
    x"3F5AFEF7",
    x"3F5AFBB6",
    x"3F5AF875",
    x"3F5AF534",
    x"3F5AF1F2",
    x"3F5AEEB1",
    x"3F5AEB6F",
    x"3F5AE82D",
    x"3F5AE4EB",
    x"3F5AE1A9",
    x"3F5ADE67",
    x"3F5ADB24",
    x"3F5AD7E2",
    x"3F5AD49F",
    x"3F5AD15C",
    x"3F5ACE1A",
    x"3F5ACAD6",
    x"3F5AC793",
    x"3F5AC450",
    x"3F5AC10D",
    x"3F5ABDC9",
    x"3F5ABA85",
    x"3F5AB741",
    x"3F5AB3FD",
    x"3F5AB0B9",
    x"3F5AAD75",
    x"3F5AAA31",
    x"3F5AA6EC",
    x"3F5AA3A8",
    x"3F5AA063",
    x"3F5A9D1E",
    x"3F5A99D9",
    x"3F5A9694",
    x"3F5A934E",
    x"3F5A9009",
    x"3F5A8CC3",
    x"3F5A897E",
    x"3F5A8638",
    x"3F5A82F2",
    x"3F5A7FAC",
    x"3F5A7C66",
    x"3F5A791F",
    x"3F5A75D9",
    x"3F5A7292",
    x"3F5A6F4C",
    x"3F5A6C05",
    x"3F5A68BE",
    x"3F5A6577",
    x"3F5A622F",
    x"3F5A5EE8",
    x"3F5A5BA0",
    x"3F5A5859",
    x"3F5A5511",
    x"3F5A51C9",
    x"3F5A4E81",
    x"3F5A4B39",
    x"3F5A47F0",
    x"3F5A44A8",
    x"3F5A415F",
    x"3F5A3E17",
    x"3F5A3ACE",
    x"3F5A3785",
    x"3F5A343C",
    x"3F5A30F2",
    x"3F5A2DA9",
    x"3F5A2A60",
    x"3F5A2716",
    x"3F5A23CC",
    x"3F5A2082",
    x"3F5A1D38",
    x"3F5A19EE",
    x"3F5A16A4",
    x"3F5A1359",
    x"3F5A100F",
    x"3F5A0CC4",
    x"3F5A0979",
    x"3F5A062E",
    x"3F5A02E3",
    x"3F59FF98",
    x"3F59FC4D",
    x"3F59F901",
    x"3F59F5B6",
    x"3F59F26A",
    x"3F59EF1E",
    x"3F59EBD2",
    x"3F59E886",
    x"3F59E53A",
    x"3F59E1ED",
    x"3F59DEA1",
    x"3F59DB54",
    x"3F59D807",
    x"3F59D4BA",
    x"3F59D16D",
    x"3F59CE20",
    x"3F59CAD3",
    x"3F59C785",
    x"3F59C438",
    x"3F59C0EA",
    x"3F59BD9C",
    x"3F59BA4E",
    x"3F59B700",
    x"3F59B3B2",
    x"3F59B064",
    x"3F59AD15",
    x"3F59A9C7",
    x"3F59A678",
    x"3F59A329",
    x"3F599FDA",
    x"3F599C8B",
    x"3F59993C",
    x"3F5995EC",
    x"3F59929D",
    x"3F598F4D",
    x"3F598BFD",
    x"3F5988AD",
    x"3F59855D",
    x"3F59820D",
    x"3F597EBD",
    x"3F597B6C",
    x"3F59781C",
    x"3F5974CB",
    x"3F59717A",
    x"3F596E29",
    x"3F596AD8",
    x"3F596787",
    x"3F596435",
    x"3F5960E4",
    x"3F595D92",
    x"3F595A40",
    x"3F5956EE",
    x"3F59539C",
    x"3F59504A",
    x"3F594CF8",
    x"3F5949A6",
    x"3F594653",
    x"3F594300",
    x"3F593FAE",
    x"3F593C5B",
    x"3F593908",
    x"3F5935B4",
    x"3F593261",
    x"3F592F0E",
    x"3F592BBA",
    x"3F592866",
    x"3F592512",
    x"3F5921BE",
    x"3F591E6A",
    x"3F591B16",
    x"3F5917C2",
    x"3F59146D",
    x"3F591118",
    x"3F590DC4",
    x"3F590A6F",
    x"3F59071A",
    x"3F5903C5",
    x"3F59006F",
    x"3F58FD1A",
    x"3F58F9C4",
    x"3F58F66F",
    x"3F58F319",
    x"3F58EFC3",
    x"3F58EC6D",
    x"3F58E916",
    x"3F58E5C0",
    x"3F58E26A",
    x"3F58DF13",
    x"3F58DBBC",
    x"3F58D865",
    x"3F58D50E",
    x"3F58D1B7",
    x"3F58CE60",
    x"3F58CB09",
    x"3F58C7B1",
    x"3F58C45A",
    x"3F58C102",
    x"3F58BDAA",
    x"3F58BA52",
    x"3F58B6FA",
    x"3F58B3A1",
    x"3F58B049",
    x"3F58ACF0",
    x"3F58A998",
    x"3F58A63F",
    x"3F58A2E6",
    x"3F589F8D",
    x"3F589C34",
    x"3F5898DA",
    x"3F589581",
    x"3F589227",
    x"3F588ECD",
    x"3F588B74",
    x"3F58881A",
    x"3F5884BF",
    x"3F588165",
    x"3F587E0B",
    x"3F587AB0",
    x"3F587756",
    x"3F5873FB",
    x"3F5870A0",
    x"3F586D45",
    x"3F5869EA",
    x"3F58668E",
    x"3F586333",
    x"3F585FD7",
    x"3F585C7C",
    x"3F585920",
    x"3F5855C4",
    x"3F585268",
    x"3F584F0C",
    x"3F584BAF",
    x"3F584853",
    x"3F5844F6",
    x"3F584199",
    x"3F583E3D",
    x"3F583AE0",
    x"3F583782",
    x"3F583425",
    x"3F5830C8",
    x"3F582D6A",
    x"3F582A0D",
    x"3F5826AF",
    x"3F582351",
    x"3F581FF3",
    x"3F581C95",
    x"3F581936",
    x"3F5815D8",
    x"3F581279",
    x"3F580F1B",
    x"3F580BBC",
    x"3F58085D",
    x"3F5804FE",
    x"3F58019F",
    x"3F57FE3F",
    x"3F57FAE0",
    x"3F57F780",
    x"3F57F421",
    x"3F57F0C1",
    x"3F57ED61",
    x"3F57EA01",
    x"3F57E6A0",
    x"3F57E340",
    x"3F57DFDF",
    x"3F57DC7F",
    x"3F57D91E",
    x"3F57D5BD",
    x"3F57D25C",
    x"3F57CEFB",
    x"3F57CB9A",
    x"3F57C838",
    x"3F57C4D7",
    x"3F57C175",
    x"3F57BE13",
    x"3F57BAB1",
    x"3F57B74F",
    x"3F57B3ED",
    x"3F57B08B",
    x"3F57AD28",
    x"3F57A9C6",
    x"3F57A663",
    x"3F57A300",
    x"3F579F9D",
    x"3F579C3A",
    x"3F5798D7",
    x"3F579573",
    x"3F579210",
    x"3F578EAC",
    x"3F578B48",
    x"3F5787E4",
    x"3F578480",
    x"3F57811C",
    x"3F577DB8",
    x"3F577A54",
    x"3F5776EF",
    x"3F57738A",
    x"3F577026",
    x"3F576CC1",
    x"3F57695C",
    x"3F5765F6",
    x"3F576291",
    x"3F575F2C",
    x"3F575BC6",
    x"3F575860",
    x"3F5754FB",
    x"3F575195",
    x"3F574E2F",
    x"3F574AC8",
    x"3F574762",
    x"3F5743FB",
    x"3F574095",
    x"3F573D2E",
    x"3F5739C7",
    x"3F573660",
    x"3F5732F9",
    x"3F572F92",
    x"3F572C2A",
    x"3F5728C3",
    x"3F57255B",
    x"3F5721F3",
    x"3F571E8C",
    x"3F571B24",
    x"3F5717BB",
    x"3F571453",
    x"3F5710EB",
    x"3F570D82",
    x"3F570A19",
    x"3F5706B1",
    x"3F570348",
    x"3F56FFDF",
    x"3F56FC75",
    x"3F56F90C",
    x"3F56F5A3",
    x"3F56F239",
    x"3F56EECF",
    x"3F56EB65",
    x"3F56E7FB",
    x"3F56E491",
    x"3F56E127",
    x"3F56DDBD",
    x"3F56DA52",
    x"3F56D6E8",
    x"3F56D37D",
    x"3F56D012",
    x"3F56CCA7",
    x"3F56C93C",
    x"3F56C5D0",
    x"3F56C265",
    x"3F56BEF9",
    x"3F56BB8E",
    x"3F56B822",
    x"3F56B4B6",
    x"3F56B14A",
    x"3F56ADDE",
    x"3F56AA72",
    x"3F56A705",
    x"3F56A399",
    x"3F56A02C",
    x"3F569CBF",
    x"3F569952",
    x"3F5695E5",
    x"3F569278",
    x"3F568F0A",
    x"3F568B9D",
    x"3F56882F",
    x"3F5684C2",
    x"3F568154",
    x"3F567DE6",
    x"3F567A78",
    x"3F567709",
    x"3F56739B",
    x"3F56702C",
    x"3F566CBE",
    x"3F56694F",
    x"3F5665E0",
    x"3F566271",
    x"3F565F02",
    x"3F565B93",
    x"3F565823",
    x"3F5654B4",
    x"3F565144",
    x"3F564DD4",
    x"3F564A64",
    x"3F5646F4",
    x"3F564384",
    x"3F564014",
    x"3F563CA3",
    x"3F563933",
    x"3F5635C2",
    x"3F563251",
    x"3F562EE0",
    x"3F562B6F",
    x"3F5627FE",
    x"3F56248D",
    x"3F56211B",
    x"3F561DA9",
    x"3F561A38",
    x"3F5616C6",
    x"3F561354",
    x"3F560FE2",
    x"3F560C70",
    x"3F5608FD",
    x"3F56058B",
    x"3F560218",
    x"3F55FEA5",
    x"3F55FB32",
    x"3F55F7BF",
    x"3F55F44C",
    x"3F55F0D9",
    x"3F55ED65",
    x"3F55E9F2",
    x"3F55E67E",
    x"3F55E30A",
    x"3F55DF96",
    x"3F55DC22",
    x"3F55D8AE",
    x"3F55D53A",
    x"3F55D1C5",
    x"3F55CE51",
    x"3F55CADC",
    x"3F55C767",
    x"3F55C3F2",
    x"3F55C07D",
    x"3F55BD08",
    x"3F55B993",
    x"3F55B61D",
    x"3F55B2A8",
    x"3F55AF32",
    x"3F55ABBC",
    x"3F55A846",
    x"3F55A4D0",
    x"3F55A15A",
    x"3F559DE3",
    x"3F559A6D",
    x"3F5596F6",
    x"3F55937F",
    x"3F559009",
    x"3F558C92",
    x"3F55891A",
    x"3F5585A3",
    x"3F55822C",
    x"3F557EB4",
    x"3F557B3D",
    x"3F5577C5",
    x"3F55744D",
    x"3F5570D5",
    x"3F556D5D",
    x"3F5569E4",
    x"3F55666C",
    x"3F5562F3",
    x"3F555F7B",
    x"3F555C02",
    x"3F555889",
    x"3F555510",
    x"3F555197",
    x"3F554E1D",
    x"3F554AA4",
    x"3F55472A",
    x"3F5543B1",
    x"3F554037",
    x"3F553CBD",
    x"3F553943",
    x"3F5535C8",
    x"3F55324E",
    x"3F552ED4",
    x"3F552B59",
    x"3F5527DE",
    x"3F552463",
    x"3F5520E8",
    x"3F551D6D",
    x"3F5519F2",
    x"3F551676",
    x"3F5512FB",
    x"3F550F7F",
    x"3F550C04",
    x"3F550888",
    x"3F55050C",
    x"3F55018F",
    x"3F54FE13",
    x"3F54FA97",
    x"3F54F71A",
    x"3F54F39E",
    x"3F54F021",
    x"3F54ECA4",
    x"3F54E927",
    x"3F54E5AA",
    x"3F54E22C",
    x"3F54DEAF",
    x"3F54DB31",
    x"3F54D7B4",
    x"3F54D436",
    x"3F54D0B8",
    x"3F54CD3A",
    x"3F54C9BC",
    x"3F54C63D",
    x"3F54C2BF",
    x"3F54BF40",
    x"3F54BBC1",
    x"3F54B843",
    x"3F54B4C4",
    x"3F54B144",
    x"3F54ADC5",
    x"3F54AA46",
    x"3F54A6C6",
    x"3F54A347",
    x"3F549FC7",
    x"3F549C47",
    x"3F5498C7",
    x"3F549547",
    x"3F5491C7",
    x"3F548E46",
    x"3F548AC6",
    x"3F548745",
    x"3F5483C4",
    x"3F548044",
    x"3F547CC3",
    x"3F547941",
    x"3F5475C0",
    x"3F54723F",
    x"3F546EBD",
    x"3F546B3B",
    x"3F5467BA",
    x"3F546438",
    x"3F5460B6",
    x"3F545D33",
    x"3F5459B1",
    x"3F54562F",
    x"3F5452AC",
    x"3F544F2A",
    x"3F544BA7",
    x"3F544824",
    x"3F5444A1",
    x"3F54411D",
    x"3F543D9A",
    x"3F543A17",
    x"3F543693",
    x"3F54330F",
    x"3F542F8C",
    x"3F542C08",
    x"3F542883",
    x"3F5424FF",
    x"3F54217B",
    x"3F541DF6",
    x"3F541A72",
    x"3F5416ED",
    x"3F541368",
    x"3F540FE3",
    x"3F540C5E",
    x"3F5408D9",
    x"3F540553",
    x"3F5401CE",
    x"3F53FE48",
    x"3F53FAC3",
    x"3F53F73D",
    x"3F53F3B7",
    x"3F53F031",
    x"3F53ECAA",
    x"3F53E924",
    x"3F53E59D",
    x"3F53E217",
    x"3F53DE90",
    x"3F53DB09",
    x"3F53D782",
    x"3F53D3FB",
    x"3F53D074",
    x"3F53CCEC",
    x"3F53C965",
    x"3F53C5DD",
    x"3F53C255",
    x"3F53BECD",
    x"3F53BB45",
    x"3F53B7BD",
    x"3F53B435",
    x"3F53B0AC",
    x"3F53AD24",
    x"3F53A99B",
    x"3F53A612",
    x"3F53A289",
    x"3F539F00",
    x"3F539B77",
    x"3F5397EE",
    x"3F539464",
    x"3F5390DB",
    x"3F538D51",
    x"3F5389C7",
    x"3F53863D",
    x"3F5382B3",
    x"3F537F29",
    x"3F537B9E",
    x"3F537814",
    x"3F537489",
    x"3F5370FF",
    x"3F536D74",
    x"3F5369E9",
    x"3F53665E",
    x"3F5362D2",
    x"3F535F47",
    x"3F535BBB",
    x"3F535830",
    x"3F5354A4",
    x"3F535118",
    x"3F534D8C",
    x"3F534A00",
    x"3F534674",
    x"3F5342E7",
    x"3F533F5B",
    x"3F533BCE",
    x"3F533841",
    x"3F5334B5",
    x"3F533128",
    x"3F532D9A",
    x"3F532A0D",
    x"3F532680",
    x"3F5322F2",
    x"3F531F65",
    x"3F531BD7",
    x"3F531849",
    x"3F5314BB",
    x"3F53112D",
    x"3F530D9E",
    x"3F530A10",
    x"3F530681",
    x"3F5302F3",
    x"3F52FF64",
    x"3F52FBD5",
    x"3F52F846",
    x"3F52F4B7",
    x"3F52F127",
    x"3F52ED98",
    x"3F52EA08",
    x"3F52E679",
    x"3F52E2E9",
    x"3F52DF59",
    x"3F52DBC9",
    x"3F52D839",
    x"3F52D4A8",
    x"3F52D118",
    x"3F52CD87",
    x"3F52C9F7",
    x"3F52C666",
    x"3F52C2D5",
    x"3F52BF44",
    x"3F52BBB2",
    x"3F52B821",
    x"3F52B490",
    x"3F52B0FE",
    x"3F52AD6C",
    x"3F52A9DA",
    x"3F52A649",
    x"3F52A2B6",
    x"3F529F24",
    x"3F529B92",
    x"3F5297FF",
    x"3F52946D",
    x"3F5290DA",
    x"3F528D47",
    x"3F5289B4",
    x"3F528621",
    x"3F52828E",
    x"3F527EFA",
    x"3F527B67",
    x"3F5277D3",
    x"3F52743F",
    x"3F5270AC",
    x"3F526D18",
    x"3F526983",
    x"3F5265EF",
    x"3F52625B",
    x"3F525EC6",
    x"3F525B32",
    x"3F52579D",
    x"3F525408",
    x"3F525073",
    x"3F524CDE",
    x"3F524949",
    x"3F5245B3",
    x"3F52421E",
    x"3F523E88",
    x"3F523AF2",
    x"3F52375C",
    x"3F5233C6",
    x"3F523030",
    x"3F522C9A",
    x"3F522903",
    x"3F52256D",
    x"3F5221D6",
    x"3F521E3F",
    x"3F521AA8",
    x"3F521711",
    x"3F52137A",
    x"3F520FE3",
    x"3F520C4C",
    x"3F5208B4",
    x"3F52051C",
    x"3F520184",
    x"3F51FDED",
    x"3F51FA54",
    x"3F51F6BC",
    x"3F51F324",
    x"3F51EF8C",
    x"3F51EBF3",
    x"3F51E85A",
    x"3F51E4C1",
    x"3F51E129",
    x"3F51DD8F",
    x"3F51D9F6",
    x"3F51D65D",
    x"3F51D2C3",
    x"3F51CF2A",
    x"3F51CB90",
    x"3F51C7F6",
    x"3F51C45C",
    x"3F51C0C2",
    x"3F51BD28",
    x"3F51B98E",
    x"3F51B5F3",
    x"3F51B259",
    x"3F51AEBE",
    x"3F51AB23",
    x"3F51A788",
    x"3F51A3ED",
    x"3F51A052",
    x"3F519CB7",
    x"3F51991B",
    x"3F51957F",
    x"3F5191E4",
    x"3F518E48",
    x"3F518AAC",
    x"3F518710",
    x"3F518374",
    x"3F517FD7",
    x"3F517C3B",
    x"3F51789E",
    x"3F517501",
    x"3F517165",
    x"3F516DC8",
    x"3F516A2A",
    x"3F51668D",
    x"3F5162F0",
    x"3F515F52",
    x"3F515BB5",
    x"3F515817",
    x"3F515479",
    x"3F5150DB",
    x"3F514D3D",
    x"3F51499F",
    x"3F514600",
    x"3F514262",
    x"3F513EC3",
    x"3F513B25",
    x"3F513786",
    x"3F5133E7",
    x"3F513047",
    x"3F512CA8",
    x"3F512909",
    x"3F512569",
    x"3F5121CA",
    x"3F511E2A",
    x"3F511A8A",
    x"3F5116EA",
    x"3F51134A",
    x"3F510FAA",
    x"3F510C09",
    x"3F510869",
    x"3F5104C8",
    x"3F510127",
    x"3F50FD86",
    x"3F50F9E5",
    x"3F50F644",
    x"3F50F2A3",
    x"3F50EF02",
    x"3F50EB60",
    x"3F50E7BE",
    x"3F50E41D",
    x"3F50E07B",
    x"3F50DCD9",
    x"3F50D937",
    x"3F50D594",
    x"3F50D1F2",
    x"3F50CE4F",
    x"3F50CAAD",
    x"3F50C70A",
    x"3F50C367",
    x"3F50BFC4",
    x"3F50BC21",
    x"3F50B87E",
    x"3F50B4DA",
    x"3F50B137",
    x"3F50AD93",
    x"3F50A9EF",
    x"3F50A64B",
    x"3F50A2A7",
    x"3F509F03",
    x"3F509B5F",
    x"3F5097BA",
    x"3F509416",
    x"3F509071",
    x"3F508CCC",
    x"3F508927",
    x"3F508582",
    x"3F5081DD",
    x"3F507E38",
    x"3F507A92",
    x"3F5076ED",
    x"3F507347",
    x"3F506FA1",
    x"3F506BFC",
    x"3F506856",
    x"3F5064AF",
    x"3F506109",
    x"3F505D63",
    x"3F5059BC",
    x"3F505615",
    x"3F50526F",
    x"3F504EC8",
    x"3F504B21",
    x"3F504779",
    x"3F5043D2",
    x"3F50402B",
    x"3F503C83",
    x"3F5038DB",
    x"3F503534",
    x"3F50318C",
    x"3F502DE4",
    x"3F502A3B",
    x"3F502693",
    x"3F5022EB",
    x"3F501F42",
    x"3F501B9A",
    x"3F5017F1",
    x"3F501448",
    x"3F50109F",
    x"3F500CF6",
    x"3F50094C",
    x"3F5005A3",
    x"3F5001F9",
    x"3F4FFE50",
    x"3F4FFAA6",
    x"3F4FF6FC",
    x"3F4FF352",
    x"3F4FEFA8",
    x"3F4FEBFD",
    x"3F4FE853",
    x"3F4FE4A8",
    x"3F4FE0FE",
    x"3F4FDD53",
    x"3F4FD9A8",
    x"3F4FD5FD",
    x"3F4FD252",
    x"3F4FCEA6",
    x"3F4FCAFB",
    x"3F4FC74F",
    x"3F4FC3A4",
    x"3F4FBFF8",
    x"3F4FBC4C",
    x"3F4FB8A0",
    x"3F4FB4F4",
    x"3F4FB147",
    x"3F4FAD9B",
    x"3F4FA9EE",
    x"3F4FA642",
    x"3F4FA295",
    x"3F4F9EE8",
    x"3F4F9B3B",
    x"3F4F978D",
    x"3F4F93E0",
    x"3F4F9033",
    x"3F4F8C85",
    x"3F4F88D7",
    x"3F4F852A",
    x"3F4F817C",
    x"3F4F7DCE",
    x"3F4F7A1F",
    x"3F4F7671",
    x"3F4F72C3",
    x"3F4F6F14",
    x"3F4F6B65",
    x"3F4F67B7",
    x"3F4F6408",
    x"3F4F6059",
    x"3F4F5CA9",
    x"3F4F58FA",
    x"3F4F554B",
    x"3F4F519B",
    x"3F4F4DEB",
    x"3F4F4A3C",
    x"3F4F468C",
    x"3F4F42DC",
    x"3F4F3F2B",
    x"3F4F3B7B",
    x"3F4F37CB",
    x"3F4F341A",
    x"3F4F3069",
    x"3F4F2CB9",
    x"3F4F2908",
    x"3F4F2557",
    x"3F4F21A5",
    x"3F4F1DF4",
    x"3F4F1A43",
    x"3F4F1691",
    x"3F4F12DF",
    x"3F4F0F2E",
    x"3F4F0B7C",
    x"3F4F07CA",
    x"3F4F0417",
    x"3F4F0065",
    x"3F4EFCB3",
    x"3F4EF900",
    x"3F4EF54D",
    x"3F4EF19B",
    x"3F4EEDE8",
    x"3F4EEA35",
    x"3F4EE681",
    x"3F4EE2CE",
    x"3F4EDF1B",
    x"3F4EDB67",
    x"3F4ED7B3",
    x"3F4ED400",
    x"3F4ED04C",
    x"3F4ECC98",
    x"3F4EC8E4",
    x"3F4EC52F",
    x"3F4EC17B",
    x"3F4EBDC6",
    x"3F4EBA12",
    x"3F4EB65D",
    x"3F4EB2A8",
    x"3F4EAEF3",
    x"3F4EAB3E",
    x"3F4EA788",
    x"3F4EA3D3",
    x"3F4EA01D",
    x"3F4E9C68",
    x"3F4E98B2",
    x"3F4E94FC",
    x"3F4E9146",
    x"3F4E8D90",
    x"3F4E89D9",
    x"3F4E8623",
    x"3F4E826C",
    x"3F4E7EB6",
    x"3F4E7AFF",
    x"3F4E7748",
    x"3F4E7391",
    x"3F4E6FDA",
    x"3F4E6C23",
    x"3F4E686B",
    x"3F4E64B4",
    x"3F4E60FC",
    x"3F4E5D44",
    x"3F4E598C",
    x"3F4E55D4",
    x"3F4E521C",
    x"3F4E4E64",
    x"3F4E4AAB",
    x"3F4E46F3",
    x"3F4E433A",
    x"3F4E3F81",
    x"3F4E3BC8",
    x"3F4E380F",
    x"3F4E3456",
    x"3F4E309D",
    x"3F4E2CE4",
    x"3F4E292A",
    x"3F4E2570",
    x"3F4E21B7",
    x"3F4E1DFD",
    x"3F4E1A43",
    x"3F4E1689",
    x"3F4E12CE",
    x"3F4E0F14",
    x"3F4E0B59",
    x"3F4E079F",
    x"3F4E03E4",
    x"3F4E0029",
    x"3F4DFC6E",
    x"3F4DF8B3",
    x"3F4DF4F8",
    x"3F4DF13C",
    x"3F4DED81",
    x"3F4DE9C5",
    x"3F4DE609",
    x"3F4DE24D",
    x"3F4DDE91",
    x"3F4DDAD5",
    x"3F4DD719",
    x"3F4DD35D",
    x"3F4DCFA0",
    x"3F4DCBE3",
    x"3F4DC827",
    x"3F4DC46A",
    x"3F4DC0AD",
    x"3F4DBCF0",
    x"3F4DB932",
    x"3F4DB575",
    x"3F4DB1B8",
    x"3F4DADFA",
    x"3F4DAA3C",
    x"3F4DA67E",
    x"3F4DA2C0",
    x"3F4D9F02",
    x"3F4D9B44",
    x"3F4D9786",
    x"3F4D93C7",
    x"3F4D9009",
    x"3F4D8C4A",
    x"3F4D888B",
    x"3F4D84CC",
    x"3F4D810D",
    x"3F4D7D4E",
    x"3F4D798E",
    x"3F4D75CF",
    x"3F4D720F",
    x"3F4D6E4F",
    x"3F4D6A90",
    x"3F4D66D0",
    x"3F4D6310",
    x"3F4D5F4F",
    x"3F4D5B8F",
    x"3F4D57CE",
    x"3F4D540E",
    x"3F4D504D",
    x"3F4D4C8C",
    x"3F4D48CB",
    x"3F4D450A",
    x"3F4D4149",
    x"3F4D3D88",
    x"3F4D39C6",
    x"3F4D3605",
    x"3F4D3243",
    x"3F4D2E81",
    x"3F4D2ABF",
    x"3F4D26FD",
    x"3F4D233B",
    x"3F4D1F79",
    x"3F4D1BB6",
    x"3F4D17F4",
    x"3F4D1431",
    x"3F4D106E",
    x"3F4D0CAB",
    x"3F4D08E8",
    x"3F4D0525",
    x"3F4D0162",
    x"3F4CFD9E",
    x"3F4CF9DB",
    x"3F4CF617",
    x"3F4CF253",
    x"3F4CEE8F",
    x"3F4CEACB",
    x"3F4CE707",
    x"3F4CE343",
    x"3F4CDF7E",
    x"3F4CDBBA",
    x"3F4CD7F5",
    x"3F4CD430",
    x"3F4CD06B",
    x"3F4CCCA6",
    x"3F4CC8E1",
    x"3F4CC51C",
    x"3F4CC156",
    x"3F4CBD91",
    x"3F4CB9CB",
    x"3F4CB605",
    x"3F4CB23F",
    x"3F4CAE79",
    x"3F4CAAB3",
    x"3F4CA6ED",
    x"3F4CA327",
    x"3F4C9F60",
    x"3F4C9B99",
    x"3F4C97D3",
    x"3F4C940C",
    x"3F4C9045",
    x"3F4C8C7E",
    x"3F4C88B6",
    x"3F4C84EF",
    x"3F4C8128",
    x"3F4C7D60",
    x"3F4C7998",
    x"3F4C75D0",
    x"3F4C7208",
    x"3F4C6E40",
    x"3F4C6A78",
    x"3F4C66B0",
    x"3F4C62E7",
    x"3F4C5F1E",
    x"3F4C5B56",
    x"3F4C578D",
    x"3F4C53C4",
    x"3F4C4FFB",
    x"3F4C4C32",
    x"3F4C4868",
    x"3F4C449F",
    x"3F4C40D5",
    x"3F4C3D0B",
    x"3F4C3942",
    x"3F4C3578",
    x"3F4C31AD",
    x"3F4C2DE3",
    x"3F4C2A19",
    x"3F4C264E",
    x"3F4C2284",
    x"3F4C1EB9",
    x"3F4C1AEE",
    x"3F4C1723",
    x"3F4C1358",
    x"3F4C0F8D",
    x"3F4C0BC2",
    x"3F4C07F6",
    x"3F4C042B",
    x"3F4C005F",
    x"3F4BFC93",
    x"3F4BF8C7",
    x"3F4BF4FB",
    x"3F4BF12F",
    x"3F4BED63",
    x"3F4BE996",
    x"3F4BE5CA",
    x"3F4BE1FD",
    x"3F4BDE30",
    x"3F4BDA63",
    x"3F4BD696",
    x"3F4BD2C9",
    x"3F4BCEFC",
    x"3F4BCB2F",
    x"3F4BC761",
    x"3F4BC393",
    x"3F4BBFC6",
    x"3F4BBBF8",
    x"3F4BB82A",
    x"3F4BB45B",
    x"3F4BB08D",
    x"3F4BACBF",
    x"3F4BA8F0",
    x"3F4BA522",
    x"3F4BA153",
    x"3F4B9D84",
    x"3F4B99B5",
    x"3F4B95E6",
    x"3F4B9217",
    x"3F4B8E47",
    x"3F4B8A78",
    x"3F4B86A8",
    x"3F4B82D8",
    x"3F4B7F09",
    x"3F4B7B39",
    x"3F4B7768",
    x"3F4B7398",
    x"3F4B6FC8",
    x"3F4B6BF7",
    x"3F4B6827",
    x"3F4B6456",
    x"3F4B6085",
    x"3F4B5CB4",
    x"3F4B58E3",
    x"3F4B5512",
    x"3F4B5141",
    x"3F4B4D6F",
    x"3F4B499E",
    x"3F4B45CC",
    x"3F4B41FA",
    x"3F4B3E28",
    x"3F4B3A56",
    x"3F4B3684",
    x"3F4B32B2",
    x"3F4B2EDF",
    x"3F4B2B0D",
    x"3F4B273A",
    x"3F4B2367",
    x"3F4B1F94",
    x"3F4B1BC1",
    x"3F4B17EE",
    x"3F4B141B",
    x"3F4B1047",
    x"3F4B0C74",
    x"3F4B08A0",
    x"3F4B04CC",
    x"3F4B00F8",
    x"3F4AFD24",
    x"3F4AF950",
    x"3F4AF57C",
    x"3F4AF1A8",
    x"3F4AEDD3",
    x"3F4AE9FE",
    x"3F4AE62A",
    x"3F4AE255",
    x"3F4ADE80",
    x"3F4ADAAB",
    x"3F4AD6D5",
    x"3F4AD300",
    x"3F4ACF2A",
    x"3F4ACB55",
    x"3F4AC77F",
    x"3F4AC3A9",
    x"3F4ABFD3",
    x"3F4ABBFD",
    x"3F4AB827",
    x"3F4AB451",
    x"3F4AB07A",
    x"3F4AACA4",
    x"3F4AA8CD",
    x"3F4AA4F6",
    x"3F4AA11F",
    x"3F4A9D48",
    x"3F4A9971",
    x"3F4A9599",
    x"3F4A91C2",
    x"3F4A8DEA",
    x"3F4A8A13",
    x"3F4A863B",
    x"3F4A8263",
    x"3F4A7E8B",
    x"3F4A7AB3",
    x"3F4A76DA",
    x"3F4A7302",
    x"3F4A6F29",
    x"3F4A6B51",
    x"3F4A6778",
    x"3F4A639F",
    x"3F4A5FC6",
    x"3F4A5BED",
    x"3F4A5814",
    x"3F4A543A",
    x"3F4A5061",
    x"3F4A4C87",
    x"3F4A48AD",
    x"3F4A44D3",
    x"3F4A40F9",
    x"3F4A3D1F",
    x"3F4A3945",
    x"3F4A356B",
    x"3F4A3190",
    x"3F4A2DB6",
    x"3F4A29DB",
    x"3F4A2600",
    x"3F4A2225",
    x"3F4A1E4A",
    x"3F4A1A6F",
    x"3F4A1693",
    x"3F4A12B8",
    x"3F4A0EDC",
    x"3F4A0B01",
    x"3F4A0725",
    x"3F4A0349",
    x"3F49FF6D",
    x"3F49FB91",
    x"3F49F7B4",
    x"3F49F3D8",
    x"3F49EFFB",
    x"3F49EC1F",
    x"3F49E842",
    x"3F49E465",
    x"3F49E088",
    x"3F49DCAB",
    x"3F49D8CD",
    x"3F49D4F0",
    x"3F49D112",
    x"3F49CD35",
    x"3F49C957",
    x"3F49C579",
    x"3F49C19B",
    x"3F49BDBD",
    x"3F49B9DF",
    x"3F49B600",
    x"3F49B222",
    x"3F49AE43",
    x"3F49AA64",
    x"3F49A685",
    x"3F49A2A6",
    x"3F499EC7",
    x"3F499AE8",
    x"3F499709",
    x"3F499329",
    x"3F498F4A",
    x"3F498B6A",
    x"3F49878A",
    x"3F4983AA",
    x"3F497FCA",
    x"3F497BEA",
    x"3F497809",
    x"3F497429",
    x"3F497048",
    x"3F496C68",
    x"3F496887",
    x"3F4964A6",
    x"3F4960C5",
    x"3F495CE4",
    x"3F495902",
    x"3F495521",
    x"3F49513F",
    x"3F494D5E",
    x"3F49497C",
    x"3F49459A",
    x"3F4941B8",
    x"3F493DD6",
    x"3F4939F4",
    x"3F493611",
    x"3F49322F",
    x"3F492E4C",
    x"3F492A69",
    x"3F492686",
    x"3F4922A3",
    x"3F491EC0",
    x"3F491ADD",
    x"3F4916FA",
    x"3F491316",
    x"3F490F33",
    x"3F490B4F",
    x"3F49076B",
    x"3F490387",
    x"3F48FFA3",
    x"3F48FBBF",
    x"3F48F7DA",
    x"3F48F3F6",
    x"3F48F011",
    x"3F48EC2D",
    x"3F48E848",
    x"3F48E463",
    x"3F48E07E",
    x"3F48DC99",
    x"3F48D8B3",
    x"3F48D4CE",
    x"3F48D0E9",
    x"3F48CD03",
    x"3F48C91D",
    x"3F48C537",
    x"3F48C151",
    x"3F48BD6B",
    x"3F48B985",
    x"3F48B59E",
    x"3F48B1B8",
    x"3F48ADD1",
    x"3F48A9EA",
    x"3F48A604",
    x"3F48A21D",
    x"3F489E36",
    x"3F489A4E",
    x"3F489667",
    x"3F48927F",
    x"3F488E98",
    x"3F488AB0",
    x"3F4886C8",
    x"3F4882E0",
    x"3F487EF8",
    x"3F487B10",
    x"3F487728",
    x"3F48733F",
    x"3F486F57",
    x"3F486B6E",
    x"3F486785",
    x"3F48639C",
    x"3F485FB3",
    x"3F485BCA",
    x"3F4857E1",
    x"3F4853F7",
    x"3F48500E",
    x"3F484C24",
    x"3F48483A",
    x"3F484451",
    x"3F484067",
    x"3F483C7C",
    x"3F483892",
    x"3F4834A8",
    x"3F4830BD",
    x"3F482CD3",
    x"3F4828E8",
    x"3F4824FD",
    x"3F482112",
    x"3F481D27",
    x"3F48193C",
    x"3F481550",
    x"3F481165",
    x"3F480D79",
    x"3F48098E",
    x"3F4805A2",
    x"3F4801B6",
    x"3F47FDCA",
    x"3F47F9DE",
    x"3F47F5F1",
    x"3F47F205",
    x"3F47EE18",
    x"3F47EA2C",
    x"3F47E63F",
    x"3F47E252",
    x"3F47DE65",
    x"3F47DA78",
    x"3F47D68B",
    x"3F47D29D",
    x"3F47CEB0",
    x"3F47CAC2",
    x"3F47C6D4",
    x"3F47C2E7",
    x"3F47BEF9",
    x"3F47BB0A",
    x"3F47B71C",
    x"3F47B32E",
    x"3F47AF3F",
    x"3F47AB51",
    x"3F47A762",
    x"3F47A373",
    x"3F479F84",
    x"3F479B95",
    x"3F4797A6",
    x"3F4793B7",
    x"3F478FC7",
    x"3F478BD8",
    x"3F4787E8",
    x"3F4783F8",
    x"3F478008",
    x"3F477C18",
    x"3F477828",
    x"3F477438",
    x"3F477048",
    x"3F476C57",
    x"3F476866",
    x"3F476476",
    x"3F476085",
    x"3F475C94",
    x"3F4758A3",
    x"3F4754B2",
    x"3F4750C0",
    x"3F474CCF",
    x"3F4748DD",
    x"3F4744EB",
    x"3F4740FA",
    x"3F473D08",
    x"3F473916",
    x"3F473523",
    x"3F473131",
    x"3F472D3F",
    x"3F47294C",
    x"3F472559",
    x"3F472167",
    x"3F471D74",
    x"3F471981",
    x"3F47158D",
    x"3F47119A",
    x"3F470DA7",
    x"3F4709B3",
    x"3F4705C0",
    x"3F4701CC",
    x"3F46FDD8",
    x"3F46F9E4",
    x"3F46F5F0",
    x"3F46F1FC",
    x"3F46EE07",
    x"3F46EA13",
    x"3F46E61E",
    x"3F46E22A",
    x"3F46DE35",
    x"3F46DA40",
    x"3F46D64B",
    x"3F46D256",
    x"3F46CE60",
    x"3F46CA6B",
    x"3F46C675",
    x"3F46C280",
    x"3F46BE8A",
    x"3F46BA94",
    x"3F46B69E",
    x"3F46B2A8",
    x"3F46AEB1",
    x"3F46AABB",
    x"3F46A6C5",
    x"3F46A2CE",
    x"3F469ED7",
    x"3F469AE0",
    x"3F4696E9",
    x"3F4692F2",
    x"3F468EFB",
    x"3F468B04",
    x"3F46870C",
    x"3F468315",
    x"3F467F1D",
    x"3F467B25",
    x"3F46772D",
    x"3F467335",
    x"3F466F3D",
    x"3F466B45",
    x"3F46674C",
    x"3F466354",
    x"3F465F5B",
    x"3F465B62",
    x"3F465769",
    x"3F465370",
    x"3F464F77",
    x"3F464B7E",
    x"3F464785",
    x"3F46438B",
    x"3F463F91",
    x"3F463B98",
    x"3F46379E",
    x"3F4633A4",
    x"3F462FAA",
    x"3F462BB0",
    x"3F4627B5",
    x"3F4623BB",
    x"3F461FC0",
    x"3F461BC6",
    x"3F4617CB",
    x"3F4613D0",
    x"3F460FD5",
    x"3F460BDA",
    x"3F4607DE",
    x"3F4603E3",
    x"3F45FFE7",
    x"3F45FBEC",
    x"3F45F7F0",
    x"3F45F3F4",
    x"3F45EFF8",
    x"3F45EBFC",
    x"3F45E800",
    x"3F45E403",
    x"3F45E007",
    x"3F45DC0A",
    x"3F45D80E",
    x"3F45D411",
    x"3F45D014",
    x"3F45CC17",
    x"3F45C819",
    x"3F45C41C",
    x"3F45C01F",
    x"3F45BC21",
    x"3F45B824",
    x"3F45B426",
    x"3F45B028",
    x"3F45AC2A",
    x"3F45A82C",
    x"3F45A42D",
    x"3F45A02F",
    x"3F459C31",
    x"3F459832",
    x"3F459433",
    x"3F459034",
    x"3F458C35",
    x"3F458836",
    x"3F458437",
    x"3F458038",
    x"3F457C38",
    x"3F457839",
    x"3F457439",
    x"3F457039",
    x"3F456C39",
    x"3F456839",
    x"3F456439",
    x"3F456039",
    x"3F455C38",
    x"3F455838",
    x"3F455437",
    x"3F455036",
    x"3F454C35",
    x"3F454834",
    x"3F454433",
    x"3F454032",
    x"3F453C31",
    x"3F45382F",
    x"3F45342E",
    x"3F45302C",
    x"3F452C2A",
    x"3F452828",
    x"3F452426",
    x"3F452024",
    x"3F451C22",
    x"3F45181F",
    x"3F45141D",
    x"3F45101A",
    x"3F450C17",
    x"3F450814",
    x"3F450411",
    x"3F45000E",
    x"3F44FC0B",
    x"3F44F807",
    x"3F44F404",
    x"3F44F000",
    x"3F44EBFD",
    x"3F44E7F9",
    x"3F44E3F5",
    x"3F44DFF1",
    x"3F44DBED",
    x"3F44D7E8",
    x"3F44D3E4",
    x"3F44CFDF",
    x"3F44CBDB",
    x"3F44C7D6",
    x"3F44C3D1",
    x"3F44BFCC",
    x"3F44BBC7",
    x"3F44B7C1",
    x"3F44B3BC",
    x"3F44AFB6",
    x"3F44ABB1",
    x"3F44A7AB",
    x"3F44A3A5",
    x"3F449F9F",
    x"3F449B99",
    x"3F449793",
    x"3F44938D",
    x"3F448F86",
    x"3F448B80",
    x"3F448779",
    x"3F448372",
    x"3F447F6B",
    x"3F447B64",
    x"3F44775D",
    x"3F447356",
    x"3F446F4E",
    x"3F446B47",
    x"3F44673F",
    x"3F446337",
    x"3F445F2F",
    x"3F445B27",
    x"3F44571F",
    x"3F445317",
    x"3F444F0F",
    x"3F444B06",
    x"3F4446FE",
    x"3F4442F5",
    x"3F443EEC",
    x"3F443AE3",
    x"3F4436DA",
    x"3F4432D1",
    x"3F442EC8",
    x"3F442ABE",
    x"3F4426B5",
    x"3F4422AB",
    x"3F441EA1",
    x"3F441A97",
    x"3F44168D",
    x"3F441283",
    x"3F440E79",
    x"3F440A6F",
    x"3F440664",
    x"3F44025A",
    x"3F43FE4F",
    x"3F43FA44",
    x"3F43F639",
    x"3F43F22E",
    x"3F43EE23",
    x"3F43EA17",
    x"3F43E60C",
    x"3F43E200",
    x"3F43DDF5",
    x"3F43D9E9",
    x"3F43D5DD",
    x"3F43D1D1",
    x"3F43CDC5",
    x"3F43C9B9",
    x"3F43C5AC",
    x"3F43C1A0",
    x"3F43BD93",
    x"3F43B987",
    x"3F43B57A",
    x"3F43B16D",
    x"3F43AD60",
    x"3F43A953",
    x"3F43A545",
    x"3F43A138",
    x"3F439D2A",
    x"3F43991D",
    x"3F43950F",
    x"3F439101",
    x"3F438CF3",
    x"3F4388E5",
    x"3F4384D6",
    x"3F4380C8",
    x"3F437CBA",
    x"3F4378AB",
    x"3F43749C",
    x"3F43708D",
    x"3F436C7F",
    x"3F43686F",
    x"3F436460",
    x"3F436051",
    x"3F435C41",
    x"3F435832",
    x"3F435422",
    x"3F435012",
    x"3F434C03",
    x"3F4347F3",
    x"3F4343E2",
    x"3F433FD2",
    x"3F433BC2",
    x"3F4337B1",
    x"3F4333A1",
    x"3F432F90",
    x"3F432B7F",
    x"3F43276E",
    x"3F43235D",
    x"3F431F4C",
    x"3F431B3B",
    x"3F431729",
    x"3F431318",
    x"3F430F06",
    x"3F430AF4",
    x"3F4306E2",
    x"3F4302D0",
    x"3F42FEBE",
    x"3F42FAAC",
    x"3F42F69A",
    x"3F42F287",
    x"3F42EE74",
    x"3F42EA62",
    x"3F42E64F",
    x"3F42E23C",
    x"3F42DE29",
    x"3F42DA16",
    x"3F42D602",
    x"3F42D1EF",
    x"3F42CDDB",
    x"3F42C9C8",
    x"3F42C5B4",
    x"3F42C1A0",
    x"3F42BD8C",
    x"3F42B978",
    x"3F42B564",
    x"3F42B14F",
    x"3F42AD3B",
    x"3F42A926",
    x"3F42A511",
    x"3F42A0FD",
    x"3F429CE8",
    x"3F4298D3",
    x"3F4294BD",
    x"3F4290A8",
    x"3F428C93",
    x"3F42887D",
    x"3F428468",
    x"3F428052",
    x"3F427C3C",
    x"3F427826",
    x"3F427410",
    x"3F426FFA",
    x"3F426BE3",
    x"3F4267CD",
    x"3F4263B6",
    x"3F425F9F",
    x"3F425B89",
    x"3F425772",
    x"3F42535B",
    x"3F424F43",
    x"3F424B2C",
    x"3F424715",
    x"3F4242FD",
    x"3F423EE5",
    x"3F423ACE",
    x"3F4236B6",
    x"3F42329E",
    x"3F422E86",
    x"3F422A6E",
    x"3F422655",
    x"3F42223D",
    x"3F421E24",
    x"3F421A0B",
    x"3F4215F3",
    x"3F4211DA",
    x"3F420DC1",
    x"3F4209A7",
    x"3F42058E",
    x"3F420175",
    x"3F41FD5B",
    x"3F41F942",
    x"3F41F528",
    x"3F41F10E",
    x"3F41ECF4",
    x"3F41E8DA",
    x"3F41E4C0",
    x"3F41E0A5",
    x"3F41DC8B",
    x"3F41D870",
    x"3F41D456",
    x"3F41D03B",
    x"3F41CC20",
    x"3F41C805",
    x"3F41C3EA",
    x"3F41BFCF",
    x"3F41BBB3",
    x"3F41B798",
    x"3F41B37C",
    x"3F41AF60",
    x"3F41AB44",
    x"3F41A728",
    x"3F41A30C",
    x"3F419EF0",
    x"3F419AD4",
    x"3F4196B7",
    x"3F41929B",
    x"3F418E7E",
    x"3F418A61",
    x"3F418645",
    x"3F418228",
    x"3F417E0A",
    x"3F4179ED",
    x"3F4175D0",
    x"3F4171B2",
    x"3F416D95",
    x"3F416977",
    x"3F416559",
    x"3F41613B",
    x"3F415D1D",
    x"3F4158FF",
    x"3F4154E1",
    x"3F4150C2",
    x"3F414CA4",
    x"3F414885",
    x"3F414466",
    x"3F414047",
    x"3F413C28",
    x"3F413809",
    x"3F4133EA",
    x"3F412FCB",
    x"3F412BAB",
    x"3F41278C",
    x"3F41236C",
    x"3F411F4C",
    x"3F411B2C",
    x"3F41170C",
    x"3F4112EC",
    x"3F410ECC",
    x"3F410AAB",
    x"3F41068B",
    x"3F41026A",
    x"3F40FE49",
    x"3F40FA29",
    x"3F40F608",
    x"3F40F1E7",
    x"3F40EDC5",
    x"3F40E9A4",
    x"3F40E583",
    x"3F40E161",
    x"3F40DD3F",
    x"3F40D91E",
    x"3F40D4FC",
    x"3F40D0DA",
    x"3F40CCB7",
    x"3F40C895",
    x"3F40C473",
    x"3F40C050",
    x"3F40BC2E",
    x"3F40B80B",
    x"3F40B3E8",
    x"3F40AFC5",
    x"3F40ABA2",
    x"3F40A77F",
    x"3F40A35C",
    x"3F409F38",
    x"3F409B15",
    x"3F4096F1",
    x"3F4092CD",
    x"3F408EA9",
    x"3F408A85",
    x"3F408661",
    x"3F40823D",
    x"3F407E19",
    x"3F4079F4",
    x"3F4075D0",
    x"3F4071AB",
    x"3F406D86",
    x"3F406961",
    x"3F40653C",
    x"3F406117",
    x"3F405CF2",
    x"3F4058CD",
    x"3F4054A7",
    x"3F405081",
    x"3F404C5C",
    x"3F404836",
    x"3F404410",
    x"3F403FEA",
    x"3F403BC4",
    x"3F40379D",
    x"3F403377",
    x"3F402F50",
    x"3F402B2A",
    x"3F402703",
    x"3F4022DC",
    x"3F401EB5",
    x"3F401A8E",
    x"3F401667",
    x"3F40123F",
    x"3F400E18",
    x"3F4009F0",
    x"3F4005C8",
    x"3F4001A1",
    x"3F3FFD79",
    x"3F3FF951",
    x"3F3FF529",
    x"3F3FF100",
    x"3F3FECD8",
    x"3F3FE8AF",
    x"3F3FE487",
    x"3F3FE05E",
    x"3F3FDC35",
    x"3F3FD80C",
    x"3F3FD3E3",
    x"3F3FCFBA",
    x"3F3FCB91",
    x"3F3FC767",
    x"3F3FC33E",
    x"3F3FBF14",
    x"3F3FBAEA",
    x"3F3FB6C0",
    x"3F3FB296",
    x"3F3FAE6C",
    x"3F3FAA42",
    x"3F3FA617",
    x"3F3FA1ED",
    x"3F3F9DC2",
    x"3F3F9998",
    x"3F3F956D",
    x"3F3F9142",
    x"3F3F8D17",
    x"3F3F88EC",
    x"3F3F84C0",
    x"3F3F8095",
    x"3F3F7C6A",
    x"3F3F783E",
    x"3F3F7412",
    x"3F3F6FE6",
    x"3F3F6BBA",
    x"3F3F678E",
    x"3F3F6362",
    x"3F3F5F36",
    x"3F3F5B09",
    x"3F3F56DD",
    x"3F3F52B0",
    x"3F3F4E83",
    x"3F3F4A56",
    x"3F3F4629",
    x"3F3F41FC",
    x"3F3F3DCF",
    x"3F3F39A2",
    x"3F3F3574",
    x"3F3F3147",
    x"3F3F2D19",
    x"3F3F28EB",
    x"3F3F24BD",
    x"3F3F208F",
    x"3F3F1C61",
    x"3F3F1833",
    x"3F3F1404",
    x"3F3F0FD6",
    x"3F3F0BA7",
    x"3F3F0778",
    x"3F3F034A",
    x"3F3EFF1B",
    x"3F3EFAEB",
    x"3F3EF6BC",
    x"3F3EF28D",
    x"3F3EEE5E",
    x"3F3EEA2E",
    x"3F3EE5FE",
    x"3F3EE1CF",
    x"3F3EDD9F",
    x"3F3ED96F",
    x"3F3ED53F",
    x"3F3ED10E",
    x"3F3ECCDE",
    x"3F3EC8AD",
    x"3F3EC47D",
    x"3F3EC04C",
    x"3F3EBC1B",
    x"3F3EB7EA",
    x"3F3EB3B9",
    x"3F3EAF88",
    x"3F3EAB57",
    x"3F3EA726",
    x"3F3EA2F4",
    x"3F3E9EC3",
    x"3F3E9A91",
    x"3F3E965F",
    x"3F3E922D",
    x"3F3E8DFB",
    x"3F3E89C9",
    x"3F3E8596",
    x"3F3E8164",
    x"3F3E7D31",
    x"3F3E78FF",
    x"3F3E74CC",
    x"3F3E7099",
    x"3F3E6C66",
    x"3F3E6833",
    x"3F3E6400",
    x"3F3E5FCD",
    x"3F3E5B99",
    x"3F3E5766",
    x"3F3E5332",
    x"3F3E4EFE",
    x"3F3E4ACA",
    x"3F3E4696",
    x"3F3E4262",
    x"3F3E3E2E",
    x"3F3E39F9",
    x"3F3E35C5",
    x"3F3E3190",
    x"3F3E2D5C",
    x"3F3E2927",
    x"3F3E24F2",
    x"3F3E20BD",
    x"3F3E1C88",
    x"3F3E1852",
    x"3F3E141D",
    x"3F3E0FE7",
    x"3F3E0BB2",
    x"3F3E077C",
    x"3F3E0346",
    x"3F3DFF10",
    x"3F3DFADA",
    x"3F3DF6A4",
    x"3F3DF26E",
    x"3F3DEE37",
    x"3F3DEA01",
    x"3F3DE5CA",
    x"3F3DE193",
    x"3F3DDD5C",
    x"3F3DD925",
    x"3F3DD4EE",
    x"3F3DD0B7",
    x"3F3DCC80",
    x"3F3DC848",
    x"3F3DC411",
    x"3F3DBFD9",
    x"3F3DBBA1",
    x"3F3DB769",
    x"3F3DB331",
    x"3F3DAEF9",
    x"3F3DAAC1",
    x"3F3DA688",
    x"3F3DA250",
    x"3F3D9E17",
    x"3F3D99DF",
    x"3F3D95A6",
    x"3F3D916D",
    x"3F3D8D34",
    x"3F3D88FB",
    x"3F3D84C1",
    x"3F3D8088",
    x"3F3D7C4E",
    x"3F3D7815",
    x"3F3D73DB",
    x"3F3D6FA1",
    x"3F3D6B67",
    x"3F3D672D",
    x"3F3D62F3",
    x"3F3D5EB9",
    x"3F3D5A7E",
    x"3F3D5644",
    x"3F3D5209",
    x"3F3D4DCE",
    x"3F3D4993",
    x"3F3D4558",
    x"3F3D411D",
    x"3F3D3CE2",
    x"3F3D38A7",
    x"3F3D346B",
    x"3F3D3030",
    x"3F3D2BF4",
    x"3F3D27B8",
    x"3F3D237C",
    x"3F3D1F40",
    x"3F3D1B04",
    x"3F3D16C8",
    x"3F3D128C",
    x"3F3D0E4F",
    x"3F3D0A12",
    x"3F3D05D6",
    x"3F3D0199",
    x"3F3CFD5C",
    x"3F3CF91F",
    x"3F3CF4E2",
    x"3F3CF0A5",
    x"3F3CEC67",
    x"3F3CE82A",
    x"3F3CE3EC",
    x"3F3CDFAE",
    x"3F3CDB70",
    x"3F3CD733",
    x"3F3CD2F4",
    x"3F3CCEB6",
    x"3F3CCA78",
    x"3F3CC63A",
    x"3F3CC1FB",
    x"3F3CBDBC",
    x"3F3CB97E",
    x"3F3CB53F",
    x"3F3CB100",
    x"3F3CACC1",
    x"3F3CA881",
    x"3F3CA442",
    x"3F3CA003",
    x"3F3C9BC3",
    x"3F3C9784",
    x"3F3C9344",
    x"3F3C8F04",
    x"3F3C8AC4",
    x"3F3C8684",
    x"3F3C8244",
    x"3F3C7E03",
    x"3F3C79C3",
    x"3F3C7582",
    x"3F3C7141",
    x"3F3C6D01",
    x"3F3C68C0",
    x"3F3C647F",
    x"3F3C603E",
    x"3F3C5BFC",
    x"3F3C57BB",
    x"3F3C5379",
    x"3F3C4F38",
    x"3F3C4AF6",
    x"3F3C46B4",
    x"3F3C4272",
    x"3F3C3E30",
    x"3F3C39EE",
    x"3F3C35AC",
    x"3F3C316A",
    x"3F3C2D27",
    x"3F3C28E4",
    x"3F3C24A2",
    x"3F3C205F",
    x"3F3C1C1C",
    x"3F3C17D9",
    x"3F3C1396",
    x"3F3C0F52",
    x"3F3C0B0F",
    x"3F3C06CB",
    x"3F3C0288",
    x"3F3BFE44",
    x"3F3BFA00",
    x"3F3BF5BC",
    x"3F3BF178",
    x"3F3BED34",
    x"3F3BE8F0",
    x"3F3BE4AB",
    x"3F3BE067",
    x"3F3BDC22",
    x"3F3BD7DD",
    x"3F3BD398",
    x"3F3BCF53",
    x"3F3BCB0E",
    x"3F3BC6C9",
    x"3F3BC284",
    x"3F3BBE3E",
    x"3F3BB9F9",
    x"3F3BB5B3",
    x"3F3BB16D",
    x"3F3BAD27",
    x"3F3BA8E1",
    x"3F3BA49B",
    x"3F3BA055",
    x"3F3B9C0F",
    x"3F3B97C8",
    x"3F3B9382",
    x"3F3B8F3B",
    x"3F3B8AF4",
    x"3F3B86AD",
    x"3F3B8266",
    x"3F3B7E1F",
    x"3F3B79D8",
    x"3F3B7590",
    x"3F3B7149",
    x"3F3B6D01",
    x"3F3B68BA",
    x"3F3B6472",
    x"3F3B602A",
    x"3F3B5BE2",
    x"3F3B579A",
    x"3F3B5351",
    x"3F3B4F09",
    x"3F3B4AC1",
    x"3F3B4678",
    x"3F3B422F",
    x"3F3B3DE6",
    x"3F3B399E",
    x"3F3B3554",
    x"3F3B310B",
    x"3F3B2CC2",
    x"3F3B2879",
    x"3F3B242F",
    x"3F3B1FE5",
    x"3F3B1B9C",
    x"3F3B1752",
    x"3F3B1308",
    x"3F3B0EBE",
    x"3F3B0A74",
    x"3F3B0629",
    x"3F3B01DF",
    x"3F3AFD94",
    x"3F3AF94A",
    x"3F3AF4FF",
    x"3F3AF0B4",
    x"3F3AEC69",
    x"3F3AE81E",
    x"3F3AE3D3",
    x"3F3ADF88",
    x"3F3ADB3C",
    x"3F3AD6F1",
    x"3F3AD2A5",
    x"3F3ACE59",
    x"3F3ACA0D",
    x"3F3AC5C1",
    x"3F3AC175",
    x"3F3ABD29",
    x"3F3AB8DD",
    x"3F3AB490",
    x"3F3AB044",
    x"3F3AABF7",
    x"3F3AA7AA",
    x"3F3AA35D",
    x"3F3A9F10",
    x"3F3A9AC3",
    x"3F3A9676",
    x"3F3A9229",
    x"3F3A8DDB",
    x"3F3A898E",
    x"3F3A8540",
    x"3F3A80F2",
    x"3F3A7CA4",
    x"3F3A7856",
    x"3F3A7408",
    x"3F3A6FBA",
    x"3F3A6B6C",
    x"3F3A671D",
    x"3F3A62CF",
    x"3F3A5E80",
    x"3F3A5A31",
    x"3F3A55E2",
    x"3F3A5193",
    x"3F3A4D44",
    x"3F3A48F5",
    x"3F3A44A6",
    x"3F3A4056",
    x"3F3A3C06",
    x"3F3A37B7",
    x"3F3A3367",
    x"3F3A2F17",
    x"3F3A2AC7",
    x"3F3A2677",
    x"3F3A2227",
    x"3F3A1DD6",
    x"3F3A1986",
    x"3F3A1535",
    x"3F3A10E4",
    x"3F3A0C94",
    x"3F3A0843",
    x"3F3A03F2",
    x"3F39FFA1",
    x"3F39FB4F",
    x"3F39F6FE",
    x"3F39F2AC",
    x"3F39EE5B",
    x"3F39EA09",
    x"3F39E5B7",
    x"3F39E165",
    x"3F39DD13",
    x"3F39D8C1",
    x"3F39D46F",
    x"3F39D01D",
    x"3F39CBCA",
    x"3F39C777",
    x"3F39C325",
    x"3F39BED2",
    x"3F39BA7F",
    x"3F39B62C",
    x"3F39B1D9",
    x"3F39AD85",
    x"3F39A932",
    x"3F39A4DF",
    x"3F39A08B",
    x"3F399C37",
    x"3F3997E3",
    x"3F39938F",
    x"3F398F3B",
    x"3F398AE7",
    x"3F398693",
    x"3F39823E",
    x"3F397DEA",
    x"3F397995",
    x"3F397541",
    x"3F3970EC",
    x"3F396C97",
    x"3F396842",
    x"3F3963ED",
    x"3F395F97",
    x"3F395B42",
    x"3F3956EC",
    x"3F395297",
    x"3F394E41",
    x"3F3949EB",
    x"3F394595",
    x"3F39413F",
    x"3F393CE9",
    x"3F393893",
    x"3F39343C",
    x"3F392FE6",
    x"3F392B8F",
    x"3F392738",
    x"3F3922E1",
    x"3F391E8B",
    x"3F391A33",
    x"3F3915DC",
    x"3F391185",
    x"3F390D2E",
    x"3F3908D6",
    x"3F39047E",
    x"3F390027",
    x"3F38FBCF",
    x"3F38F777",
    x"3F38F31F",
    x"3F38EEC7",
    x"3F38EA6E",
    x"3F38E616",
    x"3F38E1BD",
    x"3F38DD65",
    x"3F38D90C",
    x"3F38D4B3",
    x"3F38D05A",
    x"3F38CC01",
    x"3F38C7A8",
    x"3F38C34F",
    x"3F38BEF5",
    x"3F38BA9C",
    x"3F38B642",
    x"3F38B1E8",
    x"3F38AD8E",
    x"3F38A934",
    x"3F38A4DA",
    x"3F38A080",
    x"3F389C26",
    x"3F3897CB",
    x"3F389371",
    x"3F388F16",
    x"3F388ABB",
    x"3F388661",
    x"3F388206",
    x"3F387DAB",
    x"3F38794F",
    x"3F3874F4",
    x"3F387099",
    x"3F386C3D",
    x"3F3867E1",
    x"3F386386",
    x"3F385F2A",
    x"3F385ACE",
    x"3F385672",
    x"3F385216",
    x"3F384DB9",
    x"3F38495D",
    x"3F384500",
    x"3F3840A4",
    x"3F383C47",
    x"3F3837EA",
    x"3F38338D",
    x"3F382F30",
    x"3F382AD3",
    x"3F382676",
    x"3F382218",
    x"3F381DBB",
    x"3F38195D",
    x"3F3814FF",
    x"3F3810A1",
    x"3F380C43",
    x"3F3807E5",
    x"3F380387",
    x"3F37FF29",
    x"3F37FACA",
    x"3F37F66C",
    x"3F37F20D",
    x"3F37EDAF",
    x"3F37E950",
    x"3F37E4F1",
    x"3F37E092",
    x"3F37DC32",
    x"3F37D7D3",
    x"3F37D374",
    x"3F37CF14",
    x"3F37CAB5",
    x"3F37C655",
    x"3F37C1F5",
    x"3F37BD95",
    x"3F37B935",
    x"3F37B4D5",
    x"3F37B074",
    x"3F37AC14",
    x"3F37A7B4",
    x"3F37A353",
    x"3F379EF2",
    x"3F379A91",
    x"3F379630",
    x"3F3791CF",
    x"3F378D6E",
    x"3F37890D",
    x"3F3784AB",
    x"3F37804A",
    x"3F377BE8",
    x"3F377787",
    x"3F377325",
    x"3F376EC3",
    x"3F376A61",
    x"3F3765FE",
    x"3F37619C",
    x"3F375D3A",
    x"3F3758D7",
    x"3F375475",
    x"3F375012",
    x"3F374BAF",
    x"3F37474C",
    x"3F3742E9",
    x"3F373E86",
    x"3F373A23",
    x"3F3735BF",
    x"3F37315C",
    x"3F372CF8",
    x"3F372894",
    x"3F372431",
    x"3F371FCD",
    x"3F371B69",
    x"3F371704",
    x"3F3712A0",
    x"3F370E3C",
    x"3F3709D7",
    x"3F370573",
    x"3F37010E",
    x"3F36FCA9",
    x"3F36F844",
    x"3F36F3DF",
    x"3F36EF7A",
    x"3F36EB15",
    x"3F36E6AF",
    x"3F36E24A",
    x"3F36DDE4",
    x"3F36D97F",
    x"3F36D519",
    x"3F36D0B3",
    x"3F36CC4D",
    x"3F36C7E7",
    x"3F36C380",
    x"3F36BF1A",
    x"3F36BAB4",
    x"3F36B64D",
    x"3F36B1E6",
    x"3F36AD7F",
    x"3F36A919",
    x"3F36A4B2",
    x"3F36A04A",
    x"3F369BE3",
    x"3F36977C",
    x"3F369314",
    x"3F368EAD",
    x"3F368A45",
    x"3F3685DD",
    x"3F368175",
    x"3F367D0D",
    x"3F3678A5",
    x"3F36743D",
    x"3F366FD5",
    x"3F366B6C",
    x"3F366704",
    x"3F36629B",
    x"3F365E32",
    x"3F3659C9",
    x"3F365560",
    x"3F3650F7",
    x"3F364C8E",
    x"3F364825",
    x"3F3643BB",
    x"3F363F52",
    x"3F363AE8",
    x"3F36367E",
    x"3F363214",
    x"3F362DAA",
    x"3F362940",
    x"3F3624D6",
    x"3F36206C",
    x"3F361C01",
    x"3F361797",
    x"3F36132C",
    x"3F360EC1",
    x"3F360A56",
    x"3F3605EB",
    x"3F360180",
    x"3F35FD15",
    x"3F35F8AA",
    x"3F35F43E",
    x"3F35EFD3",
    x"3F35EB67",
    x"3F35E6FB",
    x"3F35E290",
    x"3F35DE24",
    x"3F35D9B8",
    x"3F35D54B",
    x"3F35D0DF",
    x"3F35CC73",
    x"3F35C806",
    x"3F35C39A",
    x"3F35BF2D",
    x"3F35BAC0",
    x"3F35B653",
    x"3F35B1E6",
    x"3F35AD79",
    x"3F35A90B",
    x"3F35A49E",
    x"3F35A031",
    x"3F359BC3",
    x"3F359755",
    x"3F3592E7",
    x"3F358E79",
    x"3F358A0B",
    x"3F35859D",
    x"3F35812F",
    x"3F357CC1",
    x"3F357852",
    x"3F3573E4",
    x"3F356F75",
    x"3F356B06",
    x"3F356697",
    x"3F356228",
    x"3F355DB9",
    x"3F35594A",
    x"3F3554DA",
    x"3F35506B",
    x"3F354BFB",
    x"3F35478C",
    x"3F35431C",
    x"3F353EAC",
    x"3F353A3C",
    x"3F3535CC",
    x"3F35315C",
    x"3F352CEB",
    x"3F35287B",
    x"3F35240A",
    x"3F351F9A",
    x"3F351B29",
    x"3F3516B8",
    x"3F351247",
    x"3F350DD6",
    x"3F350965",
    x"3F3504F3",
    x"3F350082",
    x"3F34FC10",
    x"3F34F79F",
    x"3F34F32D",
    x"3F34EEBB",
    x"3F34EA49",
    x"3F34E5D7",
    x"3F34E165",
    x"3F34DCF2",
    x"3F34D880",
    x"3F34D40D",
    x"3F34CF9B",
    x"3F34CB28",
    x"3F34C6B5",
    x"3F34C242",
    x"3F34BDCF",
    x"3F34B95C",
    x"3F34B4E9",
    x"3F34B075",
    x"3F34AC02",
    x"3F34A78E",
    x"3F34A31B",
    x"3F349EA7",
    x"3F349A33",
    x"3F3495BF",
    x"3F34914B",
    x"3F348CD6",
    x"3F348862",
    x"3F3483ED",
    x"3F347F79",
    x"3F347B04",
    x"3F34768F",
    x"3F34721A",
    x"3F346DA5",
    x"3F346930",
    x"3F3464BB",
    x"3F346046",
    x"3F345BD0",
    x"3F34575B",
    x"3F3452E5",
    x"3F344E6F",
    x"3F3449F9",
    x"3F344583",
    x"3F34410D",
    x"3F343C97",
    x"3F343821",
    x"3F3433AA",
    x"3F342F34",
    x"3F342ABD",
    x"3F342646",
    x"3F3421CF",
    x"3F341D58",
    x"3F3418E1",
    x"3F34146A",
    x"3F340FF3",
    x"3F340B7B",
    x"3F340704",
    x"3F34028C",
    x"3F33FE14",
    x"3F33F99D",
    x"3F33F525",
    x"3F33F0AD",
    x"3F33EC34",
    x"3F33E7BC",
    x"3F33E344",
    x"3F33DECB",
    x"3F33DA53",
    x"3F33D5DA",
    x"3F33D161",
    x"3F33CCE8",
    x"3F33C86F",
    x"3F33C3F6",
    x"3F33BF7D",
    x"3F33BB03",
    x"3F33B68A",
    x"3F33B210",
    x"3F33AD97",
    x"3F33A91D",
    x"3F33A4A3",
    x"3F33A029",
    x"3F339BAF",
    x"3F339735",
    x"3F3392BA",
    x"3F338E40",
    x"3F3389C5",
    x"3F33854B",
    x"3F3380D0",
    x"3F337C55",
    x"3F3377DA",
    x"3F33735F",
    x"3F336EE4",
    x"3F336A68",
    x"3F3365ED",
    x"3F336171",
    x"3F335CF6",
    x"3F33587A",
    x"3F3353FE",
    x"3F334F82",
    x"3F334B06",
    x"3F33468A",
    x"3F33420E",
    x"3F333D91",
    x"3F333915",
    x"3F333498",
    x"3F33301B",
    x"3F332B9F",
    x"3F332722",
    x"3F3322A5",
    x"3F331E27",
    x"3F3319AA",
    x"3F33152D",
    x"3F3310AF",
    x"3F330C32",
    x"3F3307B4",
    x"3F330336",
    x"3F32FEB8",
    x"3F32FA3A",
    x"3F32F5BC",
    x"3F32F13E",
    x"3F32ECC0",
    x"3F32E841",
    x"3F32E3C3",
    x"3F32DF44",
    x"3F32DAC5",
    x"3F32D646",
    x"3F32D1C7",
    x"3F32CD48",
    x"3F32C8C9",
    x"3F32C44A",
    x"3F32BFCA",
    x"3F32BB4B",
    x"3F32B6CB",
    x"3F32B24C",
    x"3F32ADCC",
    x"3F32A94C",
    x"3F32A4CC",
    x"3F32A04C",
    x"3F329BCB",
    x"3F32974B",
    x"3F3292CA",
    x"3F328E4A",
    x"3F3289C9",
    x"3F328548",
    x"3F3280C7",
    x"3F327C46",
    x"3F3277C5",
    x"3F327344",
    x"3F326EC3",
    x"3F326A41",
    x"3F3265C0",
    x"3F32613E",
    x"3F325CBC",
    x"3F32583A",
    x"3F3253B8",
    x"3F324F36",
    x"3F324AB4",
    x"3F324632",
    x"3F3241AF",
    x"3F323D2D",
    x"3F3238AA",
    x"3F323427",
    x"3F322FA5",
    x"3F322B22",
    x"3F32269E",
    x"3F32221B",
    x"3F321D98",
    x"3F321915",
    x"3F321491",
    x"3F32100E",
    x"3F320B8A",
    x"3F320706",
    x"3F320282",
    x"3F31FDFE",
    x"3F31F97A",
    x"3F31F4F6",
    x"3F31F071",
    x"3F31EBED",
    x"3F31E768",
    x"3F31E2E4",
    x"3F31DE5F",
    x"3F31D9DA",
    x"3F31D555",
    x"3F31D0D0",
    x"3F31CC4B",
    x"3F31C7C5",
    x"3F31C340",
    x"3F31BEBA",
    x"3F31BA35",
    x"3F31B5AF",
    x"3F31B129",
    x"3F31ACA3",
    x"3F31A81D",
    x"3F31A397",
    x"3F319F11",
    x"3F319A8A",
    x"3F319604",
    x"3F31917D",
    x"3F318CF6",
    x"3F318870",
    x"3F3183E9",
    x"3F317F62",
    x"3F317ADB",
    x"3F317653",
    x"3F3171CC",
    x"3F316D44",
    x"3F3168BD",
    x"3F316435",
    x"3F315FAD",
    x"3F315B26",
    x"3F31569E",
    x"3F315215",
    x"3F314D8D",
    x"3F314905",
    x"3F31447D",
    x"3F313FF4",
    x"3F313B6B",
    x"3F3136E3",
    x"3F31325A",
    x"3F312DD1",
    x"3F312948",
    x"3F3124BF",
    x"3F312035",
    x"3F311BAC",
    x"3F311722",
    x"3F311299",
    x"3F310E0F",
    x"3F310985",
    x"3F3104FB",
    x"3F310071",
    x"3F30FBE7",
    x"3F30F75D",
    x"3F30F2D3",
    x"3F30EE48",
    x"3F30E9BE",
    x"3F30E533",
    x"3F30E0A8",
    x"3F30DC1D",
    x"3F30D792",
    x"3F30D307",
    x"3F30CE7C",
    x"3F30C9F1",
    x"3F30C566",
    x"3F30C0DA",
    x"3F30BC4E",
    x"3F30B7C3",
    x"3F30B337",
    x"3F30AEAB",
    x"3F30AA1F",
    x"3F30A593",
    x"3F30A106",
    x"3F309C7A",
    x"3F3097EE",
    x"3F309361",
    x"3F308ED4",
    x"3F308A48",
    x"3F3085BB",
    x"3F30812E",
    x"3F307CA1",
    x"3F307813",
    x"3F307386",
    x"3F306EF9",
    x"3F306A6B",
    x"3F3065DD",
    x"3F306150",
    x"3F305CC2",
    x"3F305834",
    x"3F3053A6",
    x"3F304F18",
    x"3F304A89",
    x"3F3045FB",
    x"3F30416C",
    x"3F303CDE",
    x"3F30384F",
    x"3F3033C0",
    x"3F302F31",
    x"3F302AA2",
    x"3F302613",
    x"3F302184",
    x"3F301CF5",
    x"3F301865",
    x"3F3013D6",
    x"3F300F46",
    x"3F300AB6",
    x"3F300626",
    x"3F300196",
    x"3F2FFD06",
    x"3F2FF876",
    x"3F2FF3E6",
    x"3F2FEF56",
    x"3F2FEAC5",
    x"3F2FE634",
    x"3F2FE1A4",
    x"3F2FDD13",
    x"3F2FD882",
    x"3F2FD3F1",
    x"3F2FCF60",
    x"3F2FCACF",
    x"3F2FC63D",
    x"3F2FC1AC",
    x"3F2FBD1A",
    x"3F2FB888",
    x"3F2FB3F7",
    x"3F2FAF65",
    x"3F2FAAD3",
    x"3F2FA641",
    x"3F2FA1AF",
    x"3F2F9D1C",
    x"3F2F988A",
    x"3F2F93F7",
    x"3F2F8F65",
    x"3F2F8AD2",
    x"3F2F863F",
    x"3F2F81AC",
    x"3F2F7D19",
    x"3F2F7886",
    x"3F2F73F3",
    x"3F2F6F5F",
    x"3F2F6ACC",
    x"3F2F6638",
    x"3F2F61A5",
    x"3F2F5D11",
    x"3F2F587D",
    x"3F2F53E9",
    x"3F2F4F55",
    x"3F2F4AC1",
    x"3F2F462C",
    x"3F2F4198",
    x"3F2F3D03",
    x"3F2F386F",
    x"3F2F33DA",
    x"3F2F2F45",
    x"3F2F2AB0",
    x"3F2F261B",
    x"3F2F2186",
    x"3F2F1CF1",
    x"3F2F185B",
    x"3F2F13C6",
    x"3F2F0F30",
    x"3F2F0A9B",
    x"3F2F0605",
    x"3F2F016F",
    x"3F2EFCD9",
    x"3F2EF843",
    x"3F2EF3AD",
    x"3F2EEF16",
    x"3F2EEA80",
    x"3F2EE5E9",
    x"3F2EE153",
    x"3F2EDCBC",
    x"3F2ED825",
    x"3F2ED38E",
    x"3F2ECEF7",
    x"3F2ECA60",
    x"3F2EC5C9",
    x"3F2EC131",
    x"3F2EBC9A",
    x"3F2EB802",
    x"3F2EB36B",
    x"3F2EAED3",
    x"3F2EAA3B",
    x"3F2EA5A3",
    x"3F2EA10B",
    x"3F2E9C73",
    x"3F2E97DA",
    x"3F2E9342",
    x"3F2E8EA9",
    x"3F2E8A11",
    x"3F2E8578",
    x"3F2E80DF",
    x"3F2E7C46",
    x"3F2E77AD",
    x"3F2E7314",
    x"3F2E6E7B",
    x"3F2E69E1",
    x"3F2E6548",
    x"3F2E60AE",
    x"3F2E5C15",
    x"3F2E577B",
    x"3F2E52E1",
    x"3F2E4E47",
    x"3F2E49AD",
    x"3F2E4513",
    x"3F2E4078",
    x"3F2E3BDE",
    x"3F2E3743",
    x"3F2E32A9",
    x"3F2E2E0E",
    x"3F2E2973",
    x"3F2E24D8",
    x"3F2E203D",
    x"3F2E1BA2",
    x"3F2E1707",
    x"3F2E126B",
    x"3F2E0DD0",
    x"3F2E0934",
    x"3F2E0499",
    x"3F2DFFFD",
    x"3F2DFB61",
    x"3F2DF6C5",
    x"3F2DF229",
    x"3F2DED8D",
    x"3F2DE8F0",
    x"3F2DE454",
    x"3F2DDFB8",
    x"3F2DDB1B",
    x"3F2DD67E",
    x"3F2DD1E1",
    x"3F2DCD44",
    x"3F2DC8A7",
    x"3F2DC40A",
    x"3F2DBF6D",
    x"3F2DBAD0",
    x"3F2DB632",
    x"3F2DB195",
    x"3F2DACF7",
    x"3F2DA859",
    x"3F2DA3BB",
    x"3F2D9F1D",
    x"3F2D9A7F",
    x"3F2D95E1",
    x"3F2D9143",
    x"3F2D8CA4",
    x"3F2D8806",
    x"3F2D8367",
    x"3F2D7EC9",
    x"3F2D7A2A",
    x"3F2D758B",
    x"3F2D70EC",
    x"3F2D6C4D",
    x"3F2D67AD",
    x"3F2D630E",
    x"3F2D5E6F",
    x"3F2D59CF",
    x"3F2D552F",
    x"3F2D5090",
    x"3F2D4BF0",
    x"3F2D4750",
    x"3F2D42B0",
    x"3F2D3E10",
    x"3F2D396F",
    x"3F2D34CF",
    x"3F2D302E",
    x"3F2D2B8E",
    x"3F2D26ED",
    x"3F2D224C",
    x"3F2D1DAB",
    x"3F2D190A",
    x"3F2D1469",
    x"3F2D0FC8",
    x"3F2D0B27",
    x"3F2D0685",
    x"3F2D01E4",
    x"3F2CFD42",
    x"3F2CF8A0",
    x"3F2CF3FF",
    x"3F2CEF5D",
    x"3F2CEABB",
    x"3F2CE618",
    x"3F2CE176",
    x"3F2CDCD4",
    x"3F2CD831",
    x"3F2CD38F",
    x"3F2CCEEC",
    x"3F2CCA49",
    x"3F2CC5A6",
    x"3F2CC103",
    x"3F2CBC60",
    x"3F2CB7BD",
    x"3F2CB31A",
    x"3F2CAE76",
    x"3F2CA9D3",
    x"3F2CA52F",
    x"3F2CA08C",
    x"3F2C9BE8",
    x"3F2C9744",
    x"3F2C92A0",
    x"3F2C8DFC",
    x"3F2C8957",
    x"3F2C84B3",
    x"3F2C800F",
    x"3F2C7B6A",
    x"3F2C76C5",
    x"3F2C7221",
    x"3F2C6D7C",
    x"3F2C68D7",
    x"3F2C6432",
    x"3F2C5F8D",
    x"3F2C5AE7",
    x"3F2C5642",
    x"3F2C519D",
    x"3F2C4CF7",
    x"3F2C4851",
    x"3F2C43AB",
    x"3F2C3F06",
    x"3F2C3A60",
    x"3F2C35B9",
    x"3F2C3113",
    x"3F2C2C6D",
    x"3F2C27C7",
    x"3F2C2320",
    x"3F2C1E79",
    x"3F2C19D3",
    x"3F2C152C",
    x"3F2C1085",
    x"3F2C0BDE",
    x"3F2C0737",
    x"3F2C028F",
    x"3F2BFDE8",
    x"3F2BF941",
    x"3F2BF499",
    x"3F2BEFF1",
    x"3F2BEB4A",
    x"3F2BE6A2",
    x"3F2BE1FA",
    x"3F2BDD52",
    x"3F2BD8AA",
    x"3F2BD401",
    x"3F2BCF59",
    x"3F2BCAB0",
    x"3F2BC608",
    x"3F2BC15F",
    x"3F2BBCB6",
    x"3F2BB80D",
    x"3F2BB364",
    x"3F2BAEBB",
    x"3F2BAA12",
    x"3F2BA569",
    x"3F2BA0BF",
    x"3F2B9C16",
    x"3F2B976C",
    x"3F2B92C2",
    x"3F2B8E19",
    x"3F2B896F",
    x"3F2B84C5",
    x"3F2B801A",
    x"3F2B7B70",
    x"3F2B76C6",
    x"3F2B721B",
    x"3F2B6D71",
    x"3F2B68C6",
    x"3F2B641B",
    x"3F2B5F71",
    x"3F2B5AC6",
    x"3F2B561B",
    x"3F2B516F",
    x"3F2B4CC4",
    x"3F2B4819",
    x"3F2B436D",
    x"3F2B3EC2",
    x"3F2B3A16",
    x"3F2B356A",
    x"3F2B30BE",
    x"3F2B2C12",
    x"3F2B2766",
    x"3F2B22BA",
    x"3F2B1E0E",
    x"3F2B1961",
    x"3F2B14B5",
    x"3F2B1008",
    x"3F2B0B5B",
    x"3F2B06AF",
    x"3F2B0202",
    x"3F2AFD55",
    x"3F2AF8A7",
    x"3F2AF3FA",
    x"3F2AEF4D",
    x"3F2AEA9F",
    x"3F2AE5F2",
    x"3F2AE144",
    x"3F2ADC96",
    x"3F2AD7E9",
    x"3F2AD33B",
    x"3F2ACE8D",
    x"3F2AC9DE",
    x"3F2AC530",
    x"3F2AC082",
    x"3F2ABBD3",
    x"3F2AB725",
    x"3F2AB276",
    x"3F2AADC7",
    x"3F2AA918",
    x"3F2AA469",
    x"3F2A9FBA",
    x"3F2A9B0B",
    x"3F2A965C",
    x"3F2A91AC",
    x"3F2A8CFD",
    x"3F2A884D",
    x"3F2A839E",
    x"3F2A7EEE",
    x"3F2A7A3E",
    x"3F2A758E",
    x"3F2A70DE",
    x"3F2A6C2E",
    x"3F2A677D",
    x"3F2A62CD",
    x"3F2A5E1C",
    x"3F2A596C",
    x"3F2A54BB",
    x"3F2A500A",
    x"3F2A4B59",
    x"3F2A46A8",
    x"3F2A41F7",
    x"3F2A3D46",
    x"3F2A3894",
    x"3F2A33E3",
    x"3F2A2F31",
    x"3F2A2A80",
    x"3F2A25CE",
    x"3F2A211C",
    x"3F2A1C6A",
    x"3F2A17B8",
    x"3F2A1306",
    x"3F2A0E54",
    x"3F2A09A1",
    x"3F2A04EF",
    x"3F2A003C",
    x"3F29FB89",
    x"3F29F6D7",
    x"3F29F224",
    x"3F29ED71",
    x"3F29E8BE",
    x"3F29E40B",
    x"3F29DF57",
    x"3F29DAA4",
    x"3F29D5F0",
    x"3F29D13D",
    x"3F29CC89",
    x"3F29C7D5",
    x"3F29C321",
    x"3F29BE6D",
    x"3F29B9B9",
    x"3F29B505",
    x"3F29B051",
    x"3F29AB9C",
    x"3F29A6E8",
    x"3F29A233",
    x"3F299D7E",
    x"3F2998CA",
    x"3F299415",
    x"3F298F60",
    x"3F298AAA",
    x"3F2985F5",
    x"3F298140",
    x"3F297C8A",
    x"3F2977D5",
    x"3F29731F",
    x"3F296E69",
    x"3F2969B4",
    x"3F2964FE",
    x"3F296048",
    x"3F295B91",
    x"3F2956DB",
    x"3F295225",
    x"3F294D6E",
    x"3F2948B8",
    x"3F294401",
    x"3F293F4A",
    x"3F293A93",
    x"3F2935DD",
    x"3F293125",
    x"3F292C6E",
    x"3F2927B7",
    x"3F292300",
    x"3F291E48",
    x"3F291991",
    x"3F2914D9",
    x"3F291021",
    x"3F290B69",
    x"3F2906B1",
    x"3F2901F9",
    x"3F28FD41",
    x"3F28F889",
    x"3F28F3D0",
    x"3F28EF18",
    x"3F28EA5F",
    x"3F28E5A6",
    x"3F28E0EE",
    x"3F28DC35",
    x"3F28D77C",
    x"3F28D2C3",
    x"3F28CE09",
    x"3F28C950",
    x"3F28C497",
    x"3F28BFDD",
    x"3F28BB23",
    x"3F28B66A",
    x"3F28B1B0",
    x"3F28ACF6",
    x"3F28A83C",
    x"3F28A382",
    x"3F289EC8",
    x"3F289A0D",
    x"3F289553",
    x"3F289098",
    x"3F288BDE",
    x"3F288723",
    x"3F288268",
    x"3F287DAD",
    x"3F2878F2",
    x"3F287437",
    x"3F286F7C",
    x"3F286AC0",
    x"3F286605",
    x"3F286149",
    x"3F285C8E",
    x"3F2857D2",
    x"3F285316",
    x"3F284E5A",
    x"3F28499E",
    x"3F2844E2",
    x"3F284026",
    x"3F283B69",
    x"3F2836AD",
    x"3F2831F0",
    x"3F282D34",
    x"3F282877",
    x"3F2823BA",
    x"3F281EFD",
    x"3F281A40",
    x"3F281583",
    x"3F2810C6",
    x"3F280C08",
    x"3F28074B",
    x"3F28028D",
    x"3F27FDD0",
    x"3F27F912",
    x"3F27F454",
    x"3F27EF96",
    x"3F27EAD8",
    x"3F27E61A",
    x"3F27E15B",
    x"3F27DC9D",
    x"3F27D7DE",
    x"3F27D320",
    x"3F27CE61",
    x"3F27C9A2",
    x"3F27C4E4",
    x"3F27C025",
    x"3F27BB65",
    x"3F27B6A6",
    x"3F27B1E7",
    x"3F27AD28",
    x"3F27A868",
    x"3F27A3A8",
    x"3F279EE9",
    x"3F279A29",
    x"3F279569",
    x"3F2790A9",
    x"3F278BE9",
    x"3F278729",
    x"3F278268",
    x"3F277DA8",
    x"3F2778E8",
    x"3F277427",
    x"3F276F66",
    x"3F276AA5",
    x"3F2765E5",
    x"3F276123",
    x"3F275C62",
    x"3F2757A1",
    x"3F2752E0",
    x"3F274E1E",
    x"3F27495D",
    x"3F27449B",
    x"3F273FDA",
    x"3F273B18",
    x"3F273656",
    x"3F273194",
    x"3F272CD2",
    x"3F272810",
    x"3F27234D",
    x"3F271E8B",
    x"3F2719C8",
    x"3F271506",
    x"3F271043",
    x"3F270B80",
    x"3F2706BD",
    x"3F2701FA",
    x"3F26FD37",
    x"3F26F874",
    x"3F26F3B0",
    x"3F26EEED",
    x"3F26EA2A",
    x"3F26E566",
    x"3F26E0A2",
    x"3F26DBDE",
    x"3F26D71A",
    x"3F26D256",
    x"3F26CD92",
    x"3F26C8CE",
    x"3F26C40A",
    x"3F26BF45",
    x"3F26BA81",
    x"3F26B5BC",
    x"3F26B0F7",
    x"3F26AC33",
    x"3F26A76E",
    x"3F26A2A9",
    x"3F269DE3",
    x"3F26991E",
    x"3F269459",
    x"3F268F93",
    x"3F268ACE",
    x"3F268608",
    x"3F268143",
    x"3F267C7D",
    x"3F2677B7",
    x"3F2672F1",
    x"3F266E2B",
    x"3F266964",
    x"3F26649E",
    x"3F265FD8",
    x"3F265B11",
    x"3F26564A",
    x"3F265184",
    x"3F264CBD",
    x"3F2647F6",
    x"3F26432F",
    x"3F263E68",
    x"3F2639A0",
    x"3F2634D9",
    x"3F263012",
    x"3F262B4A",
    x"3F262682",
    x"3F2621BB",
    x"3F261CF3",
    x"3F26182B",
    x"3F261363",
    x"3F260E9B",
    x"3F2609D3",
    x"3F26050A",
    x"3F260042",
    x"3F25FB79",
    x"3F25F6B1",
    x"3F25F1E8",
    x"3F25ED1F",
    x"3F25E856",
    x"3F25E38D",
    x"3F25DEC4",
    x"3F25D9FB",
    x"3F25D531",
    x"3F25D068",
    x"3F25CB9E",
    x"3F25C6D5",
    x"3F25C20B",
    x"3F25BD41",
    x"3F25B877",
    x"3F25B3AD",
    x"3F25AEE3",
    x"3F25AA19",
    x"3F25A54E",
    x"3F25A084",
    x"3F259BB9",
    x"3F2596EF",
    x"3F259224",
    x"3F258D59",
    x"3F25888E",
    x"3F2583C3",
    x"3F257EF8",
    x"3F257A2D",
    x"3F257562",
    x"3F257096",
    x"3F256BCB",
    x"3F2566FF",
    x"3F256233",
    x"3F255D67",
    x"3F25589B",
    x"3F2553CF",
    x"3F254F03",
    x"3F254A37",
    x"3F25456B",
    x"3F25409E",
    x"3F253BD2",
    x"3F253705",
    x"3F253238",
    x"3F252D6C",
    x"3F25289F",
    x"3F2523D2",
    x"3F251F04",
    x"3F251A37",
    x"3F25156A",
    x"3F25109C",
    x"3F250BCF",
    x"3F250701",
    x"3F250234",
    x"3F24FD66",
    x"3F24F898",
    x"3F24F3CA",
    x"3F24EEFC",
    x"3F24EA2D",
    x"3F24E55F",
    x"3F24E091",
    x"3F24DBC2",
    x"3F24D6F4",
    x"3F24D225",
    x"3F24CD56",
    x"3F24C887",
    x"3F24C3B8",
    x"3F24BEE9",
    x"3F24BA1A",
    x"3F24B54A",
    x"3F24B07B",
    x"3F24ABAC",
    x"3F24A6DC",
    x"3F24A20C",
    x"3F249D3C",
    x"3F24986D",
    x"3F24939C",
    x"3F248ECC",
    x"3F2489FC",
    x"3F24852C",
    x"3F24805B",
    x"3F247B8B",
    x"3F2476BA",
    x"3F2471EA",
    x"3F246D19",
    x"3F246848",
    x"3F246377",
    x"3F245EA6",
    x"3F2459D5",
    x"3F245503",
    x"3F245032",
    x"3F244B60",
    x"3F24468F",
    x"3F2441BD",
    x"3F243CEB",
    x"3F24381A",
    x"3F243348",
    x"3F242E75",
    x"3F2429A3",
    x"3F2424D1",
    x"3F241FFF",
    x"3F241B2C",
    x"3F24165A",
    x"3F241187",
    x"3F240CB4",
    x"3F2407E1",
    x"3F24030E",
    x"3F23FE3B",
    x"3F23F968",
    x"3F23F495",
    x"3F23EFC1",
    x"3F23EAEE",
    x"3F23E61A",
    x"3F23E147",
    x"3F23DC73",
    x"3F23D79F",
    x"3F23D2CB",
    x"3F23CDF7",
    x"3F23C923",
    x"3F23C44F",
    x"3F23BF7A",
    x"3F23BAA6",
    x"3F23B5D1",
    x"3F23B0FC",
    x"3F23AC28",
    x"3F23A753",
    x"3F23A27E",
    x"3F239DA9",
    x"3F2398D4",
    x"3F2393FE",
    x"3F238F29",
    x"3F238A54",
    x"3F23857E",
    x"3F2380A8",
    x"3F237BD3",
    x"3F2376FD",
    x"3F237227",
    x"3F236D51",
    x"3F23687B",
    x"3F2363A5",
    x"3F235ECE",
    x"3F2359F8",
    x"3F235521",
    x"3F23504B",
    x"3F234B74",
    x"3F23469D",
    x"3F2341C6",
    x"3F233CEF",
    x"3F233818",
    x"3F233341",
    x"3F232E6A",
    x"3F232992",
    x"3F2324BB",
    x"3F231FE3",
    x"3F231B0B",
    x"3F231633",
    x"3F23115C",
    x"3F230C84",
    x"3F2307AB",
    x"3F2302D3",
    x"3F22FDFB",
    x"3F22F923",
    x"3F22F44A",
    x"3F22EF72",
    x"3F22EA99",
    x"3F22E5C0",
    x"3F22E0E7",
    x"3F22DC0E",
    x"3F22D735",
    x"3F22D25C",
    x"3F22CD83",
    x"3F22C8A9",
    x"3F22C3D0",
    x"3F22BEF6",
    x"3F22BA1D",
    x"3F22B543",
    x"3F22B069",
    x"3F22AB8F",
    x"3F22A6B5",
    x"3F22A1DB",
    x"3F229D00",
    x"3F229826",
    x"3F22934C",
    x"3F228E71",
    x"3F228996",
    x"3F2284BC",
    x"3F227FE1",
    x"3F227B06",
    x"3F22762B",
    x"3F227150",
    x"3F226C74",
    x"3F226799",
    x"3F2262BE",
    x"3F225DE2",
    x"3F225907",
    x"3F22542B",
    x"3F224F4F",
    x"3F224A73",
    x"3F224597",
    x"3F2240BB",
    x"3F223BDF",
    x"3F223702",
    x"3F223226",
    x"3F222D4A",
    x"3F22286D",
    x"3F222390",
    x"3F221EB3",
    x"3F2219D7",
    x"3F2214FA",
    x"3F22101C",
    x"3F220B3F",
    x"3F220662",
    x"3F220185",
    x"3F21FCA7",
    x"3F21F7C9",
    x"3F21F2EC",
    x"3F21EE0E",
    x"3F21E930",
    x"3F21E452",
    x"3F21DF74",
    x"3F21DA96",
    x"3F21D5B8",
    x"3F21D0D9",
    x"3F21CBFB",
    x"3F21C71C",
    x"3F21C23E",
    x"3F21BD5F",
    x"3F21B880",
    x"3F21B3A1",
    x"3F21AEC2",
    x"3F21A9E3",
    x"3F21A504",
    x"3F21A024",
    x"3F219B45",
    x"3F219665",
    x"3F219186",
    x"3F218CA6",
    x"3F2187C6",
    x"3F2182E6",
    x"3F217E06",
    x"3F217926",
    x"3F217446",
    x"3F216F66",
    x"3F216A85",
    x"3F2165A5",
    x"3F2160C4",
    x"3F215BE3",
    x"3F215703",
    x"3F215222",
    x"3F214D41",
    x"3F214860",
    x"3F21437E",
    x"3F213E9D",
    x"3F2139BC",
    x"3F2134DA",
    x"3F212FF9",
    x"3F212B17",
    x"3F212635",
    x"3F212153",
    x"3F211C71",
    x"3F21178F",
    x"3F2112AD",
    x"3F210DCB",
    x"3F2108E9",
    x"3F210406",
    x"3F20FF24",
    x"3F20FA41",
    x"3F20F55E",
    x"3F20F07B",
    x"3F20EB99",
    x"3F20E6B5",
    x"3F20E1D2",
    x"3F20DCEF",
    x"3F20D80C",
    x"3F20D328",
    x"3F20CE45",
    x"3F20C961",
    x"3F20C47E",
    x"3F20BF9A",
    x"3F20BAB6",
    x"3F20B5D2",
    x"3F20B0EE",
    x"3F20AC0A",
    x"3F20A725",
    x"3F20A241",
    x"3F209D5C",
    x"3F209878",
    x"3F209393",
    x"3F208EAE",
    x"3F2089CA",
    x"3F2084E5",
    x"3F208000",
    x"3F207B1A",
    x"3F207635",
    x"3F207150",
    x"3F206C6A",
    x"3F206785",
    x"3F20629F",
    x"3F205DB9",
    x"3F2058D4",
    x"3F2053EE",
    x"3F204F08",
    x"3F204A21",
    x"3F20453B",
    x"3F204055",
    x"3F203B6F",
    x"3F203688",
    x"3F2031A1",
    x"3F202CBB",
    x"3F2027D4",
    x"3F2022ED",
    x"3F201E06",
    x"3F20191F",
    x"3F201438",
    x"3F200F50",
    x"3F200A69",
    x"3F200582",
    x"3F20009A",
    x"3F1FFBB2",
    x"3F1FF6CB",
    x"3F1FF1E3",
    x"3F1FECFB",
    x"3F1FE813",
    x"3F1FE32B",
    x"3F1FDE42",
    x"3F1FD95A",
    x"3F1FD472",
    x"3F1FCF89",
    x"3F1FCAA0",
    x"3F1FC5B8",
    x"3F1FC0CF",
    x"3F1FBBE6",
    x"3F1FB6FD",
    x"3F1FB214",
    x"3F1FAD2B",
    x"3F1FA841",
    x"3F1FA358",
    x"3F1F9E6E",
    x"3F1F9985",
    x"3F1F949B",
    x"3F1F8FB1",
    x"3F1F8AC7",
    x"3F1F85DD",
    x"3F1F80F3",
    x"3F1F7C09",
    x"3F1F771F",
    x"3F1F7235",
    x"3F1F6D4A",
    x"3F1F6860",
    x"3F1F6375",
    x"3F1F5E8A",
    x"3F1F599F",
    x"3F1F54B4",
    x"3F1F4FC9",
    x"3F1F4ADE",
    x"3F1F45F3",
    x"3F1F4108",
    x"3F1F3C1C",
    x"3F1F3731",
    x"3F1F3245",
    x"3F1F2D59",
    x"3F1F286E",
    x"3F1F2382",
    x"3F1F1E96",
    x"3F1F19AA",
    x"3F1F14BD",
    x"3F1F0FD1",
    x"3F1F0AE5",
    x"3F1F05F8",
    x"3F1F010C",
    x"3F1EFC1F",
    x"3F1EF732",
    x"3F1EF245",
    x"3F1EED59",
    x"3F1EE86C",
    x"3F1EE37E",
    x"3F1EDE91",
    x"3F1ED9A4",
    x"3F1ED4B6",
    x"3F1ECFC9",
    x"3F1ECADB",
    x"3F1EC5ED",
    x"3F1EC100",
    x"3F1EBC12",
    x"3F1EB724",
    x"3F1EB236",
    x"3F1EAD47",
    x"3F1EA859",
    x"3F1EA36B",
    x"3F1E9E7C",
    x"3F1E998E",
    x"3F1E949F",
    x"3F1E8FB0",
    x"3F1E8AC1",
    x"3F1E85D2",
    x"3F1E80E3",
    x"3F1E7BF4",
    x"3F1E7705",
    x"3F1E7216",
    x"3F1E6D26",
    x"3F1E6837",
    x"3F1E6347",
    x"3F1E5E57",
    x"3F1E5968",
    x"3F1E5478",
    x"3F1E4F88",
    x"3F1E4A98",
    x"3F1E45A7",
    x"3F1E40B7",
    x"3F1E3BC7",
    x"3F1E36D6",
    x"3F1E31E6",
    x"3F1E2CF5",
    x"3F1E2804",
    x"3F1E2313",
    x"3F1E1E22",
    x"3F1E1931",
    x"3F1E1440",
    x"3F1E0F4F",
    x"3F1E0A5D",
    x"3F1E056C",
    x"3F1E007B",
    x"3F1DFB89",
    x"3F1DF697",
    x"3F1DF1A5",
    x"3F1DECB3",
    x"3F1DE7C1",
    x"3F1DE2CF",
    x"3F1DDDDD",
    x"3F1DD8EB",
    x"3F1DD3F8",
    x"3F1DCF06",
    x"3F1DCA13",
    x"3F1DC521",
    x"3F1DC02E",
    x"3F1DBB3B",
    x"3F1DB648",
    x"3F1DB155",
    x"3F1DAC62",
    x"3F1DA76F",
    x"3F1DA27B",
    x"3F1D9D88",
    x"3F1D9894",
    x"3F1D93A1",
    x"3F1D8EAD",
    x"3F1D89B9",
    x"3F1D84C5",
    x"3F1D7FD1",
    x"3F1D7ADD",
    x"3F1D75E9",
    x"3F1D70F5",
    x"3F1D6C00",
    x"3F1D670C",
    x"3F1D6217",
    x"3F1D5D23",
    x"3F1D582E",
    x"3F1D5339",
    x"3F1D4E44",
    x"3F1D494F",
    x"3F1D445A",
    x"3F1D3F65",
    x"3F1D3A6F",
    x"3F1D357A",
    x"3F1D3084",
    x"3F1D2B8F",
    x"3F1D2699",
    x"3F1D21A3",
    x"3F1D1CAD",
    x"3F1D17B7",
    x"3F1D12C1",
    x"3F1D0DCB",
    x"3F1D08D5",
    x"3F1D03DE",
    x"3F1CFEE8",
    x"3F1CF9F1",
    x"3F1CF4FB",
    x"3F1CF004",
    x"3F1CEB0D",
    x"3F1CE616",
    x"3F1CE11F",
    x"3F1CDC28",
    x"3F1CD731",
    x"3F1CD239",
    x"3F1CCD42",
    x"3F1CC84B",
    x"3F1CC353",
    x"3F1CBE5B",
    x"3F1CB963",
    x"3F1CB46C",
    x"3F1CAF74",
    x"3F1CAA7C",
    x"3F1CA583",
    x"3F1CA08B",
    x"3F1C9B93",
    x"3F1C969A",
    x"3F1C91A2",
    x"3F1C8CA9",
    x"3F1C87B0",
    x"3F1C82B8",
    x"3F1C7DBF",
    x"3F1C78C6",
    x"3F1C73CC",
    x"3F1C6ED3",
    x"3F1C69DA",
    x"3F1C64E1",
    x"3F1C5FE7",
    x"3F1C5AEE",
    x"3F1C55F4",
    x"3F1C50FA",
    x"3F1C4C00",
    x"3F1C4706",
    x"3F1C420C",
    x"3F1C3D12",
    x"3F1C3818",
    x"3F1C331D",
    x"3F1C2E23",
    x"3F1C2929",
    x"3F1C242E",
    x"3F1C1F33",
    x"3F1C1A38",
    x"3F1C153D",
    x"3F1C1042",
    x"3F1C0B47",
    x"3F1C064C",
    x"3F1C0151",
    x"3F1BFC56",
    x"3F1BF75A",
    x"3F1BF25F",
    x"3F1BED63",
    x"3F1BE867",
    x"3F1BE36B",
    x"3F1BDE6F",
    x"3F1BD973",
    x"3F1BD477",
    x"3F1BCF7B",
    x"3F1BCA7F",
    x"3F1BC582",
    x"3F1BC086",
    x"3F1BBB89",
    x"3F1BB68D",
    x"3F1BB190",
    x"3F1BAC93",
    x"3F1BA796",
    x"3F1BA299",
    x"3F1B9D9C",
    x"3F1B989E",
    x"3F1B93A1",
    x"3F1B8EA4",
    x"3F1B89A6",
    x"3F1B84A9",
    x"3F1B7FAB",
    x"3F1B7AAD",
    x"3F1B75AF",
    x"3F1B70B1",
    x"3F1B6BB3",
    x"3F1B66B5",
    x"3F1B61B7",
    x"3F1B5CB8",
    x"3F1B57BA",
    x"3F1B52BB",
    x"3F1B4DBD",
    x"3F1B48BE",
    x"3F1B43BF",
    x"3F1B3EC0",
    x"3F1B39C1",
    x"3F1B34C2",
    x"3F1B2FC3",
    x"3F1B2AC3",
    x"3F1B25C4",
    x"3F1B20C4",
    x"3F1B1BC5",
    x"3F1B16C5",
    x"3F1B11C5",
    x"3F1B0CC6",
    x"3F1B07C6",
    x"3F1B02C6",
    x"3F1AFDC5",
    x"3F1AF8C5",
    x"3F1AF3C5",
    x"3F1AEEC4",
    x"3F1AE9C4",
    x"3F1AE4C3",
    x"3F1ADFC3",
    x"3F1ADAC2",
    x"3F1AD5C1",
    x"3F1AD0C0",
    x"3F1ACBBF",
    x"3F1AC6BE",
    x"3F1AC1BC",
    x"3F1ABCBB",
    x"3F1AB7BA",
    x"3F1AB2B8",
    x"3F1AADB6",
    x"3F1AA8B5",
    x"3F1AA3B3",
    x"3F1A9EB1",
    x"3F1A99AF",
    x"3F1A94AD",
    x"3F1A8FAB",
    x"3F1A8AA8",
    x"3F1A85A6",
    x"3F1A80A3",
    x"3F1A7BA1",
    x"3F1A769E",
    x"3F1A719B",
    x"3F1A6C99",
    x"3F1A6796",
    x"3F1A6293",
    x"3F1A5D8F",
    x"3F1A588C",
    x"3F1A5389",
    x"3F1A4E86",
    x"3F1A4982",
    x"3F1A447E",
    x"3F1A3F7B",
    x"3F1A3A77",
    x"3F1A3573",
    x"3F1A306F",
    x"3F1A2B6B",
    x"3F1A2667",
    x"3F1A2163",
    x"3F1A1C5E",
    x"3F1A175A",
    x"3F1A1255",
    x"3F1A0D51",
    x"3F1A084C",
    x"3F1A0347",
    x"3F19FE42",
    x"3F19F93D",
    x"3F19F438",
    x"3F19EF33",
    x"3F19EA2E",
    x"3F19E529",
    x"3F19E023",
    x"3F19DB1E",
    x"3F19D618",
    x"3F19D112",
    x"3F19CC0C",
    x"3F19C706",
    x"3F19C200",
    x"3F19BCFA",
    x"3F19B7F4",
    x"3F19B2EE",
    x"3F19ADE7",
    x"3F19A8E1",
    x"3F19A3DA",
    x"3F199ED4",
    x"3F1999CD",
    x"3F1994C6",
    x"3F198FBF",
    x"3F198AB8",
    x"3F1985B1",
    x"3F1980AA",
    x"3F197BA3",
    x"3F19769B",
    x"3F197194",
    x"3F196C8C",
    x"3F196784",
    x"3F19627D",
    x"3F195D75",
    x"3F19586D",
    x"3F195365",
    x"3F194E5D",
    x"3F194955",
    x"3F19444C",
    x"3F193F44",
    x"3F193A3B",
    x"3F193533",
    x"3F19302A",
    x"3F192B21",
    x"3F192618",
    x"3F19210F",
    x"3F191C06",
    x"3F1916FD",
    x"3F1911F4",
    x"3F190CEB",
    x"3F1907E1",
    x"3F1902D8",
    x"3F18FDCE",
    x"3F18F8C4",
    x"3F18F3BB",
    x"3F18EEB1",
    x"3F18E9A7",
    x"3F18E49D",
    x"3F18DF92",
    x"3F18DA88",
    x"3F18D57E",
    x"3F18D073",
    x"3F18CB69",
    x"3F18C65E",
    x"3F18C154",
    x"3F18BC49",
    x"3F18B73E",
    x"3F18B233",
    x"3F18AD28",
    x"3F18A81D",
    x"3F18A311",
    x"3F189E06",
    x"3F1898FB",
    x"3F1893EF",
    x"3F188EE3",
    x"3F1889D8",
    x"3F1884CC",
    x"3F187FC0",
    x"3F187AB4",
    x"3F1875A8",
    x"3F18709C",
    x"3F186B8F",
    x"3F186683",
    x"3F186177",
    x"3F185C6A",
    x"3F18575D",
    x"3F185251",
    x"3F184D44",
    x"3F184837",
    x"3F18432A",
    x"3F183E1D",
    x"3F183910",
    x"3F183402",
    x"3F182EF5",
    x"3F1829E7",
    x"3F1824DA",
    x"3F181FCC",
    x"3F181ABE",
    x"3F1815B1",
    x"3F1810A3",
    x"3F180B95",
    x"3F180687",
    x"3F180178",
    x"3F17FC6A",
    x"3F17F75C",
    x"3F17F24D",
    x"3F17ED3F",
    x"3F17E830",
    x"3F17E321",
    x"3F17DE12",
    x"3F17D903",
    x"3F17D3F4",
    x"3F17CEE5",
    x"3F17C9D6",
    x"3F17C4C7",
    x"3F17BFB7",
    x"3F17BAA8",
    x"3F17B598",
    x"3F17B089",
    x"3F17AB79",
    x"3F17A669",
    x"3F17A159",
    x"3F179C49",
    x"3F179739",
    x"3F179229",
    x"3F178D18",
    x"3F178808",
    x"3F1782F8",
    x"3F177DE7",
    x"3F1778D6",
    x"3F1773C6",
    x"3F176EB5",
    x"3F1769A4",
    x"3F176493",
    x"3F175F82",
    x"3F175A70",
    x"3F17555F",
    x"3F17504E",
    x"3F174B3C",
    x"3F17462B",
    x"3F174119",
    x"3F173C07",
    x"3F1736F5",
    x"3F1731E3",
    x"3F172CD1",
    x"3F1727BF",
    x"3F1722AD",
    x"3F171D9B",
    x"3F171888",
    x"3F171376",
    x"3F170E63",
    x"3F170950",
    x"3F17043E",
    x"3F16FF2B",
    x"3F16FA18",
    x"3F16F505",
    x"3F16EFF2",
    x"3F16EADE",
    x"3F16E5CB",
    x"3F16E0B8",
    x"3F16DBA4",
    x"3F16D691",
    x"3F16D17D",
    x"3F16CC69",
    x"3F16C755",
    x"3F16C241",
    x"3F16BD2D",
    x"3F16B819",
    x"3F16B305",
    x"3F16ADF1",
    x"3F16A8DC",
    x"3F16A3C8",
    x"3F169EB3",
    x"3F16999F",
    x"3F16948A",
    x"3F168F75",
    x"3F168A60",
    x"3F16854B",
    x"3F168036",
    x"3F167B21",
    x"3F16760B",
    x"3F1670F6",
    x"3F166BE0",
    x"3F1666CB",
    x"3F1661B5",
    x"3F165C9F",
    x"3F16578A",
    x"3F165274",
    x"3F164D5E",
    x"3F164847",
    x"3F164331",
    x"3F163E1B",
    x"3F163905",
    x"3F1633EE",
    x"3F162ED8",
    x"3F1629C1",
    x"3F1624AA",
    x"3F161F93",
    x"3F161A7C",
    x"3F161565",
    x"3F16104E",
    x"3F160B37",
    x"3F160620",
    x"3F160108",
    x"3F15FBF1",
    x"3F15F6D9",
    x"3F15F1C2",
    x"3F15ECAA",
    x"3F15E792",
    x"3F15E27A",
    x"3F15DD62",
    x"3F15D84A",
    x"3F15D332",
    x"3F15CE19",
    x"3F15C901",
    x"3F15C3E9",
    x"3F15BED0",
    x"3F15B9B7",
    x"3F15B49F",
    x"3F15AF86",
    x"3F15AA6D",
    x"3F15A554",
    x"3F15A03B",
    x"3F159B21",
    x"3F159608",
    x"3F1590EF",
    x"3F158BD5",
    x"3F1586BC",
    x"3F1581A2",
    x"3F157C88",
    x"3F15776F",
    x"3F157255",
    x"3F156D3B",
    x"3F156821",
    x"3F156306",
    x"3F155DEC",
    x"3F1558D2",
    x"3F1553B7",
    x"3F154E9D",
    x"3F154982",
    x"3F154467",
    x"3F153F4D",
    x"3F153A32",
    x"3F153517",
    x"3F152FFC",
    x"3F152AE0",
    x"3F1525C5",
    x"3F1520AA",
    x"3F151B8E",
    x"3F151673",
    x"3F151157",
    x"3F150C3B",
    x"3F150720",
    x"3F150204",
    x"3F14FCE8",
    x"3F14F7CC",
    x"3F14F2B0",
    x"3F14ED93",
    x"3F14E877",
    x"3F14E35A",
    x"3F14DE3E",
    x"3F14D921",
    x"3F14D405",
    x"3F14CEE8",
    x"3F14C9CB",
    x"3F14C4AE",
    x"3F14BF91",
    x"3F14BA74",
    x"3F14B557",
    x"3F14B039",
    x"3F14AB1C",
    x"3F14A5FE",
    x"3F14A0E1",
    x"3F149BC3",
    x"3F1496A5",
    x"3F149187",
    x"3F148C69",
    x"3F14874B",
    x"3F14822D",
    x"3F147D0F",
    x"3F1477F1",
    x"3F1472D2",
    x"3F146DB4",
    x"3F146895",
    x"3F146377",
    x"3F145E58",
    x"3F145939",
    x"3F14541A",
    x"3F144EFB",
    x"3F1449DC",
    x"3F1444BD",
    x"3F143F9D",
    x"3F143A7E",
    x"3F14355E",
    x"3F14303F",
    x"3F142B1F",
    x"3F142600",
    x"3F1420E0",
    x"3F141BC0",
    x"3F1416A0",
    x"3F141180",
    x"3F140C5F",
    x"3F14073F",
    x"3F14021F",
    x"3F13FCFE",
    x"3F13F7DE",
    x"3F13F2BD",
    x"3F13ED9C",
    x"3F13E87C",
    x"3F13E35B",
    x"3F13DE3A",
    x"3F13D919",
    x"3F13D3F8",
    x"3F13CED6",
    x"3F13C9B5",
    x"3F13C493",
    x"3F13BF72",
    x"3F13BA50",
    x"3F13B52F",
    x"3F13B00D",
    x"3F13AAEB",
    x"3F13A5C9",
    x"3F13A0A7",
    x"3F139B85",
    x"3F139663",
    x"3F139140",
    x"3F138C1E",
    x"3F1386FB",
    x"3F1381D9",
    x"3F137CB6",
    x"3F137793",
    x"3F137270",
    x"3F136D4D",
    x"3F13682A",
    x"3F136307",
    x"3F135DE4",
    x"3F1358C1",
    x"3F13539D",
    x"3F134E7A",
    x"3F134956",
    x"3F134433",
    x"3F133F0F",
    x"3F1339EB",
    x"3F1334C7",
    x"3F132FA3",
    x"3F132A7F",
    x"3F13255B",
    x"3F132037",
    x"3F131B12",
    x"3F1315EE",
    x"3F1310C9",
    x"3F130BA5",
    x"3F130680",
    x"3F13015B",
    x"3F12FC36",
    x"3F12F711",
    x"3F12F1EC",
    x"3F12ECC7",
    x"3F12E7A2",
    x"3F12E27C",
    x"3F12DD57",
    x"3F12D831",
    x"3F12D30C",
    x"3F12CDE6",
    x"3F12C8C0",
    x"3F12C39A",
    x"3F12BE74",
    x"3F12B94E",
    x"3F12B428",
    x"3F12AF02",
    x"3F12A9DC",
    x"3F12A4B5",
    x"3F129F8F",
    x"3F129A68",
    x"3F129542",
    x"3F12901B",
    x"3F128AF4",
    x"3F1285CD",
    x"3F1280A6",
    x"3F127B7F",
    x"3F127658",
    x"3F127130",
    x"3F126C09",
    x"3F1266E2",
    x"3F1261BA",
    x"3F125C92",
    x"3F12576B",
    x"3F125243",
    x"3F124D1B",
    x"3F1247F3",
    x"3F1242CB",
    x"3F123DA3",
    x"3F12387A",
    x"3F123352",
    x"3F122E2A",
    x"3F122901",
    x"3F1223D9",
    x"3F121EB0",
    x"3F121987",
    x"3F12145E",
    x"3F120F35",
    x"3F120A0C",
    x"3F1204E3",
    x"3F11FFBA",
    x"3F11FA91",
    x"3F11F567",
    x"3F11F03E",
    x"3F11EB14",
    x"3F11E5EA",
    x"3F11E0C1",
    x"3F11DB97",
    x"3F11D66D",
    x"3F11D143",
    x"3F11CC19",
    x"3F11C6EF",
    x"3F11C1C4",
    x"3F11BC9A",
    x"3F11B76F",
    x"3F11B245",
    x"3F11AD1A",
    x"3F11A7F0",
    x"3F11A2C5",
    x"3F119D9A",
    x"3F11986F",
    x"3F119344",
    x"3F118E19",
    x"3F1188ED",
    x"3F1183C2",
    x"3F117E97",
    x"3F11796B",
    x"3F117440",
    x"3F116F14",
    x"3F1169E8",
    x"3F1164BC",
    x"3F115F90",
    x"3F115A64",
    x"3F115538",
    x"3F11500C",
    x"3F114AE0",
    x"3F1145B3",
    x"3F114087",
    x"3F113B5A",
    x"3F11362E",
    x"3F113101",
    x"3F112BD4",
    x"3F1126A7",
    x"3F11217A",
    x"3F111C4D",
    x"3F111720",
    x"3F1111F3",
    x"3F110CC5",
    x"3F110798",
    x"3F11026A",
    x"3F10FD3D",
    x"3F10F80F",
    x"3F10F2E1",
    x"3F10EDB3",
    x"3F10E885",
    x"3F10E357",
    x"3F10DE29",
    x"3F10D8FB",
    x"3F10D3CD",
    x"3F10CE9E",
    x"3F10C970",
    x"3F10C441",
    x"3F10BF13",
    x"3F10B9E4",
    x"3F10B4B5",
    x"3F10AF86",
    x"3F10AA57",
    x"3F10A528",
    x"3F109FF9",
    x"3F109ACA",
    x"3F10959A",
    x"3F10906B",
    x"3F108B3B",
    x"3F10860C",
    x"3F1080DC",
    x"3F107BAC",
    x"3F10767C",
    x"3F10714C",
    x"3F106C1C",
    x"3F1066EC",
    x"3F1061BC",
    x"3F105C8C",
    x"3F10575B",
    x"3F10522B",
    x"3F104CFA",
    x"3F1047CA",
    x"3F104299",
    x"3F103D68",
    x"3F103837",
    x"3F103306",
    x"3F102DD5",
    x"3F1028A4",
    x"3F102373",
    x"3F101E41",
    x"3F101910",
    x"3F1013DE",
    x"3F100EAD",
    x"3F10097B",
    x"3F100449",
    x"3F0FFF17",
    x"3F0FF9E5",
    x"3F0FF4B3",
    x"3F0FEF81",
    x"3F0FEA4F",
    x"3F0FE51D",
    x"3F0FDFEA",
    x"3F0FDAB8",
    x"3F0FD585",
    x"3F0FD053",
    x"3F0FCB20",
    x"3F0FC5ED",
    x"3F0FC0BA",
    x"3F0FBB87",
    x"3F0FB654",
    x"3F0FB121",
    x"3F0FABEE",
    x"3F0FA6BA",
    x"3F0FA187",
    x"3F0F9C53",
    x"3F0F9720",
    x"3F0F91EC",
    x"3F0F8CB8",
    x"3F0F8784",
    x"3F0F8250",
    x"3F0F7D1C",
    x"3F0F77E8",
    x"3F0F72B4",
    x"3F0F6D80",
    x"3F0F684B",
    x"3F0F6317",
    x"3F0F5DE2",
    x"3F0F58AE",
    x"3F0F5379",
    x"3F0F4E44",
    x"3F0F490F",
    x"3F0F43DA",
    x"3F0F3EA5",
    x"3F0F3970",
    x"3F0F343B",
    x"3F0F2F05",
    x"3F0F29D0",
    x"3F0F249B",
    x"3F0F1F65",
    x"3F0F1A2F",
    x"3F0F14FA",
    x"3F0F0FC4",
    x"3F0F0A8E",
    x"3F0F0558",
    x"3F0F0022",
    x"3F0EFAEB",
    x"3F0EF5B5",
    x"3F0EF07F",
    x"3F0EEB48",
    x"3F0EE612",
    x"3F0EE0DB",
    x"3F0EDBA4",
    x"3F0ED66E",
    x"3F0ED137",
    x"3F0ECC00",
    x"3F0EC6C9",
    x"3F0EC192",
    x"3F0EBC5A",
    x"3F0EB723",
    x"3F0EB1EC",
    x"3F0EACB4",
    x"3F0EA77D",
    x"3F0EA245",
    x"3F0E9D0D",
    x"3F0E97D5",
    x"3F0E929D",
    x"3F0E8D65",
    x"3F0E882D",
    x"3F0E82F5",
    x"3F0E7DBD",
    x"3F0E7885",
    x"3F0E734C",
    x"3F0E6E14",
    x"3F0E68DB",
    x"3F0E63A2",
    x"3F0E5E6A",
    x"3F0E5931",
    x"3F0E53F8",
    x"3F0E4EBF",
    x"3F0E4986",
    x"3F0E444C",
    x"3F0E3F13",
    x"3F0E39DA",
    x"3F0E34A0",
    x"3F0E2F67",
    x"3F0E2A2D",
    x"3F0E24F3",
    x"3F0E1FBA",
    x"3F0E1A80",
    x"3F0E1546",
    x"3F0E100C",
    x"3F0E0AD2",
    x"3F0E0597",
    x"3F0E005D",
    x"3F0DFB23",
    x"3F0DF5E8",
    x"3F0DF0AE",
    x"3F0DEB73",
    x"3F0DE638",
    x"3F0DE0FD",
    x"3F0DDBC2",
    x"3F0DD687",
    x"3F0DD14C",
    x"3F0DCC11",
    x"3F0DC6D6",
    x"3F0DC19B",
    x"3F0DBC5F",
    x"3F0DB724",
    x"3F0DB1E8",
    x"3F0DACAC",
    x"3F0DA771",
    x"3F0DA235",
    x"3F0D9CF9",
    x"3F0D97BD",
    x"3F0D9281",
    x"3F0D8D45",
    x"3F0D8808",
    x"3F0D82CC",
    x"3F0D7D8F",
    x"3F0D7853",
    x"3F0D7316",
    x"3F0D6DDA",
    x"3F0D689D",
    x"3F0D6360",
    x"3F0D5E23",
    x"3F0D58E6",
    x"3F0D53A9",
    x"3F0D4E6C",
    x"3F0D492E",
    x"3F0D43F1",
    x"3F0D3EB3",
    x"3F0D3976",
    x"3F0D3438",
    x"3F0D2EFA",
    x"3F0D29BD",
    x"3F0D247F",
    x"3F0D1F41",
    x"3F0D1A03",
    x"3F0D14C5",
    x"3F0D0F86",
    x"3F0D0A48",
    x"3F0D050A",
    x"3F0CFFCB",
    x"3F0CFA8D",
    x"3F0CF54E",
    x"3F0CF00F",
    x"3F0CEAD0",
    x"3F0CE591",
    x"3F0CE052",
    x"3F0CDB13",
    x"3F0CD5D4",
    x"3F0CD095",
    x"3F0CCB56",
    x"3F0CC616",
    x"3F0CC0D7",
    x"3F0CBB97",
    x"3F0CB657",
    x"3F0CB118",
    x"3F0CABD8",
    x"3F0CA698",
    x"3F0CA158",
    x"3F0C9C18",
    x"3F0C96D7",
    x"3F0C9197",
    x"3F0C8C57",
    x"3F0C8716",
    x"3F0C81D6",
    x"3F0C7C95",
    x"3F0C7755",
    x"3F0C7214",
    x"3F0C6CD3",
    x"3F0C6792",
    x"3F0C6251",
    x"3F0C5D10",
    x"3F0C57CF",
    x"3F0C528D",
    x"3F0C4D4C",
    x"3F0C480B",
    x"3F0C42C9",
    x"3F0C3D87",
    x"3F0C3846",
    x"3F0C3304",
    x"3F0C2DC2",
    x"3F0C2880",
    x"3F0C233E",
    x"3F0C1DFC",
    x"3F0C18BA",
    x"3F0C1377",
    x"3F0C0E35",
    x"3F0C08F2",
    x"3F0C03B0",
    x"3F0BFE6D",
    x"3F0BF92B",
    x"3F0BF3E8",
    x"3F0BEEA5",
    x"3F0BE962",
    x"3F0BE41F",
    x"3F0BDEDC",
    x"3F0BD998",
    x"3F0BD455",
    x"3F0BCF12",
    x"3F0BC9CE",
    x"3F0BC48B",
    x"3F0BBF47",
    x"3F0BBA03",
    x"3F0BB4BF",
    x"3F0BAF7C",
    x"3F0BAA38",
    x"3F0BA4F4",
    x"3F0B9FAF",
    x"3F0B9A6B",
    x"3F0B9527",
    x"3F0B8FE2",
    x"3F0B8A9E",
    x"3F0B8559",
    x"3F0B8015",
    x"3F0B7AD0",
    x"3F0B758B",
    x"3F0B7046",
    x"3F0B6B01",
    x"3F0B65BC",
    x"3F0B6077",
    x"3F0B5B32",
    x"3F0B55EC",
    x"3F0B50A7",
    x"3F0B4B61",
    x"3F0B461C",
    x"3F0B40D6",
    x"3F0B3B90",
    x"3F0B364B",
    x"3F0B3105",
    x"3F0B2BBF",
    x"3F0B2679",
    x"3F0B2132",
    x"3F0B1BEC",
    x"3F0B16A6",
    x"3F0B115F",
    x"3F0B0C19",
    x"3F0B06D2",
    x"3F0B018C",
    x"3F0AFC45",
    x"3F0AF6FE",
    x"3F0AF1B7",
    x"3F0AEC70",
    x"3F0AE729",
    x"3F0AE1E2",
    x"3F0ADC9B",
    x"3F0AD753",
    x"3F0AD20C",
    x"3F0ACCC4",
    x"3F0AC77D",
    x"3F0AC235",
    x"3F0ABCED",
    x"3F0AB7A5",
    x"3F0AB25E",
    x"3F0AAD16",
    x"3F0AA7CD",
    x"3F0AA285",
    x"3F0A9D3D",
    x"3F0A97F5",
    x"3F0A92AC",
    x"3F0A8D64",
    x"3F0A881B",
    x"3F0A82D2",
    x"3F0A7D8A",
    x"3F0A7841",
    x"3F0A72F8",
    x"3F0A6DAF",
    x"3F0A6866",
    x"3F0A631D",
    x"3F0A5DD3",
    x"3F0A588A",
    x"3F0A5341",
    x"3F0A4DF7",
    x"3F0A48AD",
    x"3F0A4364",
    x"3F0A3E1A",
    x"3F0A38D0",
    x"3F0A3386",
    x"3F0A2E3C",
    x"3F0A28F2",
    x"3F0A23A8",
    x"3F0A1E5E",
    x"3F0A1913",
    x"3F0A13C9",
    x"3F0A0E7E",
    x"3F0A0934",
    x"3F0A03E9",
    x"3F09FE9E",
    x"3F09F954",
    x"3F09F409",
    x"3F09EEBE",
    x"3F09E973",
    x"3F09E427",
    x"3F09DEDC",
    x"3F09D991",
    x"3F09D445",
    x"3F09CEFA",
    x"3F09C9AE",
    x"3F09C463",
    x"3F09BF17",
    x"3F09B9CB",
    x"3F09B47F",
    x"3F09AF33",
    x"3F09A9E7",
    x"3F09A49B",
    x"3F099F4E",
    x"3F099A02",
    x"3F0994B6",
    x"3F098F69",
    x"3F098A1D",
    x"3F0984D0",
    x"3F097F83",
    x"3F097A36",
    x"3F0974E9",
    x"3F096F9C",
    x"3F096A4F",
    x"3F096502",
    x"3F095FB5",
    x"3F095A68",
    x"3F09551A",
    x"3F094FCD",
    x"3F094A7F",
    x"3F094531",
    x"3F093FE4",
    x"3F093A96",
    x"3F093548",
    x"3F092FFA",
    x"3F092AAC",
    x"3F09255E",
    x"3F092010",
    x"3F091AC1",
    x"3F091573",
    x"3F091024",
    x"3F090AD6",
    x"3F090587",
    x"3F090038",
    x"3F08FAEA",
    x"3F08F59B",
    x"3F08F04C",
    x"3F08EAFD",
    x"3F08E5AD",
    x"3F08E05E",
    x"3F08DB0F",
    x"3F08D5BF",
    x"3F08D070",
    x"3F08CB20",
    x"3F08C5D1",
    x"3F08C081",
    x"3F08BB31",
    x"3F08B5E1",
    x"3F08B091",
    x"3F08AB41",
    x"3F08A5F1",
    x"3F08A0A1",
    x"3F089B51",
    x"3F089600",
    x"3F0890B0",
    x"3F088B5F",
    x"3F08860F",
    x"3F0880BE",
    x"3F087B6D",
    x"3F08761C",
    x"3F0870CB",
    x"3F086B7A",
    x"3F086629",
    x"3F0860D8",
    x"3F085B87",
    x"3F085635",
    x"3F0850E4",
    x"3F084B92",
    x"3F084641",
    x"3F0840EF",
    x"3F083B9D",
    x"3F08364B",
    x"3F0830F9",
    x"3F082BA7",
    x"3F082655",
    x"3F082103",
    x"3F081BB1",
    x"3F08165E",
    x"3F08110C",
    x"3F080BB9",
    x"3F080667",
    x"3F080114",
    x"3F07FBC1",
    x"3F07F66F",
    x"3F07F11C",
    x"3F07EBC9",
    x"3F07E676",
    x"3F07E122",
    x"3F07DBCF",
    x"3F07D67C",
    x"3F07D128",
    x"3F07CBD5",
    x"3F07C681",
    x"3F07C12E",
    x"3F07BBDA",
    x"3F07B686",
    x"3F07B132",
    x"3F07ABDE",
    x"3F07A68A",
    x"3F07A136",
    x"3F079BE2",
    x"3F07968D",
    x"3F079139",
    x"3F078BE4",
    x"3F078690",
    x"3F07813B",
    x"3F077BE6",
    x"3F077692",
    x"3F07713D",
    x"3F076BE8",
    x"3F076693",
    x"3F07613E",
    x"3F075BE8",
    x"3F075693",
    x"3F07513E",
    x"3F074BE8",
    x"3F074693",
    x"3F07413D",
    x"3F073BE7",
    x"3F073692",
    x"3F07313C",
    x"3F072BE6",
    x"3F072690",
    x"3F07213A",
    x"3F071BE3",
    x"3F07168D",
    x"3F071137",
    x"3F070BE0",
    x"3F07068A",
    x"3F070133",
    x"3F06FBDD",
    x"3F06F686",
    x"3F06F12F",
    x"3F06EBD8",
    x"3F06E681",
    x"3F06E12A",
    x"3F06DBD3",
    x"3F06D67B",
    x"3F06D124",
    x"3F06CBCD",
    x"3F06C675",
    x"3F06C11E",
    x"3F06BBC6",
    x"3F06B66E",
    x"3F06B116",
    x"3F06ABBF",
    x"3F06A667",
    x"3F06A10E",
    x"3F069BB6",
    x"3F06965E",
    x"3F069106",
    x"3F068BAD",
    x"3F068655",
    x"3F0680FC",
    x"3F067BA4",
    x"3F06764B",
    x"3F0670F2",
    x"3F066B99",
    x"3F066640",
    x"3F0660E7",
    x"3F065B8E",
    x"3F065635",
    x"3F0650DC",
    x"3F064B82",
    x"3F064629",
    x"3F0640CF",
    x"3F063B76",
    x"3F06361C",
    x"3F0630C2",
    x"3F062B69",
    x"3F06260F",
    x"3F0620B5",
    x"3F061B5B",
    x"3F061600",
    x"3F0610A6",
    x"3F060B4C",
    x"3F0605F1",
    x"3F060097",
    x"3F05FB3C",
    x"3F05F5E2",
    x"3F05F087",
    x"3F05EB2C",
    x"3F05E5D1",
    x"3F05E076",
    x"3F05DB1B",
    x"3F05D5C0",
    x"3F05D065",
    x"3F05CB0A",
    x"3F05C5AE",
    x"3F05C053",
    x"3F05BAF7",
    x"3F05B59C",
    x"3F05B040",
    x"3F05AAE4",
    x"3F05A588",
    x"3F05A02C",
    x"3F059AD0",
    x"3F059574",
    x"3F059018",
    x"3F058ABC",
    x"3F05855F",
    x"3F058003",
    x"3F057AA6",
    x"3F05754A",
    x"3F056FED",
    x"3F056A90",
    x"3F056534",
    x"3F055FD7",
    x"3F055A7A",
    x"3F05551D",
    x"3F054FBF",
    x"3F054A62",
    x"3F054505",
    x"3F053FA8",
    x"3F053A4A",
    x"3F0534EC",
    x"3F052F8F",
    x"3F052A31",
    x"3F0524D3",
    x"3F051F75",
    x"3F051A18",
    x"3F0514BA",
    x"3F050F5B",
    x"3F0509FD",
    x"3F05049F",
    x"3F04FF41",
    x"3F04F9E2",
    x"3F04F484",
    x"3F04EF25",
    x"3F04E9C6",
    x"3F04E468",
    x"3F04DF09",
    x"3F04D9AA",
    x"3F04D44B",
    x"3F04CEEC",
    x"3F04C98D",
    x"3F04C42D",
    x"3F04BECE",
    x"3F04B96F",
    x"3F04B40F",
    x"3F04AEB0",
    x"3F04A950",
    x"3F04A3F0",
    x"3F049E91",
    x"3F049931",
    x"3F0493D1",
    x"3F048E71",
    x"3F048911",
    x"3F0483B0",
    x"3F047E50",
    x"3F0478F0",
    x"3F04738F",
    x"3F046E2F",
    x"3F0468CE",
    x"3F04636E",
    x"3F045E0D",
    x"3F0458AC",
    x"3F04534B",
    x"3F044DEA",
    x"3F044889",
    x"3F044328",
    x"3F043DC7",
    x"3F043865",
    x"3F043304",
    x"3F042DA2",
    x"3F042841",
    x"3F0422DF",
    x"3F041D7E",
    x"3F04181C",
    x"3F0412BA",
    x"3F040D58",
    x"3F0407F6",
    x"3F040294",
    x"3F03FD32",
    x"3F03F7CF",
    x"3F03F26D",
    x"3F03ED0B",
    x"3F03E7A8",
    x"3F03E246",
    x"3F03DCE3",
    x"3F03D780",
    x"3F03D21D",
    x"3F03CCBA",
    x"3F03C757",
    x"3F03C1F4",
    x"3F03BC91",
    x"3F03B72E",
    x"3F03B1CB",
    x"3F03AC67",
    x"3F03A704",
    x"3F03A1A0",
    x"3F039C3D",
    x"3F0396D9",
    x"3F039175",
    x"3F038C11",
    x"3F0386AE",
    x"3F03814A",
    x"3F037BE5",
    x"3F037681",
    x"3F03711D",
    x"3F036BB9",
    x"3F036654",
    x"3F0360F0",
    x"3F035B8B",
    x"3F035627",
    x"3F0350C2",
    x"3F034B5D",
    x"3F0345F8",
    x"3F034093",
    x"3F033B2E",
    x"3F0335C9",
    x"3F033064",
    x"3F032AFF",
    x"3F032599",
    x"3F032034",
    x"3F031ACE",
    x"3F031569",
    x"3F031003",
    x"3F030A9D",
    x"3F030537",
    x"3F02FFD2",
    x"3F02FA6C",
    x"3F02F506",
    x"3F02EF9F",
    x"3F02EA39",
    x"3F02E4D3",
    x"3F02DF6C",
    x"3F02DA06",
    x"3F02D49F",
    x"3F02CF39",
    x"3F02C9D2",
    x"3F02C46B",
    x"3F02BF05",
    x"3F02B99E",
    x"3F02B437",
    x"3F02AED0",
    x"3F02A968",
    x"3F02A401",
    x"3F029E9A",
    x"3F029932",
    x"3F0293CB",
    x"3F028E63",
    x"3F0288FC",
    x"3F028394",
    x"3F027E2C",
    x"3F0278C4",
    x"3F02735C",
    x"3F026DF4",
    x"3F02688C",
    x"3F026324",
    x"3F025DBC",
    x"3F025853",
    x"3F0252EB",
    x"3F024D82",
    x"3F02481A",
    x"3F0242B1",
    x"3F023D48",
    x"3F0237E0",
    x"3F023277",
    x"3F022D0E",
    x"3F0227A5",
    x"3F02223C",
    x"3F021CD2",
    x"3F021769",
    x"3F021200",
    x"3F020C96",
    x"3F02072D",
    x"3F0201C3",
    x"3F01FC59",
    x"3F01F6F0",
    x"3F01F186",
    x"3F01EC1C",
    x"3F01E6B2",
    x"3F01E148",
    x"3F01DBDE",
    x"3F01D674",
    x"3F01D109",
    x"3F01CB9F",
    x"3F01C634",
    x"3F01C0CA",
    x"3F01BB5F",
    x"3F01B5F5",
    x"3F01B08A",
    x"3F01AB1F",
    x"3F01A5B4",
    x"3F01A049",
    x"3F019ADE",
    x"3F019573",
    x"3F019007",
    x"3F018A9C",
    x"3F018531",
    x"3F017FC5",
    x"3F017A5A",
    x"3F0174EE",
    x"3F016F82",
    x"3F016A17",
    x"3F0164AB",
    x"3F015F3F",
    x"3F0159D3",
    x"3F015467",
    x"3F014EFA",
    x"3F01498E",
    x"3F014422",
    x"3F013EB5",
    x"3F013949",
    x"3F0133DC",
    x"3F012E70",
    x"3F012903",
    x"3F012396",
    x"3F011E29",
    x"3F0118BC",
    x"3F01134F",
    x"3F010DE2",
    x"3F010875",
    x"3F010308",
    x"3F00FD9A",
    x"3F00F82D",
    x"3F00F2BF",
    x"3F00ED52",
    x"3F00E7E4",
    x"3F00E276",
    x"3F00DD09",
    x"3F00D79B",
    x"3F00D22D",
    x"3F00CCBF",
    x"3F00C751",
    x"3F00C1E2",
    x"3F00BC74",
    x"3F00B706",
    x"3F00B197",
    x"3F00AC29",
    x"3F00A6BA",
    x"3F00A14C",
    x"3F009BDD",
    x"3F00966E",
    x"3F0090FF",
    x"3F008B90",
    x"3F008621",
    x"3F0080B2",
    x"3F007B43",
    x"3F0075D4",
    x"3F007064",
    x"3F006AF5",
    x"3F006585",
    x"3F006016",
    x"3F005AA6",
    x"3F005536",
    x"3F004FC6",
    x"3F004A56",
    x"3F0044E6",
    x"3F003F76",
    x"3F003A06",
    x"3F003496",
    x"3F002F26",
    x"3F0029B5",
    x"3F002445",
    x"3F001ED4",
    x"3F001964",
    x"3F0013F3",
    x"3F000E82",
    x"3F000912",
    x"3F0003A1",
    x"3EFFFC5F",
    x"3EFFF17D",
    x"3EFFE69B",
    x"3EFFDBB8",
    x"3EFFD0D6",
    x"3EFFC5F3",
    x"3EFFBB10",
    x"3EFFB02D",
    x"3EFFA54A",
    x"3EFF9A67",
    x"3EFF8F83",
    x"3EFF849F",
    x"3EFF79BC",
    x"3EFF6ED8",
    x"3EFF63F4",
    x"3EFF590F",
    x"3EFF4E2B",
    x"3EFF4346",
    x"3EFF3862",
    x"3EFF2D7D",
    x"3EFF2298",
    x"3EFF17B2",
    x"3EFF0CCD",
    x"3EFF01E8",
    x"3EFEF702",
    x"3EFEEC1C",
    x"3EFEE136",
    x"3EFED650",
    x"3EFECB6A",
    x"3EFEC083",
    x"3EFEB59D",
    x"3EFEAAB6",
    x"3EFE9FCF",
    x"3EFE94E8",
    x"3EFE8A01",
    x"3EFE7F19",
    x"3EFE7432",
    x"3EFE694A",
    x"3EFE5E62",
    x"3EFE537A",
    x"3EFE4892",
    x"3EFE3DAA",
    x"3EFE32C2",
    x"3EFE27D9",
    x"3EFE1CF0",
    x"3EFE1207",
    x"3EFE071E",
    x"3EFDFC35",
    x"3EFDF14C",
    x"3EFDE662",
    x"3EFDDB79",
    x"3EFDD08F",
    x"3EFDC5A5",
    x"3EFDBABB",
    x"3EFDAFD1",
    x"3EFDA4E6",
    x"3EFD99FC",
    x"3EFD8F11",
    x"3EFD8426",
    x"3EFD793B",
    x"3EFD6E50",
    x"3EFD6365",
    x"3EFD5879",
    x"3EFD4D8D",
    x"3EFD42A2",
    x"3EFD37B6",
    x"3EFD2CCA",
    x"3EFD21DD",
    x"3EFD16F1",
    x"3EFD0C04",
    x"3EFD0118",
    x"3EFCF62B",
    x"3EFCEB3E",
    x"3EFCE051",
    x"3EFCD563",
    x"3EFCCA76",
    x"3EFCBF88",
    x"3EFCB49B",
    x"3EFCA9AD",
    x"3EFC9EBF",
    x"3EFC93D0",
    x"3EFC88E2",
    x"3EFC7DF3",
    x"3EFC7305",
    x"3EFC6816",
    x"3EFC5D27",
    x"3EFC5238",
    x"3EFC4748",
    x"3EFC3C59",
    x"3EFC3169",
    x"3EFC267A",
    x"3EFC1B8A",
    x"3EFC109A",
    x"3EFC05AA",
    x"3EFBFAB9",
    x"3EFBEFC9",
    x"3EFBE4D8",
    x"3EFBD9E7",
    x"3EFBCEF6",
    x"3EFBC405",
    x"3EFBB914",
    x"3EFBAE22",
    x"3EFBA331",
    x"3EFB983F",
    x"3EFB8D4D",
    x"3EFB825B",
    x"3EFB7769",
    x"3EFB6C77",
    x"3EFB6184",
    x"3EFB5692",
    x"3EFB4B9F",
    x"3EFB40AC",
    x"3EFB35B9",
    x"3EFB2AC6",
    x"3EFB1FD2",
    x"3EFB14DF",
    x"3EFB09EB",
    x"3EFAFEF7",
    x"3EFAF403",
    x"3EFAE90F",
    x"3EFADE1B",
    x"3EFAD326",
    x"3EFAC832",
    x"3EFABD3D",
    x"3EFAB248",
    x"3EFAA753",
    x"3EFA9C5E",
    x"3EFA9169",
    x"3EFA8673",
    x"3EFA7B7D",
    x"3EFA7088",
    x"3EFA6592",
    x"3EFA5A9C",
    x"3EFA4FA5",
    x"3EFA44AF",
    x"3EFA39B8",
    x"3EFA2EC2",
    x"3EFA23CB",
    x"3EFA18D4",
    x"3EFA0DDD",
    x"3EFA02E5",
    x"3EF9F7EE",
    x"3EF9ECF6",
    x"3EF9E1FE",
    x"3EF9D707",
    x"3EF9CC0E",
    x"3EF9C116",
    x"3EF9B61E",
    x"3EF9AB25",
    x"3EF9A02D",
    x"3EF99534",
    x"3EF98A3B",
    x"3EF97F42",
    x"3EF97449",
    x"3EF9694F",
    x"3EF95E56",
    x"3EF9535C",
    x"3EF94862",
    x"3EF93D68",
    x"3EF9326E",
    x"3EF92773",
    x"3EF91C79",
    x"3EF9117E",
    x"3EF90684",
    x"3EF8FB89",
    x"3EF8F08E",
    x"3EF8E592",
    x"3EF8DA97",
    x"3EF8CF9C",
    x"3EF8C4A0",
    x"3EF8B9A4",
    x"3EF8AEA8",
    x"3EF8A3AC",
    x"3EF898B0",
    x"3EF88DB3",
    x"3EF882B7",
    x"3EF877BA",
    x"3EF86CBD",
    x"3EF861C0",
    x"3EF856C3",
    x"3EF84BC6",
    x"3EF840C8",
    x"3EF835CB",
    x"3EF82ACD",
    x"3EF81FCF",
    x"3EF814D1",
    x"3EF809D3",
    x"3EF7FED4",
    x"3EF7F3D6",
    x"3EF7E8D7",
    x"3EF7DDD8",
    x"3EF7D2D9",
    x"3EF7C7DA",
    x"3EF7BCDB",
    x"3EF7B1DC",
    x"3EF7A6DC",
    x"3EF79BDC",
    x"3EF790DC",
    x"3EF785DC",
    x"3EF77ADC",
    x"3EF76FDC",
    x"3EF764DC",
    x"3EF759DB",
    x"3EF74EDA",
    x"3EF743D9",
    x"3EF738D8",
    x"3EF72DD7",
    x"3EF722D6",
    x"3EF717D4",
    x"3EF70CD3",
    x"3EF701D1",
    x"3EF6F6CF",
    x"3EF6EBCD",
    x"3EF6E0CB",
    x"3EF6D5C8",
    x"3EF6CAC6",
    x"3EF6BFC3",
    x"3EF6B4C0",
    x"3EF6A9BD",
    x"3EF69EBA",
    x"3EF693B7",
    x"3EF688B3",
    x"3EF67DB0",
    x"3EF672AC",
    x"3EF667A8",
    x"3EF65CA4",
    x"3EF651A0",
    x"3EF6469C",
    x"3EF63B97",
    x"3EF63093",
    x"3EF6258E",
    x"3EF61A89",
    x"3EF60F84",
    x"3EF6047F",
    x"3EF5F979",
    x"3EF5EE74",
    x"3EF5E36E",
    x"3EF5D868",
    x"3EF5CD62",
    x"3EF5C25C",
    x"3EF5B756",
    x"3EF5AC50",
    x"3EF5A149",
    x"3EF59643",
    x"3EF58B3C",
    x"3EF58035",
    x"3EF5752E",
    x"3EF56A26",
    x"3EF55F1F",
    x"3EF55417",
    x"3EF54910",
    x"3EF53E08",
    x"3EF53300",
    x"3EF527F8",
    x"3EF51CEF",
    x"3EF511E7",
    x"3EF506DE",
    x"3EF4FBD5",
    x"3EF4F0CC",
    x"3EF4E5C3",
    x"3EF4DABA",
    x"3EF4CFB1",
    x"3EF4C4A7",
    x"3EF4B99E",
    x"3EF4AE94",
    x"3EF4A38A",
    x"3EF49880",
    x"3EF48D76",
    x"3EF4826B",
    x"3EF47761",
    x"3EF46C56",
    x"3EF4614B",
    x"3EF45640",
    x"3EF44B35",
    x"3EF4402A",
    x"3EF4351F",
    x"3EF42A13",
    x"3EF41F07",
    x"3EF413FB",
    x"3EF408F0",
    x"3EF3FDE3",
    x"3EF3F2D7",
    x"3EF3E7CB",
    x"3EF3DCBE",
    x"3EF3D1B1",
    x"3EF3C6A4",
    x"3EF3BB97",
    x"3EF3B08A",
    x"3EF3A57D",
    x"3EF39A6F",
    x"3EF38F62",
    x"3EF38454",
    x"3EF37946",
    x"3EF36E38",
    x"3EF3632A",
    x"3EF3581C",
    x"3EF34D0D",
    x"3EF341FE",
    x"3EF336F0",
    x"3EF32BE1",
    x"3EF320D2",
    x"3EF315C2",
    x"3EF30AB3",
    x"3EF2FFA4",
    x"3EF2F494",
    x"3EF2E984",
    x"3EF2DE74",
    x"3EF2D364",
    x"3EF2C854",
    x"3EF2BD43",
    x"3EF2B233",
    x"3EF2A722",
    x"3EF29C11",
    x"3EF29100",
    x"3EF285EF",
    x"3EF27ADE",
    x"3EF26FCD",
    x"3EF264BB",
    x"3EF259A9",
    x"3EF24E97",
    x"3EF24385",
    x"3EF23873",
    x"3EF22D61",
    x"3EF2224F",
    x"3EF2173C",
    x"3EF20C29",
    x"3EF20116",
    x"3EF1F603",
    x"3EF1EAF0",
    x"3EF1DFDD",
    x"3EF1D4C9",
    x"3EF1C9B6",
    x"3EF1BEA2",
    x"3EF1B38E",
    x"3EF1A87A",
    x"3EF19D66",
    x"3EF19252",
    x"3EF1873D",
    x"3EF17C28",
    x"3EF17114",
    x"3EF165FF",
    x"3EF15AEA",
    x"3EF14FD5",
    x"3EF144BF",
    x"3EF139AA",
    x"3EF12E94",
    x"3EF1237E",
    x"3EF11868",
    x"3EF10D52",
    x"3EF1023C",
    x"3EF0F726",
    x"3EF0EC0F",
    x"3EF0E0F9",
    x"3EF0D5E2",
    x"3EF0CACB",
    x"3EF0BFB4",
    x"3EF0B49C",
    x"3EF0A985",
    x"3EF09E6E",
    x"3EF09356",
    x"3EF0883E",
    x"3EF07D26",
    x"3EF0720E",
    x"3EF066F6",
    x"3EF05BDD",
    x"3EF050C5",
    x"3EF045AC",
    x"3EF03A93",
    x"3EF02F7A",
    x"3EF02461",
    x"3EF01948",
    x"3EF00E2E",
    x"3EF00315",
    x"3EEFF7FB",
    x"3EEFECE1",
    x"3EEFE1C7",
    x"3EEFD6AD",
    x"3EEFCB93",
    x"3EEFC079",
    x"3EEFB55E",
    x"3EEFAA43",
    x"3EEF9F28",
    x"3EEF940D",
    x"3EEF88F2",
    x"3EEF7DD7",
    x"3EEF72BC",
    x"3EEF67A0",
    x"3EEF5C84",
    x"3EEF5168",
    x"3EEF464C",
    x"3EEF3B30",
    x"3EEF3014",
    x"3EEF24F7",
    x"3EEF19DB",
    x"3EEF0EBE",
    x"3EEF03A1",
    x"3EEEF884",
    x"3EEEED67",
    x"3EEEE24A",
    x"3EEED72C",
    x"3EEECC0F",
    x"3EEEC0F1",
    x"3EEEB5D3",
    x"3EEEAAB5",
    x"3EEE9F97",
    x"3EEE9479",
    x"3EEE895A",
    x"3EEE7E3C",
    x"3EEE731D",
    x"3EEE67FE",
    x"3EEE5CDF",
    x"3EEE51C0",
    x"3EEE46A0",
    x"3EEE3B81",
    x"3EEE3061",
    x"3EEE2542",
    x"3EEE1A22",
    x"3EEE0F02",
    x"3EEE03E2",
    x"3EEDF8C1",
    x"3EEDEDA1",
    x"3EEDE280",
    x"3EEDD75F",
    x"3EEDCC3E",
    x"3EEDC11D",
    x"3EEDB5FC",
    x"3EEDAADB",
    x"3EED9FB9",
    x"3EED9498",
    x"3EED8976",
    x"3EED7E54",
    x"3EED7332",
    x"3EED6810",
    x"3EED5CEE",
    x"3EED51CB",
    x"3EED46A9",
    x"3EED3B86",
    x"3EED3063",
    x"3EED2540",
    x"3EED1A1D",
    x"3EED0EF9",
    x"3EED03D6",
    x"3EECF8B2",
    x"3EECED8F",
    x"3EECE26B",
    x"3EECD747",
    x"3EECCC22",
    x"3EECC0FE",
    x"3EECB5DA",
    x"3EECAAB5",
    x"3EEC9F90",
    x"3EEC946B",
    x"3EEC8946",
    x"3EEC7E21",
    x"3EEC72FC",
    x"3EEC67D6",
    x"3EEC5CB1",
    x"3EEC518B",
    x"3EEC4665",
    x"3EEC3B3F",
    x"3EEC3019",
    x"3EEC24F3",
    x"3EEC19CC",
    x"3EEC0EA5",
    x"3EEC037F",
    x"3EEBF858",
    x"3EEBED31",
    x"3EEBE20A",
    x"3EEBD6E2",
    x"3EEBCBBB",
    x"3EEBC093",
    x"3EEBB56C",
    x"3EEBAA44",
    x"3EEB9F1C",
    x"3EEB93F3",
    x"3EEB88CB",
    x"3EEB7DA3",
    x"3EEB727A",
    x"3EEB6751",
    x"3EEB5C28",
    x"3EEB50FF",
    x"3EEB45D6",
    x"3EEB3AAD",
    x"3EEB2F84",
    x"3EEB245A",
    x"3EEB1930",
    x"3EEB0E06",
    x"3EEB02DC",
    x"3EEAF7B2",
    x"3EEAEC88",
    x"3EEAE15D",
    x"3EEAD633",
    x"3EEACB08",
    x"3EEABFDD",
    x"3EEAB4B2",
    x"3EEAA987",
    x"3EEA9E5C",
    x"3EEA9330",
    x"3EEA8805",
    x"3EEA7CD9",
    x"3EEA71AD",
    x"3EEA6681",
    x"3EEA5B55",
    x"3EEA5029",
    x"3EEA44FD",
    x"3EEA39D0",
    x"3EEA2EA3",
    x"3EEA2376",
    x"3EEA1849",
    x"3EEA0D1C",
    x"3EEA01EF",
    x"3EE9F6C2",
    x"3EE9EB94",
    x"3EE9E066",
    x"3EE9D539",
    x"3EE9CA0B",
    x"3EE9BEDD",
    x"3EE9B3AE",
    x"3EE9A880",
    x"3EE99D51",
    x"3EE99223",
    x"3EE986F4",
    x"3EE97BC5",
    x"3EE97096",
    x"3EE96567",
    x"3EE95A37",
    x"3EE94F08",
    x"3EE943D8",
    x"3EE938A8",
    x"3EE92D78",
    x"3EE92248",
    x"3EE91718",
    x"3EE90BE8",
    x"3EE900B7",
    x"3EE8F587",
    x"3EE8EA56",
    x"3EE8DF25",
    x"3EE8D3F4",
    x"3EE8C8C3",
    x"3EE8BD91",
    x"3EE8B260",
    x"3EE8A72E",
    x"3EE89BFD",
    x"3EE890CB",
    x"3EE88599",
    x"3EE87A66",
    x"3EE86F34",
    x"3EE86402",
    x"3EE858CF",
    x"3EE84D9C",
    x"3EE84269",
    x"3EE83736",
    x"3EE82C03",
    x"3EE820D0",
    x"3EE8159C",
    x"3EE80A69",
    x"3EE7FF35",
    x"3EE7F401",
    x"3EE7E8CD",
    x"3EE7DD99",
    x"3EE7D265",
    x"3EE7C731",
    x"3EE7BBFC",
    x"3EE7B0C7",
    x"3EE7A592",
    x"3EE79A5D",
    x"3EE78F28",
    x"3EE783F3",
    x"3EE778BE",
    x"3EE76D88",
    x"3EE76253",
    x"3EE7571D",
    x"3EE74BE7",
    x"3EE740B1",
    x"3EE7357A",
    x"3EE72A44",
    x"3EE71F0E",
    x"3EE713D7",
    x"3EE708A0",
    x"3EE6FD69",
    x"3EE6F232",
    x"3EE6E6FB",
    x"3EE6DBC4",
    x"3EE6D08C",
    x"3EE6C554",
    x"3EE6BA1D",
    x"3EE6AEE5",
    x"3EE6A3AD",
    x"3EE69875",
    x"3EE68D3C",
    x"3EE68204",
    x"3EE676CB",
    x"3EE66B93",
    x"3EE6605A",
    x"3EE65521",
    x"3EE649E7",
    x"3EE63EAE",
    x"3EE63375",
    x"3EE6283B",
    x"3EE61D02",
    x"3EE611C8",
    x"3EE6068E",
    x"3EE5FB54",
    x"3EE5F019",
    x"3EE5E4DF",
    x"3EE5D9A4",
    x"3EE5CE6A",
    x"3EE5C32F",
    x"3EE5B7F4",
    x"3EE5ACB9",
    x"3EE5A17E",
    x"3EE59642",
    x"3EE58B07",
    x"3EE57FCB",
    x"3EE5748F",
    x"3EE56953",
    x"3EE55E17",
    x"3EE552DB",
    x"3EE5479F",
    x"3EE53C62",
    x"3EE53126",
    x"3EE525E9",
    x"3EE51AAC",
    x"3EE50F6F",
    x"3EE50432",
    x"3EE4F8F5",
    x"3EE4EDB7",
    x"3EE4E27A",
    x"3EE4D73C",
    x"3EE4CBFE",
    x"3EE4C0C0",
    x"3EE4B582",
    x"3EE4AA44",
    x"3EE49F05",
    x"3EE493C7",
    x"3EE48888",
    x"3EE47D49",
    x"3EE4720A",
    x"3EE466CB",
    x"3EE45B8C",
    x"3EE4504D",
    x"3EE4450D",
    x"3EE439CE",
    x"3EE42E8E",
    x"3EE4234E",
    x"3EE4180E",
    x"3EE40CCE",
    x"3EE4018D",
    x"3EE3F64D",
    x"3EE3EB0C",
    x"3EE3DFCB",
    x"3EE3D48B",
    x"3EE3C94A",
    x"3EE3BE08",
    x"3EE3B2C7",
    x"3EE3A786",
    x"3EE39C44",
    x"3EE39102",
    x"3EE385C1",
    x"3EE37A7F",
    x"3EE36F3D",
    x"3EE363FA",
    x"3EE358B8",
    x"3EE34D75",
    x"3EE34233",
    x"3EE336F0",
    x"3EE32BAD",
    x"3EE3206A",
    x"3EE31527",
    x"3EE309E3",
    x"3EE2FEA0",
    x"3EE2F35C",
    x"3EE2E819",
    x"3EE2DCD5",
    x"3EE2D191",
    x"3EE2C64C",
    x"3EE2BB08",
    x"3EE2AFC4",
    x"3EE2A47F",
    x"3EE2993A",
    x"3EE28DF6",
    x"3EE282B1",
    x"3EE2776C",
    x"3EE26C26",
    x"3EE260E1",
    x"3EE2559B",
    x"3EE24A56",
    x"3EE23F10",
    x"3EE233CA",
    x"3EE22884",
    x"3EE21D3E",
    x"3EE211F7",
    x"3EE206B1",
    x"3EE1FB6A",
    x"3EE1F023",
    x"3EE1E4DD",
    x"3EE1D996",
    x"3EE1CE4E",
    x"3EE1C307",
    x"3EE1B7C0",
    x"3EE1AC78",
    x"3EE1A130",
    x"3EE195E9",
    x"3EE18AA1",
    x"3EE17F58",
    x"3EE17410",
    x"3EE168C8",
    x"3EE15D7F",
    x"3EE15237",
    x"3EE146EE",
    x"3EE13BA5",
    x"3EE1305C",
    x"3EE12513",
    x"3EE119C9",
    x"3EE10E80",
    x"3EE10336",
    x"3EE0F7ED",
    x"3EE0ECA3",
    x"3EE0E159",
    x"3EE0D60E",
    x"3EE0CAC4",
    x"3EE0BF7A",
    x"3EE0B42F",
    x"3EE0A8E5",
    x"3EE09D9A",
    x"3EE0924F",
    x"3EE08704",
    x"3EE07BB8",
    x"3EE0706D",
    x"3EE06522",
    x"3EE059D6",
    x"3EE04E8A",
    x"3EE0433E",
    x"3EE037F2",
    x"3EE02CA6",
    x"3EE0215A",
    x"3EE0160D",
    x"3EE00AC1",
    x"3EDFFF74",
    x"3EDFF427",
    x"3EDFE8DA",
    x"3EDFDD8D",
    x"3EDFD240",
    x"3EDFC6F2",
    x"3EDFBBA5",
    x"3EDFB057",
    x"3EDFA509",
    x"3EDF99BB",
    x"3EDF8E6D",
    x"3EDF831F",
    x"3EDF77D1",
    x"3EDF6C82",
    x"3EDF6134",
    x"3EDF55E5",
    x"3EDF4A96",
    x"3EDF3F47",
    x"3EDF33F8",
    x"3EDF28A9",
    x"3EDF1D59",
    x"3EDF120A",
    x"3EDF06BA",
    x"3EDEFB6A",
    x"3EDEF01A",
    x"3EDEE4CA",
    x"3EDED97A",
    x"3EDECE2A",
    x"3EDEC2D9",
    x"3EDEB789",
    x"3EDEAC38",
    x"3EDEA0E7",
    x"3EDE9596",
    x"3EDE8A45",
    x"3EDE7EF3",
    x"3EDE73A2",
    x"3EDE6851",
    x"3EDE5CFF",
    x"3EDE51AD",
    x"3EDE465B",
    x"3EDE3B09",
    x"3EDE2FB7",
    x"3EDE2464",
    x"3EDE1912",
    x"3EDE0DBF",
    x"3EDE026C",
    x"3EDDF71A",
    x"3EDDEBC7",
    x"3EDDE073",
    x"3EDDD520",
    x"3EDDC9CD",
    x"3EDDBE79",
    x"3EDDB325",
    x"3EDDA7D2",
    x"3EDD9C7E",
    x"3EDD912A",
    x"3EDD85D5",
    x"3EDD7A81",
    x"3EDD6F2C",
    x"3EDD63D8",
    x"3EDD5883",
    x"3EDD4D2E",
    x"3EDD41D9",
    x"3EDD3684",
    x"3EDD2B2F",
    x"3EDD1FD9",
    x"3EDD1484",
    x"3EDD092E",
    x"3EDCFDD8",
    x"3EDCF282",
    x"3EDCE72C",
    x"3EDCDBD6",
    x"3EDCD07F",
    x"3EDCC529",
    x"3EDCB9D2",
    x"3EDCAE7C",
    x"3EDCA325",
    x"3EDC97CE",
    x"3EDC8C76",
    x"3EDC811F",
    x"3EDC75C8",
    x"3EDC6A70",
    x"3EDC5F18",
    x"3EDC53C1",
    x"3EDC4869",
    x"3EDC3D11",
    x"3EDC31B8",
    x"3EDC2660",
    x"3EDC1B08",
    x"3EDC0FAF",
    x"3EDC0456",
    x"3EDBF8FD",
    x"3EDBEDA4",
    x"3EDBE24B",
    x"3EDBD6F2",
    x"3EDBCB98",
    x"3EDBC03F",
    x"3EDBB4E5",
    x"3EDBA98B",
    x"3EDB9E31",
    x"3EDB92D7",
    x"3EDB877D",
    x"3EDB7C23",
    x"3EDB70C8",
    x"3EDB656E",
    x"3EDB5A13",
    x"3EDB4EB8",
    x"3EDB435D",
    x"3EDB3802",
    x"3EDB2CA7",
    x"3EDB214B",
    x"3EDB15F0",
    x"3EDB0A94",
    x"3EDAFF38",
    x"3EDAF3DC",
    x"3EDAE880",
    x"3EDADD24",
    x"3EDAD1C8",
    x"3EDAC66B",
    x"3EDABB0F",
    x"3EDAAFB2",
    x"3EDAA455",
    x"3EDA98F8",
    x"3EDA8D9B",
    x"3EDA823E",
    x"3EDA76E0",
    x"3EDA6B83",
    x"3EDA6025",
    x"3EDA54C8",
    x"3EDA496A",
    x"3EDA3E0C",
    x"3EDA32AD",
    x"3EDA274F",
    x"3EDA1BF1",
    x"3EDA1092",
    x"3EDA0533",
    x"3ED9F9D5",
    x"3ED9EE76",
    x"3ED9E317",
    x"3ED9D7B7",
    x"3ED9CC58",
    x"3ED9C0F9",
    x"3ED9B599",
    x"3ED9AA39",
    x"3ED99ED9",
    x"3ED99379",
    x"3ED98819",
    x"3ED97CB9",
    x"3ED97159",
    x"3ED965F8",
    x"3ED95A97",
    x"3ED94F37",
    x"3ED943D6",
    x"3ED93875",
    x"3ED92D13",
    x"3ED921B2",
    x"3ED91651",
    x"3ED90AEF",
    x"3ED8FF8D",
    x"3ED8F42C",
    x"3ED8E8CA",
    x"3ED8DD67",
    x"3ED8D205",
    x"3ED8C6A3",
    x"3ED8BB40",
    x"3ED8AFDE",
    x"3ED8A47B",
    x"3ED89918",
    x"3ED88DB5",
    x"3ED88252",
    x"3ED876EF",
    x"3ED86B8B",
    x"3ED86028",
    x"3ED854C4",
    x"3ED84960",
    x"3ED83DFC",
    x"3ED83298",
    x"3ED82734",
    x"3ED81BD0",
    x"3ED8106B",
    x"3ED80507",
    x"3ED7F9A2",
    x"3ED7EE3D",
    x"3ED7E2D8",
    x"3ED7D773",
    x"3ED7CC0E",
    x"3ED7C0A9",
    x"3ED7B543",
    x"3ED7A9DE",
    x"3ED79E78",
    x"3ED79312",
    x"3ED787AC",
    x"3ED77C46",
    x"3ED770E0",
    x"3ED76579",
    x"3ED75A13",
    x"3ED74EAC",
    x"3ED74345",
    x"3ED737DE",
    x"3ED72C77",
    x"3ED72110",
    x"3ED715A9",
    x"3ED70A41",
    x"3ED6FEDA",
    x"3ED6F372",
    x"3ED6E80A",
    x"3ED6DCA2",
    x"3ED6D13A",
    x"3ED6C5D2",
    x"3ED6BA6A",
    x"3ED6AF01",
    x"3ED6A399",
    x"3ED69830",
    x"3ED68CC7",
    x"3ED6815E",
    x"3ED675F5",
    x"3ED66A8C",
    x"3ED65F22",
    x"3ED653B9",
    x"3ED6484F",
    x"3ED63CE5",
    x"3ED6317B",
    x"3ED62611",
    x"3ED61AA7",
    x"3ED60F3D",
    x"3ED603D3",
    x"3ED5F868",
    x"3ED5ECFD",
    x"3ED5E193",
    x"3ED5D628",
    x"3ED5CABD",
    x"3ED5BF52",
    x"3ED5B3E6",
    x"3ED5A87B",
    x"3ED59D0F",
    x"3ED591A4",
    x"3ED58638",
    x"3ED57ACC",
    x"3ED56F60",
    x"3ED563F3",
    x"3ED55887",
    x"3ED54D1B",
    x"3ED541AE",
    x"3ED53641",
    x"3ED52AD5",
    x"3ED51F68",
    x"3ED513FA",
    x"3ED5088D",
    x"3ED4FD20",
    x"3ED4F1B2",
    x"3ED4E645",
    x"3ED4DAD7",
    x"3ED4CF69",
    x"3ED4C3FB",
    x"3ED4B88D",
    x"3ED4AD1F",
    x"3ED4A1B0",
    x"3ED49642",
    x"3ED48AD3",
    x"3ED47F64",
    x"3ED473F5",
    x"3ED46886",
    x"3ED45D17",
    x"3ED451A8",
    x"3ED44639",
    x"3ED43AC9",
    x"3ED42F59",
    x"3ED423EA",
    x"3ED4187A",
    x"3ED40D0A",
    x"3ED40199",
    x"3ED3F629",
    x"3ED3EAB9",
    x"3ED3DF48",
    x"3ED3D3D7",
    x"3ED3C867",
    x"3ED3BCF6",
    x"3ED3B185",
    x"3ED3A613",
    x"3ED39AA2",
    x"3ED38F31",
    x"3ED383BF",
    x"3ED3784D",
    x"3ED36CDB",
    x"3ED3616A",
    x"3ED355F7",
    x"3ED34A85",
    x"3ED33F13",
    x"3ED333A0",
    x"3ED3282E",
    x"3ED31CBB",
    x"3ED31148",
    x"3ED305D5",
    x"3ED2FA62",
    x"3ED2EEEF",
    x"3ED2E37C",
    x"3ED2D808",
    x"3ED2CC94",
    x"3ED2C121",
    x"3ED2B5AD",
    x"3ED2AA39",
    x"3ED29EC5",
    x"3ED29350",
    x"3ED287DC",
    x"3ED27C68",
    x"3ED270F3",
    x"3ED2657E",
    x"3ED25A09",
    x"3ED24E94",
    x"3ED2431F",
    x"3ED237AA",
    x"3ED22C34",
    x"3ED220BF",
    x"3ED21549",
    x"3ED209D3",
    x"3ED1FE5E",
    x"3ED1F2E8",
    x"3ED1E771",
    x"3ED1DBFB",
    x"3ED1D085",
    x"3ED1C50E",
    x"3ED1B998",
    x"3ED1AE21",
    x"3ED1A2AA",
    x"3ED19733",
    x"3ED18BBC",
    x"3ED18044",
    x"3ED174CD",
    x"3ED16955",
    x"3ED15DDE",
    x"3ED15266",
    x"3ED146EE",
    x"3ED13B76",
    x"3ED12FFE",
    x"3ED12485",
    x"3ED1190D",
    x"3ED10D95",
    x"3ED1021C",
    x"3ED0F6A3",
    x"3ED0EB2A",
    x"3ED0DFB1",
    x"3ED0D438",
    x"3ED0C8BF",
    x"3ED0BD45",
    x"3ED0B1CC",
    x"3ED0A652",
    x"3ED09AD8",
    x"3ED08F5E",
    x"3ED083E4",
    x"3ED0786A",
    x"3ED06CF0",
    x"3ED06175",
    x"3ED055FB",
    x"3ED04A80",
    x"3ED03F05",
    x"3ED0338A",
    x"3ED0280F",
    x"3ED01C94",
    x"3ED01119",
    x"3ED0059D",
    x"3ECFFA22",
    x"3ECFEEA6",
    x"3ECFE32A",
    x"3ECFD7AE",
    x"3ECFCC32",
    x"3ECFC0B6",
    x"3ECFB53A",
    x"3ECFA9BD",
    x"3ECF9E41",
    x"3ECF92C4",
    x"3ECF8747",
    x"3ECF7BCA",
    x"3ECF704D",
    x"3ECF64D0",
    x"3ECF5953",
    x"3ECF4DD5",
    x"3ECF4258",
    x"3ECF36DA",
    x"3ECF2B5C",
    x"3ECF1FDE",
    x"3ECF1460",
    x"3ECF08E2",
    x"3ECEFD64",
    x"3ECEF1E5",
    x"3ECEE667",
    x"3ECEDAE8",
    x"3ECECF69",
    x"3ECEC3EA",
    x"3ECEB86B",
    x"3ECEACEC",
    x"3ECEA16D",
    x"3ECE95ED",
    x"3ECE8A6E",
    x"3ECE7EEE",
    x"3ECE736E",
    x"3ECE67EE",
    x"3ECE5C6E",
    x"3ECE50EE",
    x"3ECE456E",
    x"3ECE39ED",
    x"3ECE2E6D",
    x"3ECE22EC",
    x"3ECE176B",
    x"3ECE0BEA",
    x"3ECE0069",
    x"3ECDF4E8",
    x"3ECDE967",
    x"3ECDDDE5",
    x"3ECDD264",
    x"3ECDC6E2",
    x"3ECDBB60",
    x"3ECDAFDE",
    x"3ECDA45C",
    x"3ECD98DA",
    x"3ECD8D58",
    x"3ECD81D5",
    x"3ECD7653",
    x"3ECD6AD0",
    x"3ECD5F4D",
    x"3ECD53CA",
    x"3ECD4847",
    x"3ECD3CC4",
    x"3ECD3141",
    x"3ECD25BE",
    x"3ECD1A3A",
    x"3ECD0EB6",
    x"3ECD0333",
    x"3ECCF7AF",
    x"3ECCEC2B",
    x"3ECCE0A7",
    x"3ECCD522",
    x"3ECCC99E",
    x"3ECCBE19",
    x"3ECCB295",
    x"3ECCA710",
    x"3ECC9B8B",
    x"3ECC9006",
    x"3ECC8481",
    x"3ECC78FC",
    x"3ECC6D76",
    x"3ECC61F1",
    x"3ECC566B",
    x"3ECC4AE5",
    x"3ECC3F60",
    x"3ECC33DA",
    x"3ECC2853",
    x"3ECC1CCD",
    x"3ECC1147",
    x"3ECC05C0",
    x"3ECBFA3A",
    x"3ECBEEB3",
    x"3ECBE32C",
    x"3ECBD7A5",
    x"3ECBCC1E",
    x"3ECBC097",
    x"3ECBB50F",
    x"3ECBA988",
    x"3ECB9E00",
    x"3ECB9279",
    x"3ECB86F1",
    x"3ECB7B69",
    x"3ECB6FE1",
    x"3ECB6459",
    x"3ECB58D0",
    x"3ECB4D48",
    x"3ECB41BF",
    x"3ECB3637",
    x"3ECB2AAE",
    x"3ECB1F25",
    x"3ECB139C",
    x"3ECB0813",
    x"3ECAFC89",
    x"3ECAF100",
    x"3ECAE576",
    x"3ECAD9ED",
    x"3ECACE63",
    x"3ECAC2D9",
    x"3ECAB74F",
    x"3ECAABC5",
    x"3ECAA03A",
    x"3ECA94B0",
    x"3ECA8925",
    x"3ECA7D9B",
    x"3ECA7210",
    x"3ECA6685",
    x"3ECA5AFA",
    x"3ECA4F6F",
    x"3ECA43E4",
    x"3ECA3858",
    x"3ECA2CCD",
    x"3ECA2141",
    x"3ECA15B5",
    x"3ECA0A2A",
    x"3EC9FE9E",
    x"3EC9F312",
    x"3EC9E785",
    x"3EC9DBF9",
    x"3EC9D06C",
    x"3EC9C4E0",
    x"3EC9B953",
    x"3EC9ADC6",
    x"3EC9A239",
    x"3EC996AC",
    x"3EC98B1F",
    x"3EC97F92",
    x"3EC97404",
    x"3EC96877",
    x"3EC95CE9",
    x"3EC9515B",
    x"3EC945CD",
    x"3EC93A3F",
    x"3EC92EB1",
    x"3EC92323",
    x"3EC91794",
    x"3EC90C06",
    x"3EC90077",
    x"3EC8F4E8",
    x"3EC8E959",
    x"3EC8DDCA",
    x"3EC8D23B",
    x"3EC8C6AC",
    x"3EC8BB1D",
    x"3EC8AF8D",
    x"3EC8A3FD",
    x"3EC8986E",
    x"3EC88CDE",
    x"3EC8814E",
    x"3EC875BE",
    x"3EC86A2D",
    x"3EC85E9D",
    x"3EC8530D",
    x"3EC8477C",
    x"3EC83BEB",
    x"3EC8305B",
    x"3EC824CA",
    x"3EC81938",
    x"3EC80DA7",
    x"3EC80216",
    x"3EC7F685",
    x"3EC7EAF3",
    x"3EC7DF61",
    x"3EC7D3CF",
    x"3EC7C83E",
    x"3EC7BCAC",
    x"3EC7B119",
    x"3EC7A587",
    x"3EC799F5",
    x"3EC78E62",
    x"3EC782D0",
    x"3EC7773D",
    x"3EC76BAA",
    x"3EC76017",
    x"3EC75484",
    x"3EC748F0",
    x"3EC73D5D",
    x"3EC731CA",
    x"3EC72636",
    x"3EC71AA2",
    x"3EC70F0E",
    x"3EC7037B",
    x"3EC6F7E6",
    x"3EC6EC52",
    x"3EC6E0BE",
    x"3EC6D529",
    x"3EC6C995",
    x"3EC6BE00",
    x"3EC6B26B",
    x"3EC6A6D6",
    x"3EC69B41",
    x"3EC68FAC",
    x"3EC68417",
    x"3EC67882",
    x"3EC66CEC",
    x"3EC66156",
    x"3EC655C1",
    x"3EC64A2B",
    x"3EC63E95",
    x"3EC632FF",
    x"3EC62768",
    x"3EC61BD2",
    x"3EC6103C",
    x"3EC604A5",
    x"3EC5F90E",
    x"3EC5ED77",
    x"3EC5E1E1",
    x"3EC5D649",
    x"3EC5CAB2",
    x"3EC5BF1B",
    x"3EC5B384",
    x"3EC5A7EC",
    x"3EC59C54",
    x"3EC590BD",
    x"3EC58525",
    x"3EC5798D",
    x"3EC56DF4",
    x"3EC5625C",
    x"3EC556C4",
    x"3EC54B2B",
    x"3EC53F93",
    x"3EC533FA",
    x"3EC52861",
    x"3EC51CC8",
    x"3EC5112F",
    x"3EC50596",
    x"3EC4F9FD",
    x"3EC4EE63",
    x"3EC4E2C9",
    x"3EC4D730",
    x"3EC4CB96",
    x"3EC4BFFC",
    x"3EC4B462",
    x"3EC4A8C8",
    x"3EC49D2E",
    x"3EC49193",
    x"3EC485F9",
    x"3EC47A5E",
    x"3EC46EC3",
    x"3EC46328",
    x"3EC4578D",
    x"3EC44BF2",
    x"3EC44057",
    x"3EC434BC",
    x"3EC42920",
    x"3EC41D85",
    x"3EC411E9",
    x"3EC4064D",
    x"3EC3FAB1",
    x"3EC3EF15",
    x"3EC3E379",
    x"3EC3D7DD",
    x"3EC3CC40",
    x"3EC3C0A4",
    x"3EC3B507",
    x"3EC3A96A",
    x"3EC39DCE",
    x"3EC39231",
    x"3EC38693",
    x"3EC37AF6",
    x"3EC36F59",
    x"3EC363BB",
    x"3EC3581E",
    x"3EC34C80",
    x"3EC340E2",
    x"3EC33544",
    x"3EC329A6",
    x"3EC31E08",
    x"3EC3126A",
    x"3EC306CB",
    x"3EC2FB2D",
    x"3EC2EF8E",
    x"3EC2E3EF",
    x"3EC2D851",
    x"3EC2CCB2",
    x"3EC2C112",
    x"3EC2B573",
    x"3EC2A9D4",
    x"3EC29E34",
    x"3EC29295",
    x"3EC286F5",
    x"3EC27B55",
    x"3EC26FB5",
    x"3EC26415",
    x"3EC25875",
    x"3EC24CD5",
    x"3EC24135",
    x"3EC23594",
    x"3EC229F3",
    x"3EC21E53",
    x"3EC212B2",
    x"3EC20711",
    x"3EC1FB70",
    x"3EC1EFCE",
    x"3EC1E42D",
    x"3EC1D88C",
    x"3EC1CCEA",
    x"3EC1C148",
    x"3EC1B5A7",
    x"3EC1AA05",
    x"3EC19E63",
    x"3EC192C0",
    x"3EC1871E",
    x"3EC17B7C",
    x"3EC16FD9",
    x"3EC16437",
    x"3EC15894",
    x"3EC14CF1",
    x"3EC1414E",
    x"3EC135AB",
    x"3EC12A08",
    x"3EC11E64",
    x"3EC112C1",
    x"3EC1071E",
    x"3EC0FB7A",
    x"3EC0EFD6",
    x"3EC0E432",
    x"3EC0D88E",
    x"3EC0CCEA",
    x"3EC0C146",
    x"3EC0B5A1",
    x"3EC0A9FD",
    x"3EC09E58",
    x"3EC092B4",
    x"3EC0870F",
    x"3EC07B6A",
    x"3EC06FC5",
    x"3EC06420",
    x"3EC0587A",
    x"3EC04CD5",
    x"3EC0412F",
    x"3EC0358A",
    x"3EC029E4",
    x"3EC01E3E",
    x"3EC01298",
    x"3EC006F2",
    x"3EBFFB4C",
    x"3EBFEFA5",
    x"3EBFE3FF",
    x"3EBFD858",
    x"3EBFCCB2",
    x"3EBFC10B",
    x"3EBFB564",
    x"3EBFA9BD",
    x"3EBF9E16",
    x"3EBF926F",
    x"3EBF86C7",
    x"3EBF7B20",
    x"3EBF6F78",
    x"3EBF63D0",
    x"3EBF5829",
    x"3EBF4C81",
    x"3EBF40D9",
    x"3EBF3530",
    x"3EBF2988",
    x"3EBF1DE0",
    x"3EBF1237",
    x"3EBF068F",
    x"3EBEFAE6",
    x"3EBEEF3D",
    x"3EBEE394",
    x"3EBED7EB",
    x"3EBECC42",
    x"3EBEC098",
    x"3EBEB4EF",
    x"3EBEA945",
    x"3EBE9D9C",
    x"3EBE91F2",
    x"3EBE8648",
    x"3EBE7A9E",
    x"3EBE6EF4",
    x"3EBE6349",
    x"3EBE579F",
    x"3EBE4BF5",
    x"3EBE404A",
    x"3EBE349F",
    x"3EBE28F4",
    x"3EBE1D4A",
    x"3EBE119E",
    x"3EBE05F3",
    x"3EBDFA48",
    x"3EBDEE9D",
    x"3EBDE2F1",
    x"3EBDD746",
    x"3EBDCB9A",
    x"3EBDBFEE",
    x"3EBDB442",
    x"3EBDA896",
    x"3EBD9CEA",
    x"3EBD913D",
    x"3EBD8591",
    x"3EBD79E4",
    x"3EBD6E38",
    x"3EBD628B",
    x"3EBD56DE",
    x"3EBD4B31",
    x"3EBD3F84",
    x"3EBD33D7",
    x"3EBD2829",
    x"3EBD1C7C",
    x"3EBD10CE",
    x"3EBD0521",
    x"3EBCF973",
    x"3EBCEDC5",
    x"3EBCE217",
    x"3EBCD669",
    x"3EBCCABB",
    x"3EBCBF0C",
    x"3EBCB35E",
    x"3EBCA7AF",
    x"3EBC9C00",
    x"3EBC9052",
    x"3EBC84A3",
    x"3EBC78F4",
    x"3EBC6D45",
    x"3EBC6195",
    x"3EBC55E6",
    x"3EBC4A36",
    x"3EBC3E87",
    x"3EBC32D7",
    x"3EBC2727",
    x"3EBC1B77",
    x"3EBC0FC7",
    x"3EBC0417",
    x"3EBBF867",
    x"3EBBECB6",
    x"3EBBE106",
    x"3EBBD555",
    x"3EBBC9A4",
    x"3EBBBDF4",
    x"3EBBB243",
    x"3EBBA692",
    x"3EBB9AE0",
    x"3EBB8F2F",
    x"3EBB837E",
    x"3EBB77CC",
    x"3EBB6C1A",
    x"3EBB6069",
    x"3EBB54B7",
    x"3EBB4905",
    x"3EBB3D53",
    x"3EBB31A0",
    x"3EBB25EE",
    x"3EBB1A3C",
    x"3EBB0E89",
    x"3EBB02D6",
    x"3EBAF724",
    x"3EBAEB71",
    x"3EBADFBE",
    x"3EBAD40B",
    x"3EBAC857",
    x"3EBABCA4",
    x"3EBAB0F1",
    x"3EBAA53D",
    x"3EBA9989",
    x"3EBA8DD6",
    x"3EBA8222",
    x"3EBA766E",
    x"3EBA6ABA",
    x"3EBA5F05",
    x"3EBA5351",
    x"3EBA479D",
    x"3EBA3BE8",
    x"3EBA3033",
    x"3EBA247F",
    x"3EBA18CA",
    x"3EBA0D15",
    x"3EBA015F",
    x"3EB9F5AA",
    x"3EB9E9F5",
    x"3EB9DE3F",
    x"3EB9D28A",
    x"3EB9C6D4",
    x"3EB9BB1E",
    x"3EB9AF68",
    x"3EB9A3B2",
    x"3EB997FC",
    x"3EB98C46",
    x"3EB98090",
    x"3EB974D9",
    x"3EB96923",
    x"3EB95D6C",
    x"3EB951B5",
    x"3EB945FE",
    x"3EB93A47",
    x"3EB92E90",
    x"3EB922D9",
    x"3EB91721",
    x"3EB90B6A",
    x"3EB8FFB2",
    x"3EB8F3FA",
    x"3EB8E843",
    x"3EB8DC8B",
    x"3EB8D0D3",
    x"3EB8C51B",
    x"3EB8B962",
    x"3EB8ADAA",
    x"3EB8A1F1",
    x"3EB89639",
    x"3EB88A80",
    x"3EB87EC7",
    x"3EB8730E",
    x"3EB86755",
    x"3EB85B9C",
    x"3EB84FE3",
    x"3EB8442A",
    x"3EB83870",
    x"3EB82CB6",
    x"3EB820FD",
    x"3EB81543",
    x"3EB80989",
    x"3EB7FDCF",
    x"3EB7F215",
    x"3EB7E65B",
    x"3EB7DAA0",
    x"3EB7CEE6",
    x"3EB7C32B",
    x"3EB7B770",
    x"3EB7ABB6",
    x"3EB79FFB",
    x"3EB79440",
    x"3EB78884",
    x"3EB77CC9",
    x"3EB7710E",
    x"3EB76552",
    x"3EB75997",
    x"3EB74DDB",
    x"3EB7421F",
    x"3EB73663",
    x"3EB72AA7",
    x"3EB71EEB",
    x"3EB7132F",
    x"3EB70773",
    x"3EB6FBB6",
    x"3EB6EFFA",
    x"3EB6E43D",
    x"3EB6D880",
    x"3EB6CCC3",
    x"3EB6C106",
    x"3EB6B549",
    x"3EB6A98C",
    x"3EB69DCE",
    x"3EB69211",
    x"3EB68653",
    x"3EB67A96",
    x"3EB66ED8",
    x"3EB6631A",
    x"3EB6575C",
    x"3EB64B9E",
    x"3EB63FE0",
    x"3EB63421",
    x"3EB62863",
    x"3EB61CA4",
    x"3EB610E6",
    x"3EB60527",
    x"3EB5F968",
    x"3EB5EDA9",
    x"3EB5E1EA",
    x"3EB5D62B",
    x"3EB5CA6B",
    x"3EB5BEAC",
    x"3EB5B2EC",
    x"3EB5A72D",
    x"3EB59B6D",
    x"3EB58FAD",
    x"3EB583ED",
    x"3EB5782D",
    x"3EB56C6D",
    x"3EB560AC",
    x"3EB554EC",
    x"3EB5492B",
    x"3EB53D6B",
    x"3EB531AA",
    x"3EB525E9",
    x"3EB51A28",
    x"3EB50E67",
    x"3EB502A6",
    x"3EB4F6E5",
    x"3EB4EB23",
    x"3EB4DF62",
    x"3EB4D3A0",
    x"3EB4C7DE",
    x"3EB4BC1D",
    x"3EB4B05B",
    x"3EB4A499",
    x"3EB498D6",
    x"3EB48D14",
    x"3EB48152",
    x"3EB4758F",
    x"3EB469CD",
    x"3EB45E0A",
    x"3EB45247",
    x"3EB44684",
    x"3EB43AC1",
    x"3EB42EFE",
    x"3EB4233B",
    x"3EB41777",
    x"3EB40BB4",
    x"3EB3FFF0",
    x"3EB3F42D",
    x"3EB3E869",
    x"3EB3DCA5",
    x"3EB3D0E1",
    x"3EB3C51D",
    x"3EB3B959",
    x"3EB3AD94",
    x"3EB3A1D0",
    x"3EB3960B",
    x"3EB38A47",
    x"3EB37E82",
    x"3EB372BD",
    x"3EB366F8",
    x"3EB35B33",
    x"3EB34F6E",
    x"3EB343A8",
    x"3EB337E3",
    x"3EB32C1D",
    x"3EB32058",
    x"3EB31492",
    x"3EB308CC",
    x"3EB2FD06",
    x"3EB2F140",
    x"3EB2E57A",
    x"3EB2D9B4",
    x"3EB2CDED",
    x"3EB2C227",
    x"3EB2B660",
    x"3EB2AA99",
    x"3EB29ED3",
    x"3EB2930C",
    x"3EB28745",
    x"3EB27B7E",
    x"3EB26FB6",
    x"3EB263EF",
    x"3EB25827",
    x"3EB24C60",
    x"3EB24098",
    x"3EB234D0",
    x"3EB22909",
    x"3EB21D41",
    x"3EB21178",
    x"3EB205B0",
    x"3EB1F9E8",
    x"3EB1EE1F",
    x"3EB1E257",
    x"3EB1D68E",
    x"3EB1CAC5",
    x"3EB1BEFD",
    x"3EB1B334",
    x"3EB1A76B",
    x"3EB19BA1",
    x"3EB18FD8",
    x"3EB1840F",
    x"3EB17845",
    x"3EB16C7C",
    x"3EB160B2",
    x"3EB154E8",
    x"3EB1491E",
    x"3EB13D54",
    x"3EB1318A",
    x"3EB125C0",
    x"3EB119F5",
    x"3EB10E2B",
    x"3EB10260",
    x"3EB0F696",
    x"3EB0EACB",
    x"3EB0DF00",
    x"3EB0D335",
    x"3EB0C76A",
    x"3EB0BB9F",
    x"3EB0AFD3",
    x"3EB0A408",
    x"3EB0983C",
    x"3EB08C71",
    x"3EB080A5",
    x"3EB074D9",
    x"3EB0690D",
    x"3EB05D41",
    x"3EB05175",
    x"3EB045A9",
    x"3EB039DC",
    x"3EB02E10",
    x"3EB02243",
    x"3EB01677",
    x"3EB00AAA",
    x"3EAFFEDD",
    x"3EAFF310",
    x"3EAFE743",
    x"3EAFDB76",
    x"3EAFCFA8",
    x"3EAFC3DB",
    x"3EAFB80D",
    x"3EAFAC40",
    x"3EAFA072",
    x"3EAF94A4",
    x"3EAF88D6",
    x"3EAF7D08",
    x"3EAF713A",
    x"3EAF656B",
    x"3EAF599D",
    x"3EAF4DCF",
    x"3EAF4200",
    x"3EAF3631",
    x"3EAF2A62",
    x"3EAF1E94",
    x"3EAF12C5",
    x"3EAF06F5",
    x"3EAEFB26",
    x"3EAEEF57",
    x"3EAEE387",
    x"3EAED7B8",
    x"3EAECBE8",
    x"3EAEC018",
    x"3EAEB449",
    x"3EAEA879",
    x"3EAE9CA8",
    x"3EAE90D8",
    x"3EAE8508",
    x"3EAE7938",
    x"3EAE6D67",
    x"3EAE6197",
    x"3EAE55C6",
    x"3EAE49F5",
    x"3EAE3E24",
    x"3EAE3253",
    x"3EAE2682",
    x"3EAE1AB1",
    x"3EAE0EDF",
    x"3EAE030E",
    x"3EADF73C",
    x"3EADEB6B",
    x"3EADDF99",
    x"3EADD3C7",
    x"3EADC7F5",
    x"3EADBC23",
    x"3EADB051",
    x"3EADA47F",
    x"3EAD98AC",
    x"3EAD8CDA",
    x"3EAD8107",
    x"3EAD7534",
    x"3EAD6962",
    x"3EAD5D8F",
    x"3EAD51BC",
    x"3EAD45E9",
    x"3EAD3A15",
    x"3EAD2E42",
    x"3EAD226F",
    x"3EAD169B",
    x"3EAD0AC7",
    x"3EACFEF4",
    x"3EACF320",
    x"3EACE74C",
    x"3EACDB78",
    x"3EACCFA4",
    x"3EACC3CF",
    x"3EACB7FB",
    x"3EACAC27",
    x"3EACA052",
    x"3EAC947D",
    x"3EAC88A9",
    x"3EAC7CD4",
    x"3EAC70FF",
    x"3EAC652A",
    x"3EAC5954",
    x"3EAC4D7F",
    x"3EAC41AA",
    x"3EAC35D4",
    x"3EAC29FF",
    x"3EAC1E29",
    x"3EAC1253",
    x"3EAC067D",
    x"3EABFAA7",
    x"3EABEED1",
    x"3EABE2FB",
    x"3EABD724",
    x"3EABCB4E",
    x"3EABBF77",
    x"3EABB3A1",
    x"3EABA7CA",
    x"3EAB9BF3",
    x"3EAB901C",
    x"3EAB8445",
    x"3EAB786E",
    x"3EAB6C97",
    x"3EAB60BF",
    x"3EAB54E8",
    x"3EAB4910",
    x"3EAB3D39",
    x"3EAB3161",
    x"3EAB2589",
    x"3EAB19B1",
    x"3EAB0DD9",
    x"3EAB0201",
    x"3EAAF628",
    x"3EAAEA50",
    x"3EAADE77",
    x"3EAAD29F",
    x"3EAAC6C6",
    x"3EAABAED",
    x"3EAAAF14",
    x"3EAAA33B",
    x"3EAA9762",
    x"3EAA8B89",
    x"3EAA7FB0",
    x"3EAA73D6",
    x"3EAA67FD",
    x"3EAA5C23",
    x"3EAA5049",
    x"3EAA446F",
    x"3EAA3895",
    x"3EAA2CBB",
    x"3EAA20E1",
    x"3EAA1507",
    x"3EAA092D",
    x"3EA9FD52",
    x"3EA9F178",
    x"3EA9E59D",
    x"3EA9D9C2",
    x"3EA9CDE7",
    x"3EA9C20C",
    x"3EA9B631",
    x"3EA9AA56",
    x"3EA99E7B",
    x"3EA992A0",
    x"3EA986C4",
    x"3EA97AE8",
    x"3EA96F0D",
    x"3EA96331",
    x"3EA95755",
    x"3EA94B79",
    x"3EA93F9D",
    x"3EA933C1",
    x"3EA927E5",
    x"3EA91C08",
    x"3EA9102C",
    x"3EA9044F",
    x"3EA8F872",
    x"3EA8EC95",
    x"3EA8E0B9",
    x"3EA8D4DC",
    x"3EA8C8FE",
    x"3EA8BD21",
    x"3EA8B144",
    x"3EA8A567",
    x"3EA89989",
    x"3EA88DAB",
    x"3EA881CE",
    x"3EA875F0",
    x"3EA86A12",
    x"3EA85E34",
    x"3EA85256",
    x"3EA84678",
    x"3EA83A99",
    x"3EA82EBB",
    x"3EA822DC",
    x"3EA816FE",
    x"3EA80B1F",
    x"3EA7FF40",
    x"3EA7F361",
    x"3EA7E782",
    x"3EA7DBA3",
    x"3EA7CFC4",
    x"3EA7C3E4",
    x"3EA7B805",
    x"3EA7AC25",
    x"3EA7A046",
    x"3EA79466",
    x"3EA78886",
    x"3EA77CA6",
    x"3EA770C6",
    x"3EA764E6",
    x"3EA75906",
    x"3EA74D25",
    x"3EA74145",
    x"3EA73564",
    x"3EA72984",
    x"3EA71DA3",
    x"3EA711C2",
    x"3EA705E1",
    x"3EA6FA00",
    x"3EA6EE1F",
    x"3EA6E23E",
    x"3EA6D65C",
    x"3EA6CA7B",
    x"3EA6BE99",
    x"3EA6B2B8",
    x"3EA6A6D6",
    x"3EA69AF4",
    x"3EA68F12",
    x"3EA68330",
    x"3EA6774E",
    x"3EA66B6C",
    x"3EA65F89",
    x"3EA653A7",
    x"3EA647C4",
    x"3EA63BE2",
    x"3EA62FFF",
    x"3EA6241C",
    x"3EA61839",
    x"3EA60C56",
    x"3EA60073",
    x"3EA5F48F",
    x"3EA5E8AC",
    x"3EA5DCC9",
    x"3EA5D0E5",
    x"3EA5C501",
    x"3EA5B91E",
    x"3EA5AD3A",
    x"3EA5A156",
    x"3EA59572",
    x"3EA5898E",
    x"3EA57DA9",
    x"3EA571C5",
    x"3EA565E1",
    x"3EA559FC",
    x"3EA54E17",
    x"3EA54233",
    x"3EA5364E",
    x"3EA52A69",
    x"3EA51E84",
    x"3EA5129F",
    x"3EA506B9",
    x"3EA4FAD4",
    x"3EA4EEEE",
    x"3EA4E309",
    x"3EA4D723",
    x"3EA4CB3E",
    x"3EA4BF58",
    x"3EA4B372",
    x"3EA4A78C",
    x"3EA49BA6",
    x"3EA48FBF",
    x"3EA483D9",
    x"3EA477F2",
    x"3EA46C0C",
    x"3EA46025",
    x"3EA4543F",
    x"3EA44858",
    x"3EA43C71",
    x"3EA4308A",
    x"3EA424A3",
    x"3EA418BB",
    x"3EA40CD4",
    x"3EA400ED",
    x"3EA3F505",
    x"3EA3E91D",
    x"3EA3DD36",
    x"3EA3D14E",
    x"3EA3C566",
    x"3EA3B97E",
    x"3EA3AD96",
    x"3EA3A1AD",
    x"3EA395C5",
    x"3EA389DD",
    x"3EA37DF4",
    x"3EA3720C",
    x"3EA36623",
    x"3EA35A3A",
    x"3EA34E51",
    x"3EA34268",
    x"3EA3367F",
    x"3EA32A96",
    x"3EA31EAD",
    x"3EA312C3",
    x"3EA306DA",
    x"3EA2FAF0",
    x"3EA2EF06",
    x"3EA2E31C",
    x"3EA2D733",
    x"3EA2CB49",
    x"3EA2BF5E",
    x"3EA2B374",
    x"3EA2A78A",
    x"3EA29BA0",
    x"3EA28FB5",
    x"3EA283CB",
    x"3EA277E0",
    x"3EA26BF5",
    x"3EA2600A",
    x"3EA2541F",
    x"3EA24834",
    x"3EA23C49",
    x"3EA2305E",
    x"3EA22472",
    x"3EA21887",
    x"3EA20C9B",
    x"3EA200B0",
    x"3EA1F4C4",
    x"3EA1E8D8",
    x"3EA1DCEC",
    x"3EA1D100",
    x"3EA1C514",
    x"3EA1B928",
    x"3EA1AD3B",
    x"3EA1A14F",
    x"3EA19562",
    x"3EA18976",
    x"3EA17D89",
    x"3EA1719C",
    x"3EA165AF",
    x"3EA159C2",
    x"3EA14DD5",
    x"3EA141E8",
    x"3EA135FB",
    x"3EA12A0D",
    x"3EA11E20",
    x"3EA11232",
    x"3EA10644",
    x"3EA0FA57",
    x"3EA0EE69",
    x"3EA0E27B",
    x"3EA0D68D",
    x"3EA0CA9E",
    x"3EA0BEB0",
    x"3EA0B2C2",
    x"3EA0A6D3",
    x"3EA09AE5",
    x"3EA08EF6",
    x"3EA08307",
    x"3EA07718",
    x"3EA06B29",
    x"3EA05F3A",
    x"3EA0534B",
    x"3EA0475C",
    x"3EA03B6D",
    x"3EA02F7D",
    x"3EA0238E",
    x"3EA0179E",
    x"3EA00BAE",
    x"3E9FFFBE",
    x"3E9FF3CE",
    x"3E9FE7DE",
    x"3E9FDBEE",
    x"3E9FCFFE",
    x"3E9FC40E",
    x"3E9FB81D",
    x"3E9FAC2D",
    x"3E9FA03C",
    x"3E9F944C",
    x"3E9F885B",
    x"3E9F7C6A",
    x"3E9F7079",
    x"3E9F6488",
    x"3E9F5897",
    x"3E9F4CA5",
    x"3E9F40B4",
    x"3E9F34C3",
    x"3E9F28D1",
    x"3E9F1CDF",
    x"3E9F10EE",
    x"3E9F04FC",
    x"3E9EF90A",
    x"3E9EED18",
    x"3E9EE126",
    x"3E9ED533",
    x"3E9EC941",
    x"3E9EBD4F",
    x"3E9EB15C",
    x"3E9EA569",
    x"3E9E9977",
    x"3E9E8D84",
    x"3E9E8191",
    x"3E9E759E",
    x"3E9E69AB",
    x"3E9E5DB8",
    x"3E9E51C4",
    x"3E9E45D1",
    x"3E9E39DE",
    x"3E9E2DEA",
    x"3E9E21F6",
    x"3E9E1603",
    x"3E9E0A0F",
    x"3E9DFE1B",
    x"3E9DF227",
    x"3E9DE633",
    x"3E9DDA3E",
    x"3E9DCE4A",
    x"3E9DC256",
    x"3E9DB661",
    x"3E9DAA6D",
    x"3E9D9E78",
    x"3E9D9283",
    x"3E9D868E",
    x"3E9D7A99",
    x"3E9D6EA4",
    x"3E9D62AF",
    x"3E9D56BA",
    x"3E9D4AC4",
    x"3E9D3ECF",
    x"3E9D32D9",
    x"3E9D26E3",
    x"3E9D1AEE",
    x"3E9D0EF8",
    x"3E9D0302",
    x"3E9CF70C",
    x"3E9CEB16",
    x"3E9CDF20",
    x"3E9CD329",
    x"3E9CC733",
    x"3E9CBB3C",
    x"3E9CAF46",
    x"3E9CA34F",
    x"3E9C9758",
    x"3E9C8B61",
    x"3E9C7F6A",
    x"3E9C7373",
    x"3E9C677C",
    x"3E9C5B85",
    x"3E9C4F8D",
    x"3E9C4396",
    x"3E9C379E",
    x"3E9C2BA7",
    x"3E9C1FAF",
    x"3E9C13B7",
    x"3E9C07BF",
    x"3E9BFBC7",
    x"3E9BEFCF",
    x"3E9BE3D7",
    x"3E9BD7DF",
    x"3E9BCBE6",
    x"3E9BBFEE",
    x"3E9BB3F5",
    x"3E9BA7FD",
    x"3E9B9C04",
    x"3E9B900B",
    x"3E9B8412",
    x"3E9B7819",
    x"3E9B6C20",
    x"3E9B6027",
    x"3E9B542D",
    x"3E9B4834",
    x"3E9B3C3A",
    x"3E9B3041",
    x"3E9B2447",
    x"3E9B184D",
    x"3E9B0C53",
    x"3E9B0059",
    x"3E9AF45F",
    x"3E9AE865",
    x"3E9ADC6B",
    x"3E9AD070",
    x"3E9AC476",
    x"3E9AB87B",
    x"3E9AAC81",
    x"3E9AA086",
    x"3E9A948B",
    x"3E9A8890",
    x"3E9A7C95",
    x"3E9A709A",
    x"3E9A649F",
    x"3E9A58A4",
    x"3E9A4CA8",
    x"3E9A40AD",
    x"3E9A34B1",
    x"3E9A28B6",
    x"3E9A1CBA",
    x"3E9A10BE",
    x"3E9A04C2",
    x"3E99F8C6",
    x"3E99ECCA",
    x"3E99E0CE",
    x"3E99D4D1",
    x"3E99C8D5",
    x"3E99BCD9",
    x"3E99B0DC",
    x"3E99A4DF",
    x"3E9998E3",
    x"3E998CE6",
    x"3E9980E9",
    x"3E9974EC",
    x"3E9968EE",
    x"3E995CF1",
    x"3E9950F4",
    x"3E9944F7",
    x"3E9938F9",
    x"3E992CFB",
    x"3E9920FE",
    x"3E991500",
    x"3E990902",
    x"3E98FD04",
    x"3E98F106",
    x"3E98E508",
    x"3E98D90A",
    x"3E98CD0B",
    x"3E98C10D",
    x"3E98B50E",
    x"3E98A910",
    x"3E989D11",
    x"3E989112",
    x"3E988513",
    x"3E987914",
    x"3E986D15",
    x"3E986116",
    x"3E985517",
    x"3E984917",
    x"3E983D18",
    x"3E983118",
    x"3E982519",
    x"3E981919",
    x"3E980D19",
    x"3E980119",
    x"3E97F519",
    x"3E97E919",
    x"3E97DD19",
    x"3E97D119",
    x"3E97C518",
    x"3E97B918",
    x"3E97AD17",
    x"3E97A117",
    x"3E979516",
    x"3E978915",
    x"3E977D14",
    x"3E977113",
    x"3E976512",
    x"3E975911",
    x"3E974D10",
    x"3E97410E",
    x"3E97350D",
    x"3E97290B",
    x"3E971D0A",
    x"3E971108",
    x"3E970506",
    x"3E96F904",
    x"3E96ED02",
    x"3E96E100",
    x"3E96D4FE",
    x"3E96C8FC",
    x"3E96BCF9",
    x"3E96B0F7",
    x"3E96A4F4",
    x"3E9698F2",
    x"3E968CEF",
    x"3E9680EC",
    x"3E9674E9",
    x"3E9668E6",
    x"3E965CE3",
    x"3E9650E0",
    x"3E9644DD",
    x"3E9638D9",
    x"3E962CD6",
    x"3E9620D2",
    x"3E9614CF",
    x"3E9608CB",
    x"3E95FCC7",
    x"3E95F0C3",
    x"3E95E4BF",
    x"3E95D8BB",
    x"3E95CCB7",
    x"3E95C0B3",
    x"3E95B4AE",
    x"3E95A8AA",
    x"3E959CA6",
    x"3E9590A1",
    x"3E95849C",
    x"3E957897",
    x"3E956C92",
    x"3E95608D",
    x"3E955488",
    x"3E954883",
    x"3E953C7E",
    x"3E953079",
    x"3E952473",
    x"3E95186E",
    x"3E950C68",
    x"3E950062",
    x"3E94F45D",
    x"3E94E857",
    x"3E94DC51",
    x"3E94D04B",
    x"3E94C444",
    x"3E94B83E",
    x"3E94AC38",
    x"3E94A031",
    x"3E94942B",
    x"3E948824",
    x"3E947C1E",
    x"3E947017",
    x"3E946410",
    x"3E945809",
    x"3E944C02",
    x"3E943FFB",
    x"3E9433F4",
    x"3E9427EC",
    x"3E941BE5",
    x"3E940FDD",
    x"3E9403D6",
    x"3E93F7CE",
    x"3E93EBC6",
    x"3E93DFBF",
    x"3E93D3B7",
    x"3E93C7AF",
    x"3E93BBA6",
    x"3E93AF9E",
    x"3E93A396",
    x"3E93978E",
    x"3E938B85",
    x"3E937F7D",
    x"3E937374",
    x"3E93676B",
    x"3E935B62",
    x"3E934F59",
    x"3E934350",
    x"3E933747",
    x"3E932B3E",
    x"3E931F35",
    x"3E93132B",
    x"3E930722",
    x"3E92FB18",
    x"3E92EF0F",
    x"3E92E305",
    x"3E92D6FB",
    x"3E92CAF1",
    x"3E92BEE7",
    x"3E92B2DD",
    x"3E92A6D3",
    x"3E929AC9",
    x"3E928EBF",
    x"3E9282B4",
    x"3E9276AA",
    x"3E926A9F",
    x"3E925E94",
    x"3E92528A",
    x"3E92467F",
    x"3E923A74",
    x"3E922E69",
    x"3E92225E",
    x"3E921652",
    x"3E920A47",
    x"3E91FE3C",
    x"3E91F230",
    x"3E91E625",
    x"3E91DA19",
    x"3E91CE0D",
    x"3E91C201",
    x"3E91B5F5",
    x"3E91A9E9",
    x"3E919DDD",
    x"3E9191D1",
    x"3E9185C5",
    x"3E9179B9",
    x"3E916DAC",
    x"3E9161A0",
    x"3E915593",
    x"3E914986",
    x"3E913D79",
    x"3E91316D",
    x"3E912560",
    x"3E911953",
    x"3E910D45",
    x"3E910138",
    x"3E90F52B",
    x"3E90E91D",
    x"3E90DD10",
    x"3E90D102",
    x"3E90C4F5",
    x"3E90B8E7",
    x"3E90ACD9",
    x"3E90A0CB",
    x"3E9094BD",
    x"3E9088AF",
    x"3E907CA1",
    x"3E907093",
    x"3E906484",
    x"3E905876",
    x"3E904C67",
    x"3E904059",
    x"3E90344A",
    x"3E90283B",
    x"3E901C2C",
    x"3E90101D",
    x"3E90040E",
    x"3E8FF7FF",
    x"3E8FEBF0",
    x"3E8FDFE0",
    x"3E8FD3D1",
    x"3E8FC7C1",
    x"3E8FBBB2",
    x"3E8FAFA2",
    x"3E8FA392",
    x"3E8F9783",
    x"3E8F8B73",
    x"3E8F7F63",
    x"3E8F7353",
    x"3E8F6742",
    x"3E8F5B32",
    x"3E8F4F22",
    x"3E8F4311",
    x"3E8F3701",
    x"3E8F2AF0",
    x"3E8F1EDF",
    x"3E8F12CF",
    x"3E8F06BE",
    x"3E8EFAAD",
    x"3E8EEE9C",
    x"3E8EE28B",
    x"3E8ED679",
    x"3E8ECA68",
    x"3E8EBE57",
    x"3E8EB245",
    x"3E8EA634",
    x"3E8E9A22",
    x"3E8E8E10",
    x"3E8E81FE",
    x"3E8E75ED",
    x"3E8E69DB",
    x"3E8E5DC8",
    x"3E8E51B6",
    x"3E8E45A4",
    x"3E8E3992",
    x"3E8E2D7F",
    x"3E8E216D",
    x"3E8E155A",
    x"3E8E0947",
    x"3E8DFD35",
    x"3E8DF122",
    x"3E8DE50F",
    x"3E8DD8FC",
    x"3E8DCCE9",
    x"3E8DC0D6",
    x"3E8DB4C2",
    x"3E8DA8AF",
    x"3E8D9C9B",
    x"3E8D9088",
    x"3E8D8474",
    x"3E8D7861",
    x"3E8D6C4D",
    x"3E8D6039",
    x"3E8D5425",
    x"3E8D4811",
    x"3E8D3BFD",
    x"3E8D2FE9",
    x"3E8D23D4",
    x"3E8D17C0",
    x"3E8D0BAB",
    x"3E8CFF97",
    x"3E8CF382",
    x"3E8CE76D",
    x"3E8CDB59",
    x"3E8CCF44",
    x"3E8CC32F",
    x"3E8CB71A",
    x"3E8CAB05",
    x"3E8C9EEF",
    x"3E8C92DA",
    x"3E8C86C5",
    x"3E8C7AAF",
    x"3E8C6E9A",
    x"3E8C6284",
    x"3E8C566E",
    x"3E8C4A58",
    x"3E8C3E42",
    x"3E8C322C",
    x"3E8C2616",
    x"3E8C1A00",
    x"3E8C0DEA",
    x"3E8C01D4",
    x"3E8BF5BD",
    x"3E8BE9A7",
    x"3E8BDD90",
    x"3E8BD179",
    x"3E8BC563",
    x"3E8BB94C",
    x"3E8BAD35",
    x"3E8BA11E",
    x"3E8B9507",
    x"3E8B88F0",
    x"3E8B7CD8",
    x"3E8B70C1",
    x"3E8B64AA",
    x"3E8B5892",
    x"3E8B4C7A",
    x"3E8B4063",
    x"3E8B344B",
    x"3E8B2833",
    x"3E8B1C1B",
    x"3E8B1003",
    x"3E8B03EB",
    x"3E8AF7D3",
    x"3E8AEBBB",
    x"3E8ADFA2",
    x"3E8AD38A",
    x"3E8AC771",
    x"3E8ABB59",
    x"3E8AAF40",
    x"3E8AA327",
    x"3E8A970E",
    x"3E8A8AF5",
    x"3E8A7EDC",
    x"3E8A72C3",
    x"3E8A66AA",
    x"3E8A5A91",
    x"3E8A4E78",
    x"3E8A425E",
    x"3E8A3645",
    x"3E8A2A2B",
    x"3E8A1E11",
    x"3E8A11F7",
    x"3E8A05DE",
    x"3E89F9C4",
    x"3E89EDAA",
    x"3E89E190",
    x"3E89D575",
    x"3E89C95B",
    x"3E89BD41",
    x"3E89B126",
    x"3E89A50C",
    x"3E8998F1",
    x"3E898CD7",
    x"3E8980BC",
    x"3E8974A1",
    x"3E896886",
    x"3E895C6B",
    x"3E895050",
    x"3E894435",
    x"3E893819",
    x"3E892BFE",
    x"3E891FE3",
    x"3E8913C7",
    x"3E8907AC",
    x"3E88FB90",
    x"3E88EF74",
    x"3E88E358",
    x"3E88D73C",
    x"3E88CB20",
    x"3E88BF04",
    x"3E88B2E8",
    x"3E88A6CC",
    x"3E889AB0",
    x"3E888E93",
    x"3E888277",
    x"3E88765A",
    x"3E886A3D",
    x"3E885E21",
    x"3E885204",
    x"3E8845E7",
    x"3E8839CA",
    x"3E882DAD",
    x"3E882190",
    x"3E881572",
    x"3E880955",
    x"3E87FD38",
    x"3E87F11A",
    x"3E87E4FD",
    x"3E87D8DF",
    x"3E87CCC1",
    x"3E87C0A3",
    x"3E87B486",
    x"3E87A868",
    x"3E879C49",
    x"3E87902B",
    x"3E87840D",
    x"3E8777EF",
    x"3E876BD0",
    x"3E875FB2",
    x"3E875393",
    x"3E874775",
    x"3E873B56",
    x"3E872F37",
    x"3E872318",
    x"3E8716F9",
    x"3E870ADA",
    x"3E86FEBB",
    x"3E86F29C",
    x"3E86E67D",
    x"3E86DA5D",
    x"3E86CE3E",
    x"3E86C21F",
    x"3E86B5FF",
    x"3E86A9DF",
    x"3E869DBF",
    x"3E8691A0",
    x"3E868580",
    x"3E867960",
    x"3E866D40",
    x"3E86611F",
    x"3E8654FF",
    x"3E8648DF",
    x"3E863CBE",
    x"3E86309E",
    x"3E86247D",
    x"3E86185D",
    x"3E860C3C",
    x"3E86001B",
    x"3E85F3FA",
    x"3E85E7D9",
    x"3E85DBB8",
    x"3E85CF97",
    x"3E85C376",
    x"3E85B755",
    x"3E85AB33",
    x"3E859F12",
    x"3E8592F0",
    x"3E8586CE",
    x"3E857AAD",
    x"3E856E8B",
    x"3E856269",
    x"3E855647",
    x"3E854A25",
    x"3E853E03",
    x"3E8531E1",
    x"3E8525BF",
    x"3E85199C",
    x"3E850D7A",
    x"3E850157",
    x"3E84F535",
    x"3E84E912",
    x"3E84DCEF",
    x"3E84D0CC",
    x"3E84C4AA",
    x"3E84B887",
    x"3E84AC64",
    x"3E84A040",
    x"3E84941D",
    x"3E8487FA",
    x"3E847BD6",
    x"3E846FB3",
    x"3E84638F",
    x"3E84576C",
    x"3E844B48",
    x"3E843F24",
    x"3E843300",
    x"3E8426DD",
    x"3E841AB8",
    x"3E840E94",
    x"3E840270",
    x"3E83F64C",
    x"3E83EA28",
    x"3E83DE03",
    x"3E83D1DF",
    x"3E83C5BA",
    x"3E83B995",
    x"3E83AD71",
    x"3E83A14C",
    x"3E839527",
    x"3E838902",
    x"3E837CDD",
    x"3E8370B8",
    x"3E836493",
    x"3E83586D",
    x"3E834C48",
    x"3E834022",
    x"3E8333FD",
    x"3E8327D7",
    x"3E831BB2",
    x"3E830F8C",
    x"3E830366",
    x"3E82F740",
    x"3E82EB1A",
    x"3E82DEF4",
    x"3E82D2CE",
    x"3E82C6A8",
    x"3E82BA81",
    x"3E82AE5B",
    x"3E82A234",
    x"3E82960E",
    x"3E8289E7",
    x"3E827DC0",
    x"3E82719A",
    x"3E826573",
    x"3E82594C",
    x"3E824D25",
    x"3E8240FE",
    x"3E8234D7",
    x"3E8228AF",
    x"3E821C88",
    x"3E821060",
    x"3E820439",
    x"3E81F811",
    x"3E81EBEA",
    x"3E81DFC2",
    x"3E81D39A",
    x"3E81C772",
    x"3E81BB4A",
    x"3E81AF22",
    x"3E81A2FA",
    x"3E8196D2",
    x"3E818AAA",
    x"3E817E81",
    x"3E817259",
    x"3E816630",
    x"3E815A08",
    x"3E814DDF",
    x"3E8141B6",
    x"3E81358E",
    x"3E812965",
    x"3E811D3C",
    x"3E811113",
    x"3E8104E9",
    x"3E80F8C0",
    x"3E80EC97",
    x"3E80E06E",
    x"3E80D444",
    x"3E80C81B",
    x"3E80BBF1",
    x"3E80AFC7",
    x"3E80A39E",
    x"3E809774",
    x"3E808B4A",
    x"3E807F20",
    x"3E8072F6",
    x"3E8066CC",
    x"3E805AA1",
    x"3E804E77",
    x"3E80424D",
    x"3E803622",
    x"3E8029F8",
    x"3E801DCD",
    x"3E8011A2",
    x"3E800578",
    x"3E7FF29A",
    x"3E7FDA44",
    x"3E7FC1EE",
    x"3E7FA998",
    x"3E7F9141",
    x"3E7F78EB",
    x"3E7F6094",
    x"3E7F483D",
    x"3E7F2FE7",
    x"3E7F178F",
    x"3E7EFF38",
    x"3E7EE6E1",
    x"3E7ECE89",
    x"3E7EB632",
    x"3E7E9DDA",
    x"3E7E8582",
    x"3E7E6D2A",
    x"3E7E54D1",
    x"3E7E3C79",
    x"3E7E2420",
    x"3E7E0BC8",
    x"3E7DF36F",
    x"3E7DDB16",
    x"3E7DC2BC",
    x"3E7DAA63",
    x"3E7D9209",
    x"3E7D79B0",
    x"3E7D6156",
    x"3E7D48FC",
    x"3E7D30A2",
    x"3E7D1848",
    x"3E7CFFED",
    x"3E7CE793",
    x"3E7CCF38",
    x"3E7CB6DD",
    x"3E7C9E82",
    x"3E7C8627",
    x"3E7C6DCB",
    x"3E7C5570",
    x"3E7C3D14",
    x"3E7C24B8",
    x"3E7C0C5C",
    x"3E7BF400",
    x"3E7BDBA4",
    x"3E7BC348",
    x"3E7BAAEB",
    x"3E7B928E",
    x"3E7B7A31",
    x"3E7B61D4",
    x"3E7B4977",
    x"3E7B311A",
    x"3E7B18BC",
    x"3E7B005F",
    x"3E7AE801",
    x"3E7ACFA3",
    x"3E7AB745",
    x"3E7A9EE7",
    x"3E7A8688",
    x"3E7A6E2A",
    x"3E7A55CB",
    x"3E7A3D6C",
    x"3E7A250D",
    x"3E7A0CAE",
    x"3E79F44F",
    x"3E79DBF0",
    x"3E79C390",
    x"3E79AB30",
    x"3E7992D0",
    x"3E797A70",
    x"3E796210",
    x"3E7949B0",
    x"3E79314F",
    x"3E7918EF",
    x"3E79008E",
    x"3E78E82D",
    x"3E78CFCC",
    x"3E78B76B",
    x"3E789F09",
    x"3E7886A8",
    x"3E786E46",
    x"3E7855E4",
    x"3E783D82",
    x"3E782520",
    x"3E780CBE",
    x"3E77F45B",
    x"3E77DBF9",
    x"3E77C396",
    x"3E77AB33",
    x"3E7792D0",
    x"3E777A6D",
    x"3E77620A",
    x"3E7749A6",
    x"3E773142",
    x"3E7718DF",
    x"3E77007B",
    x"3E76E817",
    x"3E76CFB2",
    x"3E76B74E",
    x"3E769EEA",
    x"3E768685",
    x"3E766E20",
    x"3E7655BB",
    x"3E763D56",
    x"3E7624F1",
    x"3E760C8B",
    x"3E75F426",
    x"3E75DBC0",
    x"3E75C35A",
    x"3E75AAF4",
    x"3E75928E",
    x"3E757A28",
    x"3E7561C1",
    x"3E75495B",
    x"3E7530F4",
    x"3E75188D",
    x"3E750026",
    x"3E74E7BF",
    x"3E74CF57",
    x"3E74B6F0",
    x"3E749E88",
    x"3E748621",
    x"3E746DB9",
    x"3E745551",
    x"3E743CE8",
    x"3E742480",
    x"3E740C18",
    x"3E73F3AF",
    x"3E73DB46",
    x"3E73C2DD",
    x"3E73AA74",
    x"3E73920B",
    x"3E7379A1",
    x"3E736138",
    x"3E7348CE",
    x"3E733064",
    x"3E7317FA",
    x"3E72FF90",
    x"3E72E726",
    x"3E72CEBC",
    x"3E72B651",
    x"3E729DE6",
    x"3E72857B",
    x"3E726D10",
    x"3E7254A5",
    x"3E723C3A",
    x"3E7223CE",
    x"3E720B63",
    x"3E71F2F7",
    x"3E71DA8B",
    x"3E71C21F",
    x"3E71A9B3",
    x"3E719147",
    x"3E7178DA",
    x"3E71606E",
    x"3E714801",
    x"3E712F94",
    x"3E711727",
    x"3E70FEBA",
    x"3E70E64C",
    x"3E70CDDF",
    x"3E70B571",
    x"3E709D04",
    x"3E708496",
    x"3E706C28",
    x"3E7053B9",
    x"3E703B4B",
    x"3E7022DD",
    x"3E700A6E",
    x"3E6FF1FF",
    x"3E6FD990",
    x"3E6FC121",
    x"3E6FA8B2",
    x"3E6F9043",
    x"3E6F77D3",
    x"3E6F5F63",
    x"3E6F46F4",
    x"3E6F2E84",
    x"3E6F1614",
    x"3E6EFDA3",
    x"3E6EE533",
    x"3E6ECCC3",
    x"3E6EB452",
    x"3E6E9BE1",
    x"3E6E8370",
    x"3E6E6AFF",
    x"3E6E528E",
    x"3E6E3A1C",
    x"3E6E21AB",
    x"3E6E0939",
    x"3E6DF0C7",
    x"3E6DD856",
    x"3E6DBFE3",
    x"3E6DA771",
    x"3E6D8EFF",
    x"3E6D768C",
    x"3E6D5E1A",
    x"3E6D45A7",
    x"3E6D2D34",
    x"3E6D14C1",
    x"3E6CFC4E",
    x"3E6CE3DA",
    x"3E6CCB67",
    x"3E6CB2F3",
    x"3E6C9A7F",
    x"3E6C820B",
    x"3E6C6997",
    x"3E6C5123",
    x"3E6C38AF",
    x"3E6C203A",
    x"3E6C07C5",
    x"3E6BEF51",
    x"3E6BD6DC",
    x"3E6BBE66",
    x"3E6BA5F1",
    x"3E6B8D7C",
    x"3E6B7506",
    x"3E6B5C91",
    x"3E6B441B",
    x"3E6B2BA5",
    x"3E6B132F",
    x"3E6AFAB9",
    x"3E6AE242",
    x"3E6AC9CC",
    x"3E6AB155",
    x"3E6A98DE",
    x"3E6A8067",
    x"3E6A67F0",
    x"3E6A4F79",
    x"3E6A3702",
    x"3E6A1E8A",
    x"3E6A0613",
    x"3E69ED9B",
    x"3E69D523",
    x"3E69BCAB",
    x"3E69A433",
    x"3E698BBA",
    x"3E697342",
    x"3E695AC9",
    x"3E694251",
    x"3E6929D8",
    x"3E69115F",
    x"3E68F8E5",
    x"3E68E06C",
    x"3E68C7F3",
    x"3E68AF79",
    x"3E6896FF",
    x"3E687E85",
    x"3E68660B",
    x"3E684D91",
    x"3E683517",
    x"3E681C9C",
    x"3E680422",
    x"3E67EBA7",
    x"3E67D32C",
    x"3E67BAB1",
    x"3E67A236",
    x"3E6789BB",
    x"3E67713F",
    x"3E6758C4",
    x"3E674048",
    x"3E6727CC",
    x"3E670F50",
    x"3E66F6D4",
    x"3E66DE58",
    x"3E66C5DC",
    x"3E66AD5F",
    x"3E6694E2",
    x"3E667C66",
    x"3E6663E9",
    x"3E664B6C",
    x"3E6632EE",
    x"3E661A71",
    x"3E6601F3",
    x"3E65E976",
    x"3E65D0F8",
    x"3E65B87A",
    x"3E659FFC",
    x"3E65877E",
    x"3E656F00",
    x"3E655681",
    x"3E653E02",
    x"3E652584",
    x"3E650D05",
    x"3E64F486",
    x"3E64DC07",
    x"3E64C387",
    x"3E64AB08",
    x"3E649288",
    x"3E647A09",
    x"3E646189",
    x"3E644909",
    x"3E643089",
    x"3E641808",
    x"3E63FF88",
    x"3E63E707",
    x"3E63CE87",
    x"3E63B606",
    x"3E639D85",
    x"3E638504",
    x"3E636C83",
    x"3E635401",
    x"3E633B80",
    x"3E6322FE",
    x"3E630A7C",
    x"3E62F1FA",
    x"3E62D978",
    x"3E62C0F6",
    x"3E62A874",
    x"3E628FF1",
    x"3E62776F",
    x"3E625EEC",
    x"3E624669",
    x"3E622DE6",
    x"3E621563",
    x"3E61FCE0",
    x"3E61E45C",
    x"3E61CBD9",
    x"3E61B355",
    x"3E619AD1",
    x"3E61824D",
    x"3E6169C9",
    x"3E615145",
    x"3E6138C1",
    x"3E61203C",
    x"3E6107B8",
    x"3E60EF33",
    x"3E60D6AE",
    x"3E60BE29",
    x"3E60A5A4",
    x"3E608D1E",
    x"3E607499",
    x"3E605C13",
    x"3E60438E",
    x"3E602B08",
    x"3E601282",
    x"3E5FF9FC",
    x"3E5FE175",
    x"3E5FC8EF",
    x"3E5FB068",
    x"3E5F97E2",
    x"3E5F7F5B",
    x"3E5F66D4",
    x"3E5F4E4D",
    x"3E5F35C6",
    x"3E5F1D3E",
    x"3E5F04B7",
    x"3E5EEC2F",
    x"3E5ED3A8",
    x"3E5EBB20",
    x"3E5EA298",
    x"3E5E8A10",
    x"3E5E7187",
    x"3E5E58FF",
    x"3E5E4076",
    x"3E5E27EE",
    x"3E5E0F65",
    x"3E5DF6DC",
    x"3E5DDE53",
    x"3E5DC5CA",
    x"3E5DAD40",
    x"3E5D94B7",
    x"3E5D7C2D",
    x"3E5D63A4",
    x"3E5D4B1A",
    x"3E5D3290",
    x"3E5D1A05",
    x"3E5D017B",
    x"3E5CE8F1",
    x"3E5CD066",
    x"3E5CB7DC",
    x"3E5C9F51",
    x"3E5C86C6",
    x"3E5C6E3B",
    x"3E5C55B0",
    x"3E5C3D24",
    x"3E5C2499",
    x"3E5C0C0D",
    x"3E5BF381",
    x"3E5BDAF6",
    x"3E5BC26A",
    x"3E5BA9DD",
    x"3E5B9151",
    x"3E5B78C5",
    x"3E5B6038",
    x"3E5B47AC",
    x"3E5B2F1F",
    x"3E5B1692",
    x"3E5AFE05",
    x"3E5AE578",
    x"3E5ACCEA",
    x"3E5AB45D",
    x"3E5A9BCF",
    x"3E5A8341",
    x"3E5A6AB4",
    x"3E5A5226",
    x"3E5A3997",
    x"3E5A2109",
    x"3E5A087B",
    x"3E59EFEC",
    x"3E59D75E",
    x"3E59BECF",
    x"3E59A640",
    x"3E598DB1",
    x"3E597522",
    x"3E595C93",
    x"3E594403",
    x"3E592B74",
    x"3E5912E4",
    x"3E58FA54",
    x"3E58E1C4",
    x"3E58C934",
    x"3E58B0A4",
    x"3E589813",
    x"3E587F83",
    x"3E5866F2",
    x"3E584E62",
    x"3E5835D1",
    x"3E581D40",
    x"3E5804AF",
    x"3E57EC1D",
    x"3E57D38C",
    x"3E57BAFB",
    x"3E57A269",
    x"3E5789D7",
    x"3E577145",
    x"3E5758B3",
    x"3E574021",
    x"3E57278F",
    x"3E570EFC",
    x"3E56F66A",
    x"3E56DDD7",
    x"3E56C544",
    x"3E56ACB1",
    x"3E56941E",
    x"3E567B8B",
    x"3E5662F8",
    x"3E564A64",
    x"3E5631D1",
    x"3E56193D",
    x"3E5600A9",
    x"3E55E815",
    x"3E55CF81",
    x"3E55B6ED",
    x"3E559E58",
    x"3E5585C4",
    x"3E556D2F",
    x"3E55549B",
    x"3E553C06",
    x"3E552371",
    x"3E550ADC",
    x"3E54F246",
    x"3E54D9B1",
    x"3E54C11B",
    x"3E54A886",
    x"3E548FF0",
    x"3E54775A",
    x"3E545EC4",
    x"3E54462E",
    x"3E542D98",
    x"3E541501",
    x"3E53FC6B",
    x"3E53E3D4",
    x"3E53CB3D",
    x"3E53B2A6",
    x"3E539A0F",
    x"3E538178",
    x"3E5368E1",
    x"3E535049",
    x"3E5337B2",
    x"3E531F1A",
    x"3E530682",
    x"3E52EDEA",
    x"3E52D552",
    x"3E52BCBA",
    x"3E52A422",
    x"3E528B89",
    x"3E5272F1",
    x"3E525A58",
    x"3E5241BF",
    x"3E522926",
    x"3E52108D",
    x"3E51F7F4",
    x"3E51DF5B",
    x"3E51C6C1",
    x"3E51AE28",
    x"3E51958E",
    x"3E517CF4",
    x"3E51645A",
    x"3E514BC0",
    x"3E513326",
    x"3E511A8B",
    x"3E5101F1",
    x"3E50E956",
    x"3E50D0BC",
    x"3E50B821",
    x"3E509F86",
    x"3E5086EB",
    x"3E506E4F",
    x"3E5055B4",
    x"3E503D19",
    x"3E50247D",
    x"3E500BE1",
    x"3E4FF345",
    x"3E4FDAA9",
    x"3E4FC20D",
    x"3E4FA971",
    x"3E4F90D5",
    x"3E4F7838",
    x"3E4F5F9C",
    x"3E4F46FF",
    x"3E4F2E62",
    x"3E4F15C5",
    x"3E4EFD28",
    x"3E4EE48B",
    x"3E4ECBED",
    x"3E4EB350",
    x"3E4E9AB2",
    x"3E4E8215",
    x"3E4E6977",
    x"3E4E50D9",
    x"3E4E383B",
    x"3E4E1F9C",
    x"3E4E06FE",
    x"3E4DEE60",
    x"3E4DD5C1",
    x"3E4DBD22",
    x"3E4DA483",
    x"3E4D8BE4",
    x"3E4D7345",
    x"3E4D5AA6",
    x"3E4D4207",
    x"3E4D2967",
    x"3E4D10C8",
    x"3E4CF828",
    x"3E4CDF88",
    x"3E4CC6E8",
    x"3E4CAE48",
    x"3E4C95A8",
    x"3E4C7D08",
    x"3E4C6467",
    x"3E4C4BC7",
    x"3E4C3326",
    x"3E4C1A85",
    x"3E4C01E4",
    x"3E4BE943",
    x"3E4BD0A2",
    x"3E4BB801",
    x"3E4B9F5F",
    x"3E4B86BE",
    x"3E4B6E1C",
    x"3E4B557A",
    x"3E4B3CD8",
    x"3E4B2436",
    x"3E4B0B94",
    x"3E4AF2F2",
    x"3E4ADA4F",
    x"3E4AC1AD",
    x"3E4AA90A",
    x"3E4A9067",
    x"3E4A77C4",
    x"3E4A5F21",
    x"3E4A467E",
    x"3E4A2DDB",
    x"3E4A1538",
    x"3E49FC94",
    x"3E49E3F0",
    x"3E49CB4D",
    x"3E49B2A9",
    x"3E499A05",
    x"3E498161",
    x"3E4968BC",
    x"3E495018",
    x"3E493774",
    x"3E491ECF",
    x"3E49062A",
    x"3E48ED85",
    x"3E48D4E0",
    x"3E48BC3B",
    x"3E48A396",
    x"3E488AF1",
    x"3E48724B",
    x"3E4859A6",
    x"3E484100",
    x"3E48285A",
    x"3E480FB4",
    x"3E47F70E",
    x"3E47DE68",
    x"3E47C5C2",
    x"3E47AD1B",
    x"3E479475",
    x"3E477BCE",
    x"3E476328",
    x"3E474A81",
    x"3E4731DA",
    x"3E471932",
    x"3E47008B",
    x"3E46E7E4",
    x"3E46CF3C",
    x"3E46B695",
    x"3E469DED",
    x"3E468545",
    x"3E466C9D",
    x"3E4653F5",
    x"3E463B4D",
    x"3E4622A5",
    x"3E4609FC",
    x"3E45F153",
    x"3E45D8AB",
    x"3E45C002",
    x"3E45A759",
    x"3E458EB0",
    x"3E457607",
    x"3E455D5E",
    x"3E4544B4",
    x"3E452C0B",
    x"3E451361",
    x"3E44FAB7",
    x"3E44E20D",
    x"3E44C963",
    x"3E44B0B9",
    x"3E44980F",
    x"3E447F65",
    x"3E4466BA",
    x"3E444E10",
    x"3E443565",
    x"3E441CBA",
    x"3E44040F",
    x"3E43EB64",
    x"3E43D2B9",
    x"3E43BA0E",
    x"3E43A162",
    x"3E4388B7",
    x"3E43700B",
    x"3E43575F",
    x"3E433EB3",
    x"3E432607",
    x"3E430D5B",
    x"3E42F4AF",
    x"3E42DC03",
    x"3E42C356",
    x"3E42AAAA",
    x"3E4291FD",
    x"3E427950",
    x"3E4260A3",
    x"3E4247F6",
    x"3E422F49",
    x"3E42169B",
    x"3E41FDEE",
    x"3E41E541",
    x"3E41CC93",
    x"3E41B3E5",
    x"3E419B37",
    x"3E418289",
    x"3E4169DB",
    x"3E41512D",
    x"3E41387F",
    x"3E411FD0",
    x"3E410722",
    x"3E40EE73",
    x"3E40D5C4",
    x"3E40BD15",
    x"3E40A466",
    x"3E408BB7",
    x"3E407308",
    x"3E405A58",
    x"3E4041A9",
    x"3E4028F9",
    x"3E401049",
    x"3E3FF79A",
    x"3E3FDEEA",
    x"3E3FC639",
    x"3E3FAD89",
    x"3E3F94D9",
    x"3E3F7C29",
    x"3E3F6378",
    x"3E3F4AC7",
    x"3E3F3217",
    x"3E3F1966",
    x"3E3F00B5",
    x"3E3EE804",
    x"3E3ECF52",
    x"3E3EB6A1",
    x"3E3E9DEF",
    x"3E3E853E",
    x"3E3E6C8C",
    x"3E3E53DA",
    x"3E3E3B28",
    x"3E3E2276",
    x"3E3E09C4",
    x"3E3DF112",
    x"3E3DD860",
    x"3E3DBFAD",
    x"3E3DA6FA",
    x"3E3D8E48",
    x"3E3D7595",
    x"3E3D5CE2",
    x"3E3D442F",
    x"3E3D2B7C",
    x"3E3D12C8",
    x"3E3CFA15",
    x"3E3CE161",
    x"3E3CC8AE",
    x"3E3CAFFA",
    x"3E3C9746",
    x"3E3C7E92",
    x"3E3C65DE",
    x"3E3C4D2A",
    x"3E3C3476",
    x"3E3C1BC1",
    x"3E3C030D",
    x"3E3BEA58",
    x"3E3BD1A3",
    x"3E3BB8EE",
    x"3E3BA039",
    x"3E3B8784",
    x"3E3B6ECF",
    x"3E3B561A",
    x"3E3B3D64",
    x"3E3B24AF",
    x"3E3B0BF9",
    x"3E3AF343",
    x"3E3ADA8D",
    x"3E3AC1D7",
    x"3E3AA921",
    x"3E3A906B",
    x"3E3A77B4",
    x"3E3A5EFE",
    x"3E3A4647",
    x"3E3A2D91",
    x"3E3A14DA",
    x"3E39FC23",
    x"3E39E36C",
    x"3E39CAB5",
    x"3E39B1FE",
    x"3E399946",
    x"3E39808F",
    x"3E3967D7",
    x"3E394F20",
    x"3E393668",
    x"3E391DB0",
    x"3E3904F8",
    x"3E38EC40",
    x"3E38D387",
    x"3E38BACF",
    x"3E38A217",
    x"3E38895E",
    x"3E3870A5",
    x"3E3857EC",
    x"3E383F33",
    x"3E38267A",
    x"3E380DC1",
    x"3E37F508",
    x"3E37DC4F",
    x"3E37C395",
    x"3E37AADC",
    x"3E379222",
    x"3E377968",
    x"3E3760AE",
    x"3E3747F4",
    x"3E372F3A",
    x"3E371680",
    x"3E36FDC5",
    x"3E36E50B",
    x"3E36CC50",
    x"3E36B396",
    x"3E369ADB",
    x"3E368220",
    x"3E366965",
    x"3E3650AA",
    x"3E3637EF",
    x"3E361F33",
    x"3E360678",
    x"3E35EDBC",
    x"3E35D501",
    x"3E35BC45",
    x"3E35A389",
    x"3E358ACD",
    x"3E357211",
    x"3E355954",
    x"3E354098",
    x"3E3527DC",
    x"3E350F1F",
    x"3E34F662",
    x"3E34DDA6",
    x"3E34C4E9",
    x"3E34AC2C",
    x"3E34936F",
    x"3E347AB2",
    x"3E3461F4",
    x"3E344937",
    x"3E343079",
    x"3E3417BC",
    x"3E33FEFE",
    x"3E33E640",
    x"3E33CD82",
    x"3E33B4C4",
    x"3E339C06",
    x"3E338348",
    x"3E336A89",
    x"3E3351CB",
    x"3E33390C",
    x"3E33204D",
    x"3E33078E",
    x"3E32EECF",
    x"3E32D610",
    x"3E32BD51",
    x"3E32A492",
    x"3E328BD3",
    x"3E327313",
    x"3E325A54",
    x"3E324194",
    x"3E3228D4",
    x"3E321014",
    x"3E31F754",
    x"3E31DE94",
    x"3E31C5D4",
    x"3E31AD13",
    x"3E319453",
    x"3E317B92",
    x"3E3162D2",
    x"3E314A11",
    x"3E313150",
    x"3E31188F",
    x"3E30FFCE",
    x"3E30E70D",
    x"3E30CE4C",
    x"3E30B58A",
    x"3E309CC9",
    x"3E308407",
    x"3E306B45",
    x"3E305284",
    x"3E3039C2",
    x"3E302100",
    x"3E30083D",
    x"3E2FEF7B",
    x"3E2FD6B9",
    x"3E2FBDF6",
    x"3E2FA534",
    x"3E2F8C71",
    x"3E2F73AE",
    x"3E2F5AEB",
    x"3E2F4228",
    x"3E2F2965",
    x"3E2F10A2",
    x"3E2EF7DF",
    x"3E2EDF1B",
    x"3E2EC658",
    x"3E2EAD94",
    x"3E2E94D1",
    x"3E2E7C0D",
    x"3E2E6349",
    x"3E2E4A85",
    x"3E2E31C1",
    x"3E2E18FC",
    x"3E2E0038",
    x"3E2DE773",
    x"3E2DCEAF",
    x"3E2DB5EA",
    x"3E2D9D25",
    x"3E2D8461",
    x"3E2D6B9C",
    x"3E2D52D6",
    x"3E2D3A11",
    x"3E2D214C",
    x"3E2D0887",
    x"3E2CEFC1",
    x"3E2CD6FB",
    x"3E2CBE36",
    x"3E2CA570",
    x"3E2C8CAA",
    x"3E2C73E4",
    x"3E2C5B1E",
    x"3E2C4258",
    x"3E2C2991",
    x"3E2C10CB",
    x"3E2BF804",
    x"3E2BDF3E",
    x"3E2BC677",
    x"3E2BADB0",
    x"3E2B94E9",
    x"3E2B7C22",
    x"3E2B635B",
    x"3E2B4A93",
    x"3E2B31CC",
    x"3E2B1905",
    x"3E2B003D",
    x"3E2AE775",
    x"3E2ACEAE",
    x"3E2AB5E6",
    x"3E2A9D1E",
    x"3E2A8456",
    x"3E2A6B8D",
    x"3E2A52C5",
    x"3E2A39FD",
    x"3E2A2134",
    x"3E2A086B",
    x"3E29EFA3",
    x"3E29D6DA",
    x"3E29BE11",
    x"3E29A548",
    x"3E298C7F",
    x"3E2973B6",
    x"3E295AEC",
    x"3E294223",
    x"3E292959",
    x"3E291090",
    x"3E28F7C6",
    x"3E28DEFC",
    x"3E28C632",
    x"3E28AD68",
    x"3E28949E",
    x"3E287BD4",
    x"3E286309",
    x"3E284A3F",
    x"3E283174",
    x"3E2818AA",
    x"3E27FFDF",
    x"3E27E714",
    x"3E27CE49",
    x"3E27B57E",
    x"3E279CB3",
    x"3E2783E8",
    x"3E276B1C",
    x"3E275251",
    x"3E273985",
    x"3E2720BA",
    x"3E2707EE",
    x"3E26EF22",
    x"3E26D656",
    x"3E26BD8A",
    x"3E26A4BE",
    x"3E268BF2",
    x"3E267325",
    x"3E265A59",
    x"3E26418C",
    x"3E2628C0",
    x"3E260FF3",
    x"3E25F726",
    x"3E25DE59",
    x"3E25C58C",
    x"3E25ACBF",
    x"3E2593F2",
    x"3E257B24",
    x"3E256257",
    x"3E254989",
    x"3E2530BC",
    x"3E2517EE",
    x"3E24FF20",
    x"3E24E652",
    x"3E24CD84",
    x"3E24B4B6",
    x"3E249BE7",
    x"3E248319",
    x"3E246A4B",
    x"3E24517C",
    x"3E2438AD",
    x"3E241FDF",
    x"3E240710",
    x"3E23EE41",
    x"3E23D572",
    x"3E23BCA3",
    x"3E23A3D3",
    x"3E238B04",
    x"3E237235",
    x"3E235965",
    x"3E234095",
    x"3E2327C6",
    x"3E230EF6",
    x"3E22F626",
    x"3E22DD56",
    x"3E22C486",
    x"3E22ABB6",
    x"3E2292E5",
    x"3E227A15",
    x"3E226144",
    x"3E224874",
    x"3E222FA3",
    x"3E2216D2",
    x"3E21FE01",
    x"3E21E530",
    x"3E21CC5F",
    x"3E21B38E",
    x"3E219ABD",
    x"3E2181EB",
    x"3E21691A",
    x"3E215048",
    x"3E213776",
    x"3E211EA5",
    x"3E2105D3",
    x"3E20ED01",
    x"3E20D42F",
    x"3E20BB5C",
    x"3E20A28A",
    x"3E2089B8",
    x"3E2070E5",
    x"3E205813",
    x"3E203F40",
    x"3E20266D",
    x"3E200D9A",
    x"3E1FF4C8",
    x"3E1FDBF4",
    x"3E1FC321",
    x"3E1FAA4E",
    x"3E1F917B",
    x"3E1F78A7",
    x"3E1F5FD4",
    x"3E1F4700",
    x"3E1F2E2C",
    x"3E1F1559",
    x"3E1EFC85",
    x"3E1EE3B1",
    x"3E1ECADD",
    x"3E1EB208",
    x"3E1E9934",
    x"3E1E8060",
    x"3E1E678B",
    x"3E1E4EB7",
    x"3E1E35E2",
    x"3E1E1D0D",
    x"3E1E0438",
    x"3E1DEB63",
    x"3E1DD28E",
    x"3E1DB9B9",
    x"3E1DA0E4",
    x"3E1D880F",
    x"3E1D6F39",
    x"3E1D5664",
    x"3E1D3D8E",
    x"3E1D24B8",
    x"3E1D0BE2",
    x"3E1CF30D",
    x"3E1CDA36",
    x"3E1CC160",
    x"3E1CA88A",
    x"3E1C8FB4",
    x"3E1C76DE",
    x"3E1C5E07",
    x"3E1C4530",
    x"3E1C2C5A",
    x"3E1C1383",
    x"3E1BFAAC",
    x"3E1BE1D5",
    x"3E1BC8FE",
    x"3E1BB027",
    x"3E1B9750",
    x"3E1B7E79",
    x"3E1B65A1",
    x"3E1B4CCA",
    x"3E1B33F2",
    x"3E1B1B1A",
    x"3E1B0242",
    x"3E1AE96B",
    x"3E1AD093",
    x"3E1AB7BB",
    x"3E1A9EE2",
    x"3E1A860A",
    x"3E1A6D32",
    x"3E1A5459",
    x"3E1A3B81",
    x"3E1A22A8",
    x"3E1A09CF",
    x"3E19F0F7",
    x"3E19D81E",
    x"3E19BF45",
    x"3E19A66C",
    x"3E198D92",
    x"3E1974B9",
    x"3E195BE0",
    x"3E194306",
    x"3E192A2D",
    x"3E191153",
    x"3E18F879",
    x"3E18DFA0",
    x"3E18C6C6",
    x"3E18ADEC",
    x"3E189511",
    x"3E187C37",
    x"3E18635D",
    x"3E184A83",
    x"3E1831A8",
    x"3E1818CE",
    x"3E17FFF3",
    x"3E17E718",
    x"3E17CE3D",
    x"3E17B562",
    x"3E179C87",
    x"3E1783AC",
    x"3E176AD1",
    x"3E1751F6",
    x"3E17391A",
    x"3E17203F",
    x"3E170763",
    x"3E16EE88",
    x"3E16D5AC",
    x"3E16BCD0",
    x"3E16A3F4",
    x"3E168B18",
    x"3E16723C",
    x"3E165960",
    x"3E164083",
    x"3E1627A7",
    x"3E160ECB",
    x"3E15F5EE",
    x"3E15DD11",
    x"3E15C435",
    x"3E15AB58",
    x"3E15927B",
    x"3E15799E",
    x"3E1560C1",
    x"3E1547E4",
    x"3E152F06",
    x"3E151629",
    x"3E14FD4B",
    x"3E14E46E",
    x"3E14CB90",
    x"3E14B2B2",
    x"3E1499D5",
    x"3E1480F7",
    x"3E146819",
    x"3E144F3B",
    x"3E14365C",
    x"3E141D7E",
    x"3E1404A0",
    x"3E13EBC1",
    x"3E13D2E3",
    x"3E13BA04",
    x"3E13A125",
    x"3E138847",
    x"3E136F68",
    x"3E135689",
    x"3E133DAA",
    x"3E1324CA",
    x"3E130BEB",
    x"3E12F30C",
    x"3E12DA2C",
    x"3E12C14D",
    x"3E12A86D",
    x"3E128F8E",
    x"3E1276AE",
    x"3E125DCE",
    x"3E1244EE",
    x"3E122C0E",
    x"3E12132E",
    x"3E11FA4E",
    x"3E11E16D",
    x"3E11C88D",
    x"3E11AFAC",
    x"3E1196CC",
    x"3E117DEB",
    x"3E11650A",
    x"3E114C2A",
    x"3E113349",
    x"3E111A68",
    x"3E110186",
    x"3E10E8A5",
    x"3E10CFC4",
    x"3E10B6E3",
    x"3E109E01",
    x"3E108520",
    x"3E106C3E",
    x"3E10535C",
    x"3E103A7B",
    x"3E102199",
    x"3E1008B7",
    x"3E0FEFD5",
    x"3E0FD6F2",
    x"3E0FBE10",
    x"3E0FA52E",
    x"3E0F8C4B",
    x"3E0F7369",
    x"3E0F5A86",
    x"3E0F41A4",
    x"3E0F28C1",
    x"3E0F0FDE",
    x"3E0EF6FB",
    x"3E0EDE18",
    x"3E0EC535",
    x"3E0EAC52",
    x"3E0E936F",
    x"3E0E7A8B",
    x"3E0E61A8",
    x"3E0E48C4",
    x"3E0E2FE1",
    x"3E0E16FD",
    x"3E0DFE19",
    x"3E0DE535",
    x"3E0DCC51",
    x"3E0DB36D",
    x"3E0D9A89",
    x"3E0D81A5",
    x"3E0D68C1",
    x"3E0D4FDC",
    x"3E0D36F8",
    x"3E0D1E13",
    x"3E0D052F",
    x"3E0CEC4A",
    x"3E0CD365",
    x"3E0CBA80",
    x"3E0CA19B",
    x"3E0C88B6",
    x"3E0C6FD1",
    x"3E0C56EC",
    x"3E0C3E07",
    x"3E0C2521",
    x"3E0C0C3C",
    x"3E0BF356",
    x"3E0BDA71",
    x"3E0BC18B",
    x"3E0BA8A5",
    x"3E0B8FBF",
    x"3E0B76D9",
    x"3E0B5DF3",
    x"3E0B450D",
    x"3E0B2C27",
    x"3E0B1340",
    x"3E0AFA5A",
    x"3E0AE173",
    x"3E0AC88D",
    x"3E0AAFA6",
    x"3E0A96BF",
    x"3E0A7DD9",
    x"3E0A64F2",
    x"3E0A4C0B",
    x"3E0A3324",
    x"3E0A1A3C",
    x"3E0A0155",
    x"3E09E86E",
    x"3E09CF86",
    x"3E09B69F",
    x"3E099DB7",
    x"3E0984D0",
    x"3E096BE8",
    x"3E095300",
    x"3E093A18",
    x"3E092130",
    x"3E090848",
    x"3E08EF60",
    x"3E08D678",
    x"3E08BD90",
    x"3E08A4A7",
    x"3E088BBF",
    x"3E0872D6",
    x"3E0859ED",
    x"3E084105",
    x"3E08281C",
    x"3E080F33",
    x"3E07F64A",
    x"3E07DD61",
    x"3E07C478",
    x"3E07AB8F",
    x"3E0792A5",
    x"3E0779BC",
    x"3E0760D2",
    x"3E0747E9",
    x"3E072EFF",
    x"3E071616",
    x"3E06FD2C",
    x"3E06E442",
    x"3E06CB58",
    x"3E06B26E",
    x"3E069984",
    x"3E06809A",
    x"3E0667AF",
    x"3E064EC5",
    x"3E0635DB",
    x"3E061CF0",
    x"3E060405",
    x"3E05EB1B",
    x"3E05D230",
    x"3E05B945",
    x"3E05A05A",
    x"3E05876F",
    x"3E056E84",
    x"3E055599",
    x"3E053CAE",
    x"3E0523C2",
    x"3E050AD7",
    x"3E04F1EB",
    x"3E04D900",
    x"3E04C014",
    x"3E04A729",
    x"3E048E3D",
    x"3E047551",
    x"3E045C65",
    x"3E044379",
    x"3E042A8D",
    x"3E0411A0",
    x"3E03F8B4",
    x"3E03DFC8",
    x"3E03C6DB",
    x"3E03ADEF",
    x"3E039502",
    x"3E037C16",
    x"3E036329",
    x"3E034A3C",
    x"3E03314F",
    x"3E031862",
    x"3E02FF75",
    x"3E02E688",
    x"3E02CD9B",
    x"3E02B4AD",
    x"3E029BC0",
    x"3E0282D2",
    x"3E0269E5",
    x"3E0250F7",
    x"3E02380A",
    x"3E021F1C",
    x"3E02062E",
    x"3E01ED40",
    x"3E01D452",
    x"3E01BB64",
    x"3E01A276",
    x"3E018987",
    x"3E017099",
    x"3E0157AB",
    x"3E013EBC",
    x"3E0125CE",
    x"3E010CDF",
    x"3E00F3F0",
    x"3E00DB01",
    x"3E00C213",
    x"3E00A924",
    x"3E009035",
    x"3E007745",
    x"3E005E56",
    x"3E004567",
    x"3E002C78",
    x"3E001388",
    x"3DFFF531",
    x"3DFFC352",
    x"3DFF9173",
    x"3DFF5F94",
    x"3DFF2DB4",
    x"3DFEFBD4",
    x"3DFEC9F4",
    x"3DFE9814",
    x"3DFE6634",
    x"3DFE3454",
    x"3DFE0273",
    x"3DFDD092",
    x"3DFD9EB2",
    x"3DFD6CD1",
    x"3DFD3AEF",
    x"3DFD090E",
    x"3DFCD72D",
    x"3DFCA54B",
    x"3DFC7369",
    x"3DFC4187",
    x"3DFC0FA5",
    x"3DFBDDC3",
    x"3DFBABE1",
    x"3DFB79FE",
    x"3DFB481C",
    x"3DFB1639",
    x"3DFAE456",
    x"3DFAB273",
    x"3DFA808F",
    x"3DFA4EAC",
    x"3DFA1CC8",
    x"3DF9EAE5",
    x"3DF9B901",
    x"3DF9871D",
    x"3DF95539",
    x"3DF92354",
    x"3DF8F170",
    x"3DF8BF8B",
    x"3DF88DA7",
    x"3DF85BC2",
    x"3DF829DD",
    x"3DF7F7F7",
    x"3DF7C612",
    x"3DF7942C",
    x"3DF76247",
    x"3DF73061",
    x"3DF6FE7B",
    x"3DF6CC95",
    x"3DF69AAF",
    x"3DF668C8",
    x"3DF636E2",
    x"3DF604FB",
    x"3DF5D314",
    x"3DF5A12D",
    x"3DF56F46",
    x"3DF53D5F",
    x"3DF50B77",
    x"3DF4D990",
    x"3DF4A7A8",
    x"3DF475C0",
    x"3DF443D8",
    x"3DF411F0",
    x"3DF3E007",
    x"3DF3AE1F",
    x"3DF37C36",
    x"3DF34A4E",
    x"3DF31865",
    x"3DF2E67C",
    x"3DF2B492",
    x"3DF282A9",
    x"3DF250BF",
    x"3DF21ED6",
    x"3DF1ECEC",
    x"3DF1BB02",
    x"3DF18918",
    x"3DF1572E",
    x"3DF12543",
    x"3DF0F359",
    x"3DF0C16E",
    x"3DF08F83",
    x"3DF05D98",
    x"3DF02BAD",
    x"3DEFF9C2",
    x"3DEFC7D7",
    x"3DEF95EB",
    x"3DEF63FF",
    x"3DEF3214",
    x"3DEF0028",
    x"3DEECE3C",
    x"3DEE9C4F",
    x"3DEE6A63",
    x"3DEE3876",
    x"3DEE068A",
    x"3DEDD49D",
    x"3DEDA2B0",
    x"3DED70C3",
    x"3DED3ED5",
    x"3DED0CE8",
    x"3DECDAFB",
    x"3DECA90D",
    x"3DEC771F",
    x"3DEC4531",
    x"3DEC1343",
    x"3DEBE155",
    x"3DEBAF66",
    x"3DEB7D78",
    x"3DEB4B89",
    x"3DEB199A",
    x"3DEAE7AB",
    x"3DEAB5BC",
    x"3DEA83CD",
    x"3DEA51DE",
    x"3DEA1FEE",
    x"3DE9EDFE",
    x"3DE9BC0E",
    x"3DE98A1F",
    x"3DE9582E",
    x"3DE9263E",
    x"3DE8F44E",
    x"3DE8C25D",
    x"3DE8906D",
    x"3DE85E7C",
    x"3DE82C8B",
    x"3DE7FA9A",
    x"3DE7C8A9",
    x"3DE796B7",
    x"3DE764C6",
    x"3DE732D4",
    x"3DE700E2",
    x"3DE6CEF0",
    x"3DE69CFE",
    x"3DE66B0C",
    x"3DE6391A",
    x"3DE60727",
    x"3DE5D535",
    x"3DE5A342",
    x"3DE5714F",
    x"3DE53F5C",
    x"3DE50D69",
    x"3DE4DB76",
    x"3DE4A982",
    x"3DE4778F",
    x"3DE4459B",
    x"3DE413A7",
    x"3DE3E1B3",
    x"3DE3AFBF",
    x"3DE37DCB",
    x"3DE34BD6",
    x"3DE319E2",
    x"3DE2E7ED",
    x"3DE2B5F8",
    x"3DE28403",
    x"3DE2520E",
    x"3DE22019",
    x"3DE1EE24",
    x"3DE1BC2E",
    x"3DE18A39",
    x"3DE15843",
    x"3DE1264D",
    x"3DE0F457",
    x"3DE0C261",
    x"3DE0906A",
    x"3DE05E74",
    x"3DE02C7D",
    x"3DDFFA87",
    x"3DDFC890",
    x"3DDF9699",
    x"3DDF64A2",
    x"3DDF32AB",
    x"3DDF00B3",
    x"3DDECEBC",
    x"3DDE9CC4",
    x"3DDE6ACC",
    x"3DDE38D4",
    x"3DDE06DC",
    x"3DDDD4E4",
    x"3DDDA2EC",
    x"3DDD70F3",
    x"3DDD3EFB",
    x"3DDD0D02",
    x"3DDCDB09",
    x"3DDCA910",
    x"3DDC7717",
    x"3DDC451E",
    x"3DDC1324",
    x"3DDBE12B",
    x"3DDBAF31",
    x"3DDB7D37",
    x"3DDB4B3D",
    x"3DDB1943",
    x"3DDAE749",
    x"3DDAB54F",
    x"3DDA8354",
    x"3DDA515A",
    x"3DDA1F5F",
    x"3DD9ED64",
    x"3DD9BB69",
    x"3DD9896E",
    x"3DD95773",
    x"3DD92578",
    x"3DD8F37C",
    x"3DD8C181",
    x"3DD88F85",
    x"3DD85D89",
    x"3DD82B8D",
    x"3DD7F991",
    x"3DD7C795",
    x"3DD79598",
    x"3DD7639C",
    x"3DD7319F",
    x"3DD6FFA2",
    x"3DD6CDA5",
    x"3DD69BA8",
    x"3DD669AB",
    x"3DD637AE",
    x"3DD605B0",
    x"3DD5D3B3",
    x"3DD5A1B5",
    x"3DD56FB7",
    x"3DD53DB9",
    x"3DD50BBB",
    x"3DD4D9BD",
    x"3DD4A7BE",
    x"3DD475C0",
    x"3DD443C1",
    x"3DD411C3",
    x"3DD3DFC4",
    x"3DD3ADC5",
    x"3DD37BC6",
    x"3DD349C7",
    x"3DD317C7",
    x"3DD2E5C8",
    x"3DD2B3C8",
    x"3DD281C8",
    x"3DD24FC8",
    x"3DD21DC8",
    x"3DD1EBC8",
    x"3DD1B9C8",
    x"3DD187C8",
    x"3DD155C7",
    x"3DD123C7",
    x"3DD0F1C6",
    x"3DD0BFC5",
    x"3DD08DC4",
    x"3DD05BC3",
    x"3DD029C2",
    x"3DCFF7C0",
    x"3DCFC5BF",
    x"3DCF93BD",
    x"3DCF61BB",
    x"3DCF2FB9",
    x"3DCEFDB7",
    x"3DCECBB5",
    x"3DCE99B3",
    x"3DCE67B1",
    x"3DCE35AE",
    x"3DCE03AB",
    x"3DCDD1A9",
    x"3DCD9FA6",
    x"3DCD6DA3",
    x"3DCD3BA0",
    x"3DCD099C",
    x"3DCCD799",
    x"3DCCA596",
    x"3DCC7392",
    x"3DCC418E",
    x"3DCC0F8A",
    x"3DCBDD86",
    x"3DCBAB82",
    x"3DCB797E",
    x"3DCB477A",
    x"3DCB1575",
    x"3DCAE371",
    x"3DCAB16C",
    x"3DCA7F67",
    x"3DCA4D62",
    x"3DCA1B5D",
    x"3DC9E958",
    x"3DC9B752",
    x"3DC9854D",
    x"3DC95347",
    x"3DC92142",
    x"3DC8EF3C",
    x"3DC8BD36",
    x"3DC88B30",
    x"3DC8592A",
    x"3DC82723",
    x"3DC7F51D",
    x"3DC7C316",
    x"3DC79110",
    x"3DC75F09",
    x"3DC72D02",
    x"3DC6FAFB",
    x"3DC6C8F4",
    x"3DC696ED",
    x"3DC664E5",
    x"3DC632DE",
    x"3DC600D6",
    x"3DC5CECE",
    x"3DC59CC6",
    x"3DC56ABE",
    x"3DC538B6",
    x"3DC506AE",
    x"3DC4D4A6",
    x"3DC4A29D",
    x"3DC47095",
    x"3DC43E8C",
    x"3DC40C83",
    x"3DC3DA7A",
    x"3DC3A871",
    x"3DC37668",
    x"3DC3445F",
    x"3DC31255",
    x"3DC2E04C",
    x"3DC2AE42",
    x"3DC27C39",
    x"3DC24A2F",
    x"3DC21825",
    x"3DC1E61B",
    x"3DC1B410",
    x"3DC18206",
    x"3DC14FFC",
    x"3DC11DF1",
    x"3DC0EBE6",
    x"3DC0B9DC",
    x"3DC087D1",
    x"3DC055C6",
    x"3DC023BA",
    x"3DBFF1AF",
    x"3DBFBFA4",
    x"3DBF8D98",
    x"3DBF5B8D",
    x"3DBF2981",
    x"3DBEF775",
    x"3DBEC569",
    x"3DBE935D",
    x"3DBE6151",
    x"3DBE2F45",
    x"3DBDFD38",
    x"3DBDCB2C",
    x"3DBD991F",
    x"3DBD6712",
    x"3DBD3505",
    x"3DBD02F8",
    x"3DBCD0EB",
    x"3DBC9EDE",
    x"3DBC6CD1",
    x"3DBC3AC3",
    x"3DBC08B6",
    x"3DBBD6A8",
    x"3DBBA49A",
    x"3DBB728C",
    x"3DBB407E",
    x"3DBB0E70",
    x"3DBADC62",
    x"3DBAAA54",
    x"3DBA7845",
    x"3DBA4637",
    x"3DBA1428",
    x"3DB9E219",
    x"3DB9B00A",
    x"3DB97DFB",
    x"3DB94BEC",
    x"3DB919DD",
    x"3DB8E7CE",
    x"3DB8B5BE",
    x"3DB883AF",
    x"3DB8519F",
    x"3DB81F8F",
    x"3DB7ED7F",
    x"3DB7BB6F",
    x"3DB7895F",
    x"3DB7574F",
    x"3DB7253E",
    x"3DB6F32E",
    x"3DB6C11D",
    x"3DB68F0D",
    x"3DB65CFC",
    x"3DB62AEB",
    x"3DB5F8DA",
    x"3DB5C6C9",
    x"3DB594B8",
    x"3DB562A6",
    x"3DB53095",
    x"3DB4FE83",
    x"3DB4CC72",
    x"3DB49A60",
    x"3DB4684E",
    x"3DB4363C",
    x"3DB4042A",
    x"3DB3D218",
    x"3DB3A005",
    x"3DB36DF3",
    x"3DB33BE0",
    x"3DB309CE",
    x"3DB2D7BB",
    x"3DB2A5A8",
    x"3DB27395",
    x"3DB24182",
    x"3DB20F6F",
    x"3DB1DD5C",
    x"3DB1AB48",
    x"3DB17935",
    x"3DB14721",
    x"3DB1150D",
    x"3DB0E2FA",
    x"3DB0B0E6",
    x"3DB07ED2",
    x"3DB04CBD",
    x"3DB01AA9",
    x"3DAFE895",
    x"3DAFB680",
    x"3DAF846C",
    x"3DAF5257",
    x"3DAF2042",
    x"3DAEEE2D",
    x"3DAEBC18",
    x"3DAE8A03",
    x"3DAE57EE",
    x"3DAE25D9",
    x"3DADF3C3",
    x"3DADC1AE",
    x"3DAD8F98",
    x"3DAD5D83",
    x"3DAD2B6D",
    x"3DACF957",
    x"3DACC741",
    x"3DAC952B",
    x"3DAC6314",
    x"3DAC30FE",
    x"3DABFEE8",
    x"3DABCCD1",
    x"3DAB9ABA",
    x"3DAB68A4",
    x"3DAB368D",
    x"3DAB0476",
    x"3DAAD25F",
    x"3DAAA048",
    x"3DAA6E30",
    x"3DAA3C19",
    x"3DAA0A01",
    x"3DA9D7EA",
    x"3DA9A5D2",
    x"3DA973BA",
    x"3DA941A2",
    x"3DA90F8A",
    x"3DA8DD72",
    x"3DA8AB5A",
    x"3DA87942",
    x"3DA84729",
    x"3DA81511",
    x"3DA7E2F8",
    x"3DA7B0E0",
    x"3DA77EC7",
    x"3DA74CAE",
    x"3DA71A95",
    x"3DA6E87C",
    x"3DA6B663",
    x"3DA68449",
    x"3DA65230",
    x"3DA62016",
    x"3DA5EDFD",
    x"3DA5BBE3",
    x"3DA589C9",
    x"3DA557AF",
    x"3DA52595",
    x"3DA4F37B",
    x"3DA4C161",
    x"3DA48F47",
    x"3DA45D2C",
    x"3DA42B12",
    x"3DA3F8F7",
    x"3DA3C6DC",
    x"3DA394C2",
    x"3DA362A7",
    x"3DA3308C",
    x"3DA2FE71",
    x"3DA2CC55",
    x"3DA29A3A",
    x"3DA2681F",
    x"3DA23603",
    x"3DA203E8",
    x"3DA1D1CC",
    x"3DA19FB0",
    x"3DA16D94",
    x"3DA13B78",
    x"3DA1095C",
    x"3DA0D740",
    x"3DA0A524",
    x"3DA07308",
    x"3DA040EB",
    x"3DA00ECF",
    x"3D9FDCB2",
    x"3D9FAA95",
    x"3D9F7878",
    x"3D9F465B",
    x"3D9F143E",
    x"3D9EE221",
    x"3D9EB004",
    x"3D9E7DE7",
    x"3D9E4BC9",
    x"3D9E19AC",
    x"3D9DE78E",
    x"3D9DB570",
    x"3D9D8353",
    x"3D9D5135",
    x"3D9D1F17",
    x"3D9CECF9",
    x"3D9CBADA",
    x"3D9C88BC",
    x"3D9C569E",
    x"3D9C247F",
    x"3D9BF261",
    x"3D9BC042",
    x"3D9B8E23",
    x"3D9B5C05",
    x"3D9B29E6",
    x"3D9AF7C7",
    x"3D9AC5A7",
    x"3D9A9388",
    x"3D9A6169",
    x"3D9A2F4A",
    x"3D99FD2A",
    x"3D99CB0A",
    x"3D9998EB",
    x"3D9966CB",
    x"3D9934AB",
    x"3D99028B",
    x"3D98D06B",
    x"3D989E4B",
    x"3D986C2B",
    x"3D983A0A",
    x"3D9807EA",
    x"3D97D5CA",
    x"3D97A3A9",
    x"3D977188",
    x"3D973F67",
    x"3D970D47",
    x"3D96DB26",
    x"3D96A905",
    x"3D9676E3",
    x"3D9644C2",
    x"3D9612A1",
    x"3D95E07F",
    x"3D95AE5E",
    x"3D957C3C",
    x"3D954A1B",
    x"3D9517F9",
    x"3D94E5D7",
    x"3D94B3B5",
    x"3D948193",
    x"3D944F71",
    x"3D941D4F",
    x"3D93EB2C",
    x"3D93B90A",
    x"3D9386E7",
    x"3D9354C5",
    x"3D9322A2",
    x"3D92F07F",
    x"3D92BE5D",
    x"3D928C3A",
    x"3D925A17",
    x"3D9227F4",
    x"3D91F5D0",
    x"3D91C3AD",
    x"3D91918A",
    x"3D915F66",
    x"3D912D43",
    x"3D90FB1F",
    x"3D90C8FB",
    x"3D9096D8",
    x"3D9064B4",
    x"3D903290",
    x"3D90006C",
    x"3D8FCE47",
    x"3D8F9C23",
    x"3D8F69FF",
    x"3D8F37DA",
    x"3D8F05B6",
    x"3D8ED391",
    x"3D8EA16D",
    x"3D8E6F48",
    x"3D8E3D23",
    x"3D8E0AFE",
    x"3D8DD8D9",
    x"3D8DA6B4",
    x"3D8D748F",
    x"3D8D426A",
    x"3D8D1044",
    x"3D8CDE1F",
    x"3D8CABF9",
    x"3D8C79D4",
    x"3D8C47AE",
    x"3D8C1588",
    x"3D8BE362",
    x"3D8BB13C",
    x"3D8B7F16",
    x"3D8B4CF0",
    x"3D8B1ACA",
    x"3D8AE8A4",
    x"3D8AB67D",
    x"3D8A8457",
    x"3D8A5230",
    x"3D8A200A",
    x"3D89EDE3",
    x"3D89BBBC",
    x"3D898995",
    x"3D89576E",
    x"3D892547",
    x"3D88F320",
    x"3D88C0F9",
    x"3D888ED2",
    x"3D885CAA",
    x"3D882A83",
    x"3D87F85B",
    x"3D87C634",
    x"3D87940C",
    x"3D8761E4",
    x"3D872FBC",
    x"3D86FD94",
    x"3D86CB6C",
    x"3D869944",
    x"3D86671C",
    x"3D8634F4",
    x"3D8602CC",
    x"3D85D0A3",
    x"3D859E7B",
    x"3D856C52",
    x"3D853A29",
    x"3D850801",
    x"3D84D5D8",
    x"3D84A3AF",
    x"3D847186",
    x"3D843F5D",
    x"3D840D34",
    x"3D83DB0A",
    x"3D83A8E1",
    x"3D8376B8",
    x"3D83448E",
    x"3D831265",
    x"3D82E03B",
    x"3D82AE11",
    x"3D827BE8",
    x"3D8249BE",
    x"3D821794",
    x"3D81E56A",
    x"3D81B340",
    x"3D818116",
    x"3D814EEB",
    x"3D811CC1",
    x"3D80EA97",
    x"3D80B86C",
    x"3D808642",
    x"3D805417",
    x"3D8021EC",
    x"3D7FDF83",
    x"3D7F7B2D",
    x"3D7F16D7",
    x"3D7EB281",
    x"3D7E4E2B",
    x"3D7DE9D5",
    x"3D7D857E",
    x"3D7D2127",
    x"3D7CBCD1",
    x"3D7C587A",
    x"3D7BF422",
    x"3D7B8FCB",
    x"3D7B2B74",
    x"3D7AC71C",
    x"3D7A62C5",
    x"3D79FE6D",
    x"3D799A15",
    x"3D7935BC",
    x"3D78D164",
    x"3D786D0C",
    x"3D7808B3",
    x"3D77A45A",
    x"3D774001",
    x"3D76DBA8",
    x"3D76774F",
    x"3D7612F6",
    x"3D75AE9C",
    x"3D754A42",
    x"3D74E5E9",
    x"3D74818F",
    x"3D741D35",
    x"3D73B8DA",
    x"3D735480",
    x"3D72F025",
    x"3D728BCB",
    x"3D722770",
    x"3D71C315",
    x"3D715EBA",
    x"3D70FA5E",
    x"3D709603",
    x"3D7031A8",
    x"3D6FCD4C",
    x"3D6F68F0",
    x"3D6F0494",
    x"3D6EA038",
    x"3D6E3BDC",
    x"3D6DD77F",
    x"3D6D7323",
    x"3D6D0EC6",
    x"3D6CAA69",
    x"3D6C460C",
    x"3D6BE1AF",
    x"3D6B7D51",
    x"3D6B18F4",
    x"3D6AB496",
    x"3D6A5039",
    x"3D69EBDB",
    x"3D69877D",
    x"3D69231F",
    x"3D68BEC1",
    x"3D685A62",
    x"3D67F604",
    x"3D6791A5",
    x"3D672D46",
    x"3D66C8E7",
    x"3D666488",
    x"3D660029",
    x"3D659BC9",
    x"3D65376A",
    x"3D64D30A",
    x"3D646EAA",
    x"3D640A4A",
    x"3D63A5EA",
    x"3D63418A",
    x"3D62DD2A",
    x"3D6278C9",
    x"3D621469",
    x"3D61B008",
    x"3D614BA7",
    x"3D60E746",
    x"3D6082E5",
    x"3D601E83",
    x"3D5FBA22",
    x"3D5F55C0",
    x"3D5EF15F",
    x"3D5E8CFD",
    x"3D5E289B",
    x"3D5DC439",
    x"3D5D5FD7",
    x"3D5CFB74",
    x"3D5C9712",
    x"3D5C32AF",
    x"3D5BCE4C",
    x"3D5B69E9",
    x"3D5B0586",
    x"3D5AA123",
    x"3D5A3CC0",
    x"3D59D85C",
    x"3D5973F9",
    x"3D590F95",
    x"3D58AB31",
    x"3D5846CD",
    x"3D57E269",
    x"3D577E05",
    x"3D5719A1",
    x"3D56B53C",
    x"3D5650D8",
    x"3D55EC73",
    x"3D55880E",
    x"3D5523A9",
    x"3D54BF44",
    x"3D545ADF",
    x"3D53F679",
    x"3D539214",
    x"3D532DAE",
    x"3D52C948",
    x"3D5264E2",
    x"3D52007C",
    x"3D519C16",
    x"3D5137B0",
    x"3D50D34A",
    x"3D506EE3",
    x"3D500A7C",
    x"3D4FA616",
    x"3D4F41AF",
    x"3D4EDD48",
    x"3D4E78E1",
    x"3D4E1479",
    x"3D4DB012",
    x"3D4D4BAA",
    x"3D4CE743",
    x"3D4C82DB",
    x"3D4C1E73",
    x"3D4BBA0B",
    x"3D4B55A3",
    x"3D4AF13B",
    x"3D4A8CD2",
    x"3D4A286A",
    x"3D49C401",
    x"3D495F98",
    x"3D48FB30",
    x"3D4896C7",
    x"3D48325D",
    x"3D47CDF4",
    x"3D47698B",
    x"3D470521",
    x"3D46A0B8",
    x"3D463C4E",
    x"3D45D7E4",
    x"3D45737A",
    x"3D450F10",
    x"3D44AAA6",
    x"3D44463C",
    x"3D43E1D1",
    x"3D437D67",
    x"3D4318FC",
    x"3D42B491",
    x"3D425026",
    x"3D41EBBB",
    x"3D418750",
    x"3D4122E5",
    x"3D40BE7A",
    x"3D405A0E",
    x"3D3FF5A3",
    x"3D3F9137",
    x"3D3F2CCB",
    x"3D3EC85F",
    x"3D3E63F3",
    x"3D3DFF87",
    x"3D3D9B1B",
    x"3D3D36AE",
    x"3D3CD242",
    x"3D3C6DD5",
    x"3D3C0968",
    x"3D3BA4FC",
    x"3D3B408F",
    x"3D3ADC22",
    x"3D3A77B4",
    x"3D3A1347",
    x"3D39AEDA",
    x"3D394A6C",
    x"3D38E5FE",
    x"3D388191",
    x"3D381D23",
    x"3D37B8B5",
    x"3D375447",
    x"3D36EFD9",
    x"3D368B6A",
    x"3D3626FC",
    x"3D35C28D",
    x"3D355E1F",
    x"3D34F9B0",
    x"3D349541",
    x"3D3430D2",
    x"3D33CC63",
    x"3D3367F4",
    x"3D330385",
    x"3D329F15",
    x"3D323AA6",
    x"3D31D636",
    x"3D3171C6",
    x"3D310D57",
    x"3D30A8E7",
    x"3D304477",
    x"3D2FE007",
    x"3D2F7B96",
    x"3D2F1726",
    x"3D2EB2B6",
    x"3D2E4E45",
    x"3D2DE9D4",
    x"3D2D8564",
    x"3D2D20F3",
    x"3D2CBC82",
    x"3D2C5811",
    x"3D2BF39F",
    x"3D2B8F2E",
    x"3D2B2ABD",
    x"3D2AC64B",
    x"3D2A61DA",
    x"3D29FD68",
    x"3D2998F6",
    x"3D293484",
    x"3D28D012",
    x"3D286BA0",
    x"3D28072E",
    x"3D27A2BC",
    x"3D273E49",
    x"3D26D9D7",
    x"3D267564",
    x"3D2610F1",
    x"3D25AC7E",
    x"3D25480C",
    x"3D24E399",
    x"3D247F25",
    x"3D241AB2",
    x"3D23B63F",
    x"3D2351CB",
    x"3D22ED58",
    x"3D2288E4",
    x"3D222471",
    x"3D21BFFD",
    x"3D215B89",
    x"3D20F715",
    x"3D2092A1",
    x"3D202E2D",
    x"3D1FC9B8",
    x"3D1F6544",
    x"3D1F00D0",
    x"3D1E9C5B",
    x"3D1E37E6",
    x"3D1DD372",
    x"3D1D6EFD",
    x"3D1D0A88",
    x"3D1CA613",
    x"3D1C419D",
    x"3D1BDD28",
    x"3D1B78B3",
    x"3D1B143D",
    x"3D1AAFC8",
    x"3D1A4B52",
    x"3D19E6DD",
    x"3D198267",
    x"3D191DF1",
    x"3D18B97B",
    x"3D185505",
    x"3D17F08F",
    x"3D178C18",
    x"3D1727A2",
    x"3D16C32C",
    x"3D165EB5",
    x"3D15FA3F",
    x"3D1595C8",
    x"3D153151",
    x"3D14CCDA",
    x"3D146863",
    x"3D1403EC",
    x"3D139F75",
    x"3D133AFE",
    x"3D12D686",
    x"3D12720F",
    x"3D120D97",
    x"3D11A920",
    x"3D1144A8",
    x"3D10E030",
    x"3D107BB8",
    x"3D101740",
    x"3D0FB2C8",
    x"3D0F4E50",
    x"3D0EE9D8",
    x"3D0E8560",
    x"3D0E20E7",
    x"3D0DBC6F",
    x"3D0D57F6",
    x"3D0CF37E",
    x"3D0C8F05",
    x"3D0C2A8C",
    x"3D0BC613",
    x"3D0B619A",
    x"3D0AFD21",
    x"3D0A98A8",
    x"3D0A342F",
    x"3D09CFB6",
    x"3D096B3C",
    x"3D0906C3",
    x"3D08A249",
    x"3D083DCF",
    x"3D07D956",
    x"3D0774DC",
    x"3D071062",
    x"3D06ABE8",
    x"3D06476E",
    x"3D05E2F4",
    x"3D057E7A",
    x"3D0519FF",
    x"3D04B585",
    x"3D04510B",
    x"3D03EC90",
    x"3D038815",
    x"3D03239B",
    x"3D02BF20",
    x"3D025AA5",
    x"3D01F62A",
    x"3D0191AF",
    x"3D012D34",
    x"3D00C8B9",
    x"3D00643E",
    x"3CFFFF85",
    x"3CFF368E",
    x"3CFE6D97",
    x"3CFDA4A0",
    x"3CFCDBA9",
    x"3CFC12B1",
    x"3CFB49BA",
    x"3CFA80C2",
    x"3CF9B7CA",
    x"3CF8EED2",
    x"3CF825DA",
    x"3CF75CE2",
    x"3CF693E9",
    x"3CF5CAF0",
    x"3CF501F8",
    x"3CF438FF",
    x"3CF37006",
    x"3CF2A70D",
    x"3CF1DE13",
    x"3CF1151A",
    x"3CF04C20",
    x"3CEF8326",
    x"3CEEBA2C",
    x"3CEDF132",
    x"3CED2838",
    x"3CEC5F3E",
    x"3CEB9643",
    x"3CEACD49",
    x"3CEA044E",
    x"3CE93B53",
    x"3CE87258",
    x"3CE7A95D",
    x"3CE6E061",
    x"3CE61766",
    x"3CE54E6A",
    x"3CE4856E",
    x"3CE3BC73",
    x"3CE2F377",
    x"3CE22A7A",
    x"3CE1617E",
    x"3CE09882",
    x"3CDFCF85",
    x"3CDF0688",
    x"3CDE3D8C",
    x"3CDD748F",
    x"3CDCAB91",
    x"3CDBE294",
    x"3CDB1997",
    x"3CDA5099",
    x"3CD9879C",
    x"3CD8BE9E",
    x"3CD7F5A0",
    x"3CD72CA2",
    x"3CD663A4",
    x"3CD59AA6",
    x"3CD4D1A7",
    x"3CD408A9",
    x"3CD33FAA",
    x"3CD276AB",
    x"3CD1ADAC",
    x"3CD0E4AD",
    x"3CD01BAE",
    x"3CCF52AF",
    x"3CCE89AF",
    x"3CCDC0B0",
    x"3CCCF7B0",
    x"3CCC2EB0",
    x"3CCB65B0",
    x"3CCA9CB0",
    x"3CC9D3B0",
    x"3CC90AB0",
    x"3CC841AF",
    x"3CC778AF",
    x"3CC6AFAE",
    x"3CC5E6AD",
    x"3CC51DAC",
    x"3CC454AB",
    x"3CC38BAA",
    x"3CC2C2A9",
    x"3CC1F9A8",
    x"3CC130A6",
    x"3CC067A5",
    x"3CBF9EA3",
    x"3CBED5A1",
    x"3CBE0C9F",
    x"3CBD439D",
    x"3CBC7A9B",
    x"3CBBB199",
    x"3CBAE896",
    x"3CBA1F94",
    x"3CB95691",
    x"3CB88D8E",
    x"3CB7C48C",
    x"3CB6FB89",
    x"3CB63286",
    x"3CB56982",
    x"3CB4A07F",
    x"3CB3D77C",
    x"3CB30E78",
    x"3CB24575",
    x"3CB17C71",
    x"3CB0B36D",
    x"3CAFEA69",
    x"3CAF2165",
    x"3CAE5861",
    x"3CAD8F5D",
    x"3CACC658",
    x"3CABFD54",
    x"3CAB344F",
    x"3CAA6B4B",
    x"3CA9A246",
    x"3CA8D941",
    x"3CA8103C",
    x"3CA74737",
    x"3CA67E32",
    x"3CA5B52C",
    x"3CA4EC27",
    x"3CA42322",
    x"3CA35A1C",
    x"3CA29116",
    x"3CA1C811",
    x"3CA0FF0B",
    x"3CA03605",
    x"3C9F6CFF",
    x"3C9EA3F9",
    x"3C9DDAF2",
    x"3C9D11EC",
    x"3C9C48E6",
    x"3C9B7FDF",
    x"3C9AB6D8",
    x"3C99EDD2",
    x"3C9924CB",
    x"3C985BC4",
    x"3C9792BD",
    x"3C96C9B6",
    x"3C9600AF",
    x"3C9537A7",
    x"3C946EA0",
    x"3C93A599",
    x"3C92DC91",
    x"3C921389",
    x"3C914A82",
    x"3C90817A",
    x"3C8FB872",
    x"3C8EEF6A",
    x"3C8E2662",
    x"3C8D5D5A",
    x"3C8C9452",
    x"3C8BCB49",
    x"3C8B0241",
    x"3C8A3938",
    x"3C897030",
    x"3C88A727",
    x"3C87DE1E",
    x"3C871516",
    x"3C864C0D",
    x"3C858304",
    x"3C84B9FB",
    x"3C83F0F2",
    x"3C8327E8",
    x"3C825EDF",
    x"3C8195D6",
    x"3C80CCCC",
    x"3C8003C3",
    x"3C7E7572",
    x"3C7CE35F",
    x"3C7B514B",
    x"3C79BF38",
    x"3C782D24",
    x"3C769B10",
    x"3C7508FC",
    x"3C7376E7",
    x"3C71E4D3",
    x"3C7052BF",
    x"3C6EC0AA",
    x"3C6D2E95",
    x"3C6B9C80",
    x"3C6A0A6B",
    x"3C687856",
    x"3C66E640",
    x"3C65542B",
    x"3C63C215",
    x"3C622FFF",
    x"3C609DE9",
    x"3C5F0BD3",
    x"3C5D79BD",
    x"3C5BE7A6",
    x"3C5A5590",
    x"3C58C379",
    x"3C573162",
    x"3C559F4C",
    x"3C540D35",
    x"3C527B1D",
    x"3C50E906",
    x"3C4F56EF",
    x"3C4DC4D7",
    x"3C4C32C0",
    x"3C4AA0A8",
    x"3C490E90",
    x"3C477C78",
    x"3C45EA60",
    x"3C445847",
    x"3C42C62F",
    x"3C413417",
    x"3C3FA1FE",
    x"3C3E0FE5",
    x"3C3C7DCC",
    x"3C3AEBB4",
    x"3C39599A",
    x"3C37C781",
    x"3C363568",
    x"3C34A34F",
    x"3C331135",
    x"3C317F1B",
    x"3C2FED02",
    x"3C2E5AE8",
    x"3C2CC8CE",
    x"3C2B36B4",
    x"3C29A49A",
    x"3C281280",
    x"3C268065",
    x"3C24EE4B",
    x"3C235C30",
    x"3C21CA16",
    x"3C2037FB",
    x"3C1EA5E0",
    x"3C1D13C5",
    x"3C1B81AA",
    x"3C19EF8F",
    x"3C185D74",
    x"3C16CB58",
    x"3C15393D",
    x"3C13A722",
    x"3C121506",
    x"3C1082EA",
    x"3C0EF0CF",
    x"3C0D5EB3",
    x"3C0BCC97",
    x"3C0A3A7B",
    x"3C08A85F",
    x"3C071643",
    x"3C058426",
    x"3C03F20A",
    x"3C025FEE",
    x"3C00CDD1",
    x"3BFE7769",
    x"3BFB5330",
    x"3BF82EF6",
    x"3BF50ABD",
    x"3BF1E683",
    x"3BEEC249",
    x"3BEB9E0F",
    x"3BE879D5",
    x"3BE5559B",
    x"3BE23160",
    x"3BDF0D26",
    x"3BDBE8EB",
    x"3BD8C4B0",
    x"3BD5A075",
    x"3BD27C3A",
    x"3BCF57FF",
    x"3BCC33C3",
    x"3BC90F88",
    x"3BC5EB4C",
    x"3BC2C711",
    x"3BBFA2D5",
    x"3BBC7E99",
    x"3BB95A5D",
    x"3BB63621",
    x"3BB311E4",
    x"3BAFEDA8",
    x"3BACC96B",
    x"3BA9A52F",
    x"3BA680F2",
    x"3BA35CB5",
    x"3BA03878",
    x"3B9D143B",
    x"3B99EFFE",
    x"3B96CBC1",
    x"3B93A784",
    x"3B908346",
    x"3B8D5F09",
    x"3B8A3ACB",
    x"3B87168E",
    x"3B83F250",
    x"3B80CE12",
    x"3B7B53A9",
    x"3B750B2D",
    x"3B6EC2B1",
    x"3B687A35",
    x"3B6231B9",
    x"3B5BE93C",
    x"3B55A0C0",
    x"3B4F5843",
    x"3B490FC6",
    x"3B42C749",
    x"3B3C7ECC",
    x"3B36364F",
    x"3B2FEDD1",
    x"3B29A554",
    x"3B235CD7",
    x"3B1D1459",
    x"3B16CBDB",
    x"3B10835D",
    x"3B0A3AE0",
    x"3B03F262",
    x"3AFB53C7",
    x"3AEEC2CB",
    x"3AE231CF",
    x"3AD5A0D2",
    x"3AC90FD5",
    x"3ABC7ED9",
    x"3AAFEDDC",
    x"3AA35CDF",
    x"3A96CBE2",
    x"3A8A3AE5",
    x"3A7B53CF",
    x"3A6231D4",
    x"3A490FD9",
    x"3A2FEDDE",
    x"3A16CBE3",
    x"39FB53D1",
    x"39C90FDA",
    x"3996CBE4",
    x"39490FDB",
    x"38C90FDB",
    x"250D3132",
    x"B8C90FDB",
    x"B9490FDB",
    x"B996CBE4",
    x"B9C90FDA",
    x"B9FB53D1",
    x"BA16CBE3",
    x"BA2FEDDE",
    x"BA490FD9",
    x"BA6231D4",
    x"BA7B53CF",
    x"BA8A3AE5",
    x"BA96CBE2",
    x"BAA35CDF",
    x"BAAFEDDC",
    x"BABC7ED9",
    x"BAC90FD5",
    x"BAD5A0D2",
    x"BAE231CF",
    x"BAEEC2CB",
    x"BAFB53C7",
    x"BB03F262",
    x"BB0A3AE0",
    x"BB10835D",
    x"BB16CBDB",
    x"BB1D1459",
    x"BB235CD7",
    x"BB29A554",
    x"BB2FEDD1",
    x"BB36364F",
    x"BB3C7ECC",
    x"BB42C749",
    x"BB490FC6",
    x"BB4F5843",
    x"BB55A0C0",
    x"BB5BE93C",
    x"BB6231B9",
    x"BB687A35",
    x"BB6EC2B1",
    x"BB750B2D",
    x"BB7B53A9",
    x"BB80CE12",
    x"BB83F250",
    x"BB87168E",
    x"BB8A3ACB",
    x"BB8D5F09",
    x"BB908346",
    x"BB93A784",
    x"BB96CBC1",
    x"BB99EFFE",
    x"BB9D143B",
    x"BBA03878",
    x"BBA35CB5",
    x"BBA680F2",
    x"BBA9A52F",
    x"BBACC96B",
    x"BBAFEDA8",
    x"BBB311E4",
    x"BBB63621",
    x"BBB95A5D",
    x"BBBC7E99",
    x"BBBFA2D5",
    x"BBC2C711",
    x"BBC5EB4C",
    x"BBC90F88",
    x"BBCC33C3",
    x"BBCF57FF",
    x"BBD27C3A",
    x"BBD5A075",
    x"BBD8C4B0",
    x"BBDBE8EB",
    x"BBDF0D26",
    x"BBE23160",
    x"BBE5559B",
    x"BBE879D5",
    x"BBEB9E0F",
    x"BBEEC249",
    x"BBF1E683",
    x"BBF50ABD",
    x"BBF82EF6",
    x"BBFB5330",
    x"BBFE7769",
    x"BC00CDD1",
    x"BC025FEE",
    x"BC03F20A",
    x"BC058426",
    x"BC071643",
    x"BC08A85F",
    x"BC0A3A7B",
    x"BC0BCC97",
    x"BC0D5EB3",
    x"BC0EF0CF",
    x"BC1082EA",
    x"BC121506",
    x"BC13A722",
    x"BC15393D",
    x"BC16CB58",
    x"BC185D74",
    x"BC19EF8F",
    x"BC1B81AA",
    x"BC1D13C5",
    x"BC1EA5E0",
    x"BC2037FB",
    x"BC21CA16",
    x"BC235C30",
    x"BC24EE4B",
    x"BC268065",
    x"BC281280",
    x"BC29A49A",
    x"BC2B36B4",
    x"BC2CC8CE",
    x"BC2E5AE8",
    x"BC2FED02",
    x"BC317F1B",
    x"BC331135",
    x"BC34A34F",
    x"BC363568",
    x"BC37C781",
    x"BC39599A",
    x"BC3AEBB4",
    x"BC3C7DCC",
    x"BC3E0FE5",
    x"BC3FA1FE",
    x"BC413417",
    x"BC42C62F",
    x"BC445847",
    x"BC45EA60",
    x"BC477C78",
    x"BC490E90",
    x"BC4AA0A8",
    x"BC4C32C0",
    x"BC4DC4D7",
    x"BC4F56EF",
    x"BC50E906",
    x"BC527B1D",
    x"BC540D35",
    x"BC559F4C",
    x"BC573162",
    x"BC58C379",
    x"BC5A5590",
    x"BC5BE7A6",
    x"BC5D79BD",
    x"BC5F0BD3",
    x"BC609DE9",
    x"BC622FFF",
    x"BC63C215",
    x"BC65542B",
    x"BC66E640",
    x"BC687856",
    x"BC6A0A6B",
    x"BC6B9C80",
    x"BC6D2E95",
    x"BC6EC0AA",
    x"BC7052BF",
    x"BC71E4D3",
    x"BC7376E7",
    x"BC7508FC",
    x"BC769B10",
    x"BC782D24",
    x"BC79BF38",
    x"BC7B514B",
    x"BC7CE35F",
    x"BC7E7572",
    x"BC8003C3",
    x"BC80CCCC",
    x"BC8195D6",
    x"BC825EDF",
    x"BC8327E8",
    x"BC83F0F2",
    x"BC84B9FB",
    x"BC858304",
    x"BC864C0D",
    x"BC871516",
    x"BC87DE1E",
    x"BC88A727",
    x"BC897030",
    x"BC8A3938",
    x"BC8B0241",
    x"BC8BCB49",
    x"BC8C9452",
    x"BC8D5D5A",
    x"BC8E2662",
    x"BC8EEF6A",
    x"BC8FB872",
    x"BC90817A",
    x"BC914A82",
    x"BC921389",
    x"BC92DC91",
    x"BC93A599",
    x"BC946EA0",
    x"BC9537A7",
    x"BC9600AF",
    x"BC96C9B6",
    x"BC9792BD",
    x"BC985BC4",
    x"BC9924CB",
    x"BC99EDD2",
    x"BC9AB6D8",
    x"BC9B7FDF",
    x"BC9C48E6",
    x"BC9D11EC",
    x"BC9DDAF2",
    x"BC9EA3F9",
    x"BC9F6CFF",
    x"BCA03605",
    x"BCA0FF0B",
    x"BCA1C811",
    x"BCA29116",
    x"BCA35A1C",
    x"BCA42322",
    x"BCA4EC27",
    x"BCA5B52C",
    x"BCA67E32",
    x"BCA74737",
    x"BCA8103C",
    x"BCA8D941",
    x"BCA9A246",
    x"BCAA6B4B",
    x"BCAB344F",
    x"BCABFD54",
    x"BCACC658",
    x"BCAD8F5D",
    x"BCAE5861",
    x"BCAF2165",
    x"BCAFEA69",
    x"BCB0B36D",
    x"BCB17C71",
    x"BCB24575",
    x"BCB30E78",
    x"BCB3D77C",
    x"BCB4A07F",
    x"BCB56982",
    x"BCB63286",
    x"BCB6FB89",
    x"BCB7C48C",
    x"BCB88D8E",
    x"BCB95691",
    x"BCBA1F94",
    x"BCBAE896",
    x"BCBBB199",
    x"BCBC7A9B",
    x"BCBD439D",
    x"BCBE0C9F",
    x"BCBED5A1",
    x"BCBF9EA3",
    x"BCC067A5",
    x"BCC130A6",
    x"BCC1F9A8",
    x"BCC2C2A9",
    x"BCC38BAA",
    x"BCC454AB",
    x"BCC51DAC",
    x"BCC5E6AD",
    x"BCC6AFAE",
    x"BCC778AF",
    x"BCC841AF",
    x"BCC90AB0",
    x"BCC9D3B0",
    x"BCCA9CB0",
    x"BCCB65B0",
    x"BCCC2EB0",
    x"BCCCF7B0",
    x"BCCDC0B0",
    x"BCCE89AF",
    x"BCCF52AF",
    x"BCD01BAE",
    x"BCD0E4AD",
    x"BCD1ADAC",
    x"BCD276AB",
    x"BCD33FAA",
    x"BCD408A9",
    x"BCD4D1A7",
    x"BCD59AA6",
    x"BCD663A4",
    x"BCD72CA2",
    x"BCD7F5A0",
    x"BCD8BE9E",
    x"BCD9879C",
    x"BCDA5099",
    x"BCDB1997",
    x"BCDBE294",
    x"BCDCAB91",
    x"BCDD748F",
    x"BCDE3D8C",
    x"BCDF0688",
    x"BCDFCF85",
    x"BCE09882",
    x"BCE1617E",
    x"BCE22A7A",
    x"BCE2F377",
    x"BCE3BC73",
    x"BCE4856E",
    x"BCE54E6A",
    x"BCE61766",
    x"BCE6E061",
    x"BCE7A95D",
    x"BCE87258",
    x"BCE93B53",
    x"BCEA044E",
    x"BCEACD49",
    x"BCEB9643",
    x"BCEC5F3E",
    x"BCED2838",
    x"BCEDF132",
    x"BCEEBA2C",
    x"BCEF8326",
    x"BCF04C20",
    x"BCF1151A",
    x"BCF1DE13",
    x"BCF2A70D",
    x"BCF37006",
    x"BCF438FF",
    x"BCF501F8",
    x"BCF5CAF0",
    x"BCF693E9",
    x"BCF75CE2",
    x"BCF825DA",
    x"BCF8EED2",
    x"BCF9B7CA",
    x"BCFA80C2",
    x"BCFB49BA",
    x"BCFC12B1",
    x"BCFCDBA9",
    x"BCFDA4A0",
    x"BCFE6D97",
    x"BCFF368E",
    x"BCFFFF85",
    x"BD00643E",
    x"BD00C8B9",
    x"BD012D34",
    x"BD0191AF",
    x"BD01F62A",
    x"BD025AA5",
    x"BD02BF20",
    x"BD03239B",
    x"BD038815",
    x"BD03EC90",
    x"BD04510B",
    x"BD04B585",
    x"BD0519FF",
    x"BD057E7A",
    x"BD05E2F4",
    x"BD06476E",
    x"BD06ABE8",
    x"BD071062",
    x"BD0774DC",
    x"BD07D956",
    x"BD083DCF",
    x"BD08A249",
    x"BD0906C3",
    x"BD096B3C",
    x"BD09CFB6",
    x"BD0A342F",
    x"BD0A98A8",
    x"BD0AFD21",
    x"BD0B619A",
    x"BD0BC613",
    x"BD0C2A8C",
    x"BD0C8F05",
    x"BD0CF37E",
    x"BD0D57F6",
    x"BD0DBC6F",
    x"BD0E20E7",
    x"BD0E8560",
    x"BD0EE9D8",
    x"BD0F4E50",
    x"BD0FB2C8",
    x"BD101740",
    x"BD107BB8",
    x"BD10E030",
    x"BD1144A8",
    x"BD11A920",
    x"BD120D97",
    x"BD12720F",
    x"BD12D686",
    x"BD133AFE",
    x"BD139F75",
    x"BD1403EC",
    x"BD146863",
    x"BD14CCDA",
    x"BD153151",
    x"BD1595C8",
    x"BD15FA3F",
    x"BD165EB5",
    x"BD16C32C",
    x"BD1727A2",
    x"BD178C18",
    x"BD17F08F",
    x"BD185505",
    x"BD18B97B",
    x"BD191DF1",
    x"BD198267",
    x"BD19E6DD",
    x"BD1A4B52",
    x"BD1AAFC8",
    x"BD1B143D",
    x"BD1B78B3",
    x"BD1BDD28",
    x"BD1C419D",
    x"BD1CA613",
    x"BD1D0A88",
    x"BD1D6EFD",
    x"BD1DD372",
    x"BD1E37E6",
    x"BD1E9C5B",
    x"BD1F00D0",
    x"BD1F6544",
    x"BD1FC9B8",
    x"BD202E2D",
    x"BD2092A1",
    x"BD20F715",
    x"BD215B89",
    x"BD21BFFD",
    x"BD222471",
    x"BD2288E4",
    x"BD22ED58",
    x"BD2351CB",
    x"BD23B63F",
    x"BD241AB2",
    x"BD247F25",
    x"BD24E399",
    x"BD25480C",
    x"BD25AC7E",
    x"BD2610F1",
    x"BD267564",
    x"BD26D9D7",
    x"BD273E49",
    x"BD27A2BC",
    x"BD28072E",
    x"BD286BA0",
    x"BD28D012",
    x"BD293484",
    x"BD2998F6",
    x"BD29FD68",
    x"BD2A61DA",
    x"BD2AC64B",
    x"BD2B2ABD",
    x"BD2B8F2E",
    x"BD2BF39F",
    x"BD2C5811",
    x"BD2CBC82",
    x"BD2D20F3",
    x"BD2D8564",
    x"BD2DE9D4",
    x"BD2E4E45",
    x"BD2EB2B6",
    x"BD2F1726",
    x"BD2F7B96",
    x"BD2FE007",
    x"BD304477",
    x"BD30A8E7",
    x"BD310D57",
    x"BD3171C6",
    x"BD31D636",
    x"BD323AA6",
    x"BD329F15",
    x"BD330385",
    x"BD3367F4",
    x"BD33CC63",
    x"BD3430D2",
    x"BD349541",
    x"BD34F9B0",
    x"BD355E1F",
    x"BD35C28D",
    x"BD3626FC",
    x"BD368B6A",
    x"BD36EFD9",
    x"BD375447",
    x"BD37B8B5",
    x"BD381D23",
    x"BD388191",
    x"BD38E5FE",
    x"BD394A6C",
    x"BD39AEDA",
    x"BD3A1347",
    x"BD3A77B4",
    x"BD3ADC22",
    x"BD3B408F",
    x"BD3BA4FC",
    x"BD3C0968",
    x"BD3C6DD5",
    x"BD3CD242",
    x"BD3D36AE",
    x"BD3D9B1B",
    x"BD3DFF87",
    x"BD3E63F3",
    x"BD3EC85F",
    x"BD3F2CCB",
    x"BD3F9137",
    x"BD3FF5A3",
    x"BD405A0E",
    x"BD40BE7A",
    x"BD4122E5",
    x"BD418750",
    x"BD41EBBB",
    x"BD425026",
    x"BD42B491",
    x"BD4318FC",
    x"BD437D67",
    x"BD43E1D1",
    x"BD44463C",
    x"BD44AAA6",
    x"BD450F10",
    x"BD45737A",
    x"BD45D7E4",
    x"BD463C4E",
    x"BD46A0B8",
    x"BD470521",
    x"BD47698B",
    x"BD47CDF4",
    x"BD48325D",
    x"BD4896C7",
    x"BD48FB30",
    x"BD495F98",
    x"BD49C401",
    x"BD4A286A",
    x"BD4A8CD2",
    x"BD4AF13B",
    x"BD4B55A3",
    x"BD4BBA0B",
    x"BD4C1E73",
    x"BD4C82DB",
    x"BD4CE743",
    x"BD4D4BAA",
    x"BD4DB012",
    x"BD4E1479",
    x"BD4E78E1",
    x"BD4EDD48",
    x"BD4F41AF",
    x"BD4FA616",
    x"BD500A7C",
    x"BD506EE3",
    x"BD50D34A",
    x"BD5137B0",
    x"BD519C16",
    x"BD52007C",
    x"BD5264E2",
    x"BD52C948",
    x"BD532DAE",
    x"BD539214",
    x"BD53F679",
    x"BD545ADF",
    x"BD54BF44",
    x"BD5523A9",
    x"BD55880E",
    x"BD55EC73",
    x"BD5650D8",
    x"BD56B53C",
    x"BD5719A1",
    x"BD577E05",
    x"BD57E269",
    x"BD5846CD",
    x"BD58AB31",
    x"BD590F95",
    x"BD5973F9",
    x"BD59D85C",
    x"BD5A3CC0",
    x"BD5AA123",
    x"BD5B0586",
    x"BD5B69E9",
    x"BD5BCE4C",
    x"BD5C32AF",
    x"BD5C9712",
    x"BD5CFB74",
    x"BD5D5FD7",
    x"BD5DC439",
    x"BD5E289B",
    x"BD5E8CFD",
    x"BD5EF15F",
    x"BD5F55C0",
    x"BD5FBA22",
    x"BD601E83",
    x"BD6082E5",
    x"BD60E746",
    x"BD614BA7",
    x"BD61B008",
    x"BD621469",
    x"BD6278C9",
    x"BD62DD2A",
    x"BD63418A",
    x"BD63A5EA",
    x"BD640A4A",
    x"BD646EAA",
    x"BD64D30A",
    x"BD65376A",
    x"BD659BC9",
    x"BD660029",
    x"BD666488",
    x"BD66C8E7",
    x"BD672D46",
    x"BD6791A5",
    x"BD67F604",
    x"BD685A62",
    x"BD68BEC1",
    x"BD69231F",
    x"BD69877D",
    x"BD69EBDB",
    x"BD6A5039",
    x"BD6AB496",
    x"BD6B18F4",
    x"BD6B7D51",
    x"BD6BE1AF",
    x"BD6C460C",
    x"BD6CAA69",
    x"BD6D0EC6",
    x"BD6D7323",
    x"BD6DD77F",
    x"BD6E3BDC",
    x"BD6EA038",
    x"BD6F0494",
    x"BD6F68F0",
    x"BD6FCD4C",
    x"BD7031A8",
    x"BD709603",
    x"BD70FA5E",
    x"BD715EBA",
    x"BD71C315",
    x"BD722770",
    x"BD728BCB",
    x"BD72F025",
    x"BD735480",
    x"BD73B8DA",
    x"BD741D35",
    x"BD74818F",
    x"BD74E5E9",
    x"BD754A42",
    x"BD75AE9C",
    x"BD7612F6",
    x"BD76774F",
    x"BD76DBA8",
    x"BD774001",
    x"BD77A45A",
    x"BD7808B3",
    x"BD786D0C",
    x"BD78D164",
    x"BD7935BC",
    x"BD799A15",
    x"BD79FE6D",
    x"BD7A62C5",
    x"BD7AC71C",
    x"BD7B2B74",
    x"BD7B8FCB",
    x"BD7BF422",
    x"BD7C587A",
    x"BD7CBCD1",
    x"BD7D2127",
    x"BD7D857E",
    x"BD7DE9D5",
    x"BD7E4E2B",
    x"BD7EB281",
    x"BD7F16D7",
    x"BD7F7B2D",
    x"BD7FDF83",
    x"BD8021EC",
    x"BD805417",
    x"BD808642",
    x"BD80B86C",
    x"BD80EA97",
    x"BD811CC1",
    x"BD814EEB",
    x"BD818116",
    x"BD81B340",
    x"BD81E56A",
    x"BD821794",
    x"BD8249BE",
    x"BD827BE8",
    x"BD82AE11",
    x"BD82E03B",
    x"BD831265",
    x"BD83448E",
    x"BD8376B8",
    x"BD83A8E1",
    x"BD83DB0A",
    x"BD840D34",
    x"BD843F5D",
    x"BD847186",
    x"BD84A3AF",
    x"BD84D5D8",
    x"BD850801",
    x"BD853A29",
    x"BD856C52",
    x"BD859E7B",
    x"BD85D0A3",
    x"BD8602CC",
    x"BD8634F4",
    x"BD86671C",
    x"BD869944",
    x"BD86CB6C",
    x"BD86FD94",
    x"BD872FBC",
    x"BD8761E4",
    x"BD87940C",
    x"BD87C634",
    x"BD87F85B",
    x"BD882A83",
    x"BD885CAA",
    x"BD888ED2",
    x"BD88C0F9",
    x"BD88F320",
    x"BD892547",
    x"BD89576E",
    x"BD898995",
    x"BD89BBBC",
    x"BD89EDE3",
    x"BD8A200A",
    x"BD8A5230",
    x"BD8A8457",
    x"BD8AB67D",
    x"BD8AE8A4",
    x"BD8B1ACA",
    x"BD8B4CF0",
    x"BD8B7F16",
    x"BD8BB13C",
    x"BD8BE362",
    x"BD8C1588",
    x"BD8C47AE",
    x"BD8C79D4",
    x"BD8CABF9",
    x"BD8CDE1F",
    x"BD8D1044",
    x"BD8D426A",
    x"BD8D748F",
    x"BD8DA6B4",
    x"BD8DD8D9",
    x"BD8E0AFE",
    x"BD8E3D23",
    x"BD8E6F48",
    x"BD8EA16D",
    x"BD8ED391",
    x"BD8F05B6",
    x"BD8F37DA",
    x"BD8F69FF",
    x"BD8F9C23",
    x"BD8FCE47",
    x"BD90006C",
    x"BD903290",
    x"BD9064B4",
    x"BD9096D8",
    x"BD90C8FB",
    x"BD90FB1F",
    x"BD912D43",
    x"BD915F66",
    x"BD91918A",
    x"BD91C3AD",
    x"BD91F5D0",
    x"BD9227F4",
    x"BD925A17",
    x"BD928C3A",
    x"BD92BE5D",
    x"BD92F07F",
    x"BD9322A2",
    x"BD9354C5",
    x"BD9386E7",
    x"BD93B90A",
    x"BD93EB2C",
    x"BD941D4F",
    x"BD944F71",
    x"BD948193",
    x"BD94B3B5",
    x"BD94E5D7",
    x"BD9517F9",
    x"BD954A1B",
    x"BD957C3C",
    x"BD95AE5E",
    x"BD95E07F",
    x"BD9612A1",
    x"BD9644C2",
    x"BD9676E3",
    x"BD96A905",
    x"BD96DB26",
    x"BD970D47",
    x"BD973F67",
    x"BD977188",
    x"BD97A3A9",
    x"BD97D5CA",
    x"BD9807EA",
    x"BD983A0A",
    x"BD986C2B",
    x"BD989E4B",
    x"BD98D06B",
    x"BD99028B",
    x"BD9934AB",
    x"BD9966CB",
    x"BD9998EB",
    x"BD99CB0A",
    x"BD99FD2A",
    x"BD9A2F4A",
    x"BD9A6169",
    x"BD9A9388",
    x"BD9AC5A7",
    x"BD9AF7C7",
    x"BD9B29E6",
    x"BD9B5C05",
    x"BD9B8E23",
    x"BD9BC042",
    x"BD9BF261",
    x"BD9C247F",
    x"BD9C569E",
    x"BD9C88BC",
    x"BD9CBADA",
    x"BD9CECF9",
    x"BD9D1F17",
    x"BD9D5135",
    x"BD9D8353",
    x"BD9DB570",
    x"BD9DE78E",
    x"BD9E19AC",
    x"BD9E4BC9",
    x"BD9E7DE7",
    x"BD9EB004",
    x"BD9EE221",
    x"BD9F143E",
    x"BD9F465B",
    x"BD9F7878",
    x"BD9FAA95",
    x"BD9FDCB2",
    x"BDA00ECF",
    x"BDA040EB",
    x"BDA07308",
    x"BDA0A524",
    x"BDA0D740",
    x"BDA1095C",
    x"BDA13B78",
    x"BDA16D94",
    x"BDA19FB0",
    x"BDA1D1CC",
    x"BDA203E8",
    x"BDA23603",
    x"BDA2681F",
    x"BDA29A3A",
    x"BDA2CC55",
    x"BDA2FE71",
    x"BDA3308C",
    x"BDA362A7",
    x"BDA394C2",
    x"BDA3C6DC",
    x"BDA3F8F7",
    x"BDA42B12",
    x"BDA45D2C",
    x"BDA48F47",
    x"BDA4C161",
    x"BDA4F37B",
    x"BDA52595",
    x"BDA557AF",
    x"BDA589C9",
    x"BDA5BBE3",
    x"BDA5EDFD",
    x"BDA62016",
    x"BDA65230",
    x"BDA68449",
    x"BDA6B663",
    x"BDA6E87C",
    x"BDA71A95",
    x"BDA74CAE",
    x"BDA77EC7",
    x"BDA7B0E0",
    x"BDA7E2F8",
    x"BDA81511",
    x"BDA84729",
    x"BDA87942",
    x"BDA8AB5A",
    x"BDA8DD72",
    x"BDA90F8A",
    x"BDA941A2",
    x"BDA973BA",
    x"BDA9A5D2",
    x"BDA9D7EA",
    x"BDAA0A01",
    x"BDAA3C19",
    x"BDAA6E30",
    x"BDAAA048",
    x"BDAAD25F",
    x"BDAB0476",
    x"BDAB368D",
    x"BDAB68A4",
    x"BDAB9ABA",
    x"BDABCCD1",
    x"BDABFEE8",
    x"BDAC30FE",
    x"BDAC6314",
    x"BDAC952B",
    x"BDACC741",
    x"BDACF957",
    x"BDAD2B6D",
    x"BDAD5D83",
    x"BDAD8F98",
    x"BDADC1AE",
    x"BDADF3C3",
    x"BDAE25D9",
    x"BDAE57EE",
    x"BDAE8A03",
    x"BDAEBC18",
    x"BDAEEE2D",
    x"BDAF2042",
    x"BDAF5257",
    x"BDAF846C",
    x"BDAFB680",
    x"BDAFE895",
    x"BDB01AA9",
    x"BDB04CBD",
    x"BDB07ED2",
    x"BDB0B0E6",
    x"BDB0E2FA",
    x"BDB1150D",
    x"BDB14721",
    x"BDB17935",
    x"BDB1AB48",
    x"BDB1DD5C",
    x"BDB20F6F",
    x"BDB24182",
    x"BDB27395",
    x"BDB2A5A8",
    x"BDB2D7BB",
    x"BDB309CE",
    x"BDB33BE0",
    x"BDB36DF3",
    x"BDB3A005",
    x"BDB3D218",
    x"BDB4042A",
    x"BDB4363C",
    x"BDB4684E",
    x"BDB49A60",
    x"BDB4CC72",
    x"BDB4FE83",
    x"BDB53095",
    x"BDB562A6",
    x"BDB594B8",
    x"BDB5C6C9",
    x"BDB5F8DA",
    x"BDB62AEB",
    x"BDB65CFC",
    x"BDB68F0D",
    x"BDB6C11D",
    x"BDB6F32E",
    x"BDB7253E",
    x"BDB7574F",
    x"BDB7895F",
    x"BDB7BB6F",
    x"BDB7ED7F",
    x"BDB81F8F",
    x"BDB8519F",
    x"BDB883AF",
    x"BDB8B5BE",
    x"BDB8E7CE",
    x"BDB919DD",
    x"BDB94BEC",
    x"BDB97DFB",
    x"BDB9B00A",
    x"BDB9E219",
    x"BDBA1428",
    x"BDBA4637",
    x"BDBA7845",
    x"BDBAAA54",
    x"BDBADC62",
    x"BDBB0E70",
    x"BDBB407E",
    x"BDBB728C",
    x"BDBBA49A",
    x"BDBBD6A8",
    x"BDBC08B6",
    x"BDBC3AC3",
    x"BDBC6CD1",
    x"BDBC9EDE",
    x"BDBCD0EB",
    x"BDBD02F8",
    x"BDBD3505",
    x"BDBD6712",
    x"BDBD991F",
    x"BDBDCB2C",
    x"BDBDFD38",
    x"BDBE2F45",
    x"BDBE6151",
    x"BDBE935D",
    x"BDBEC569",
    x"BDBEF775",
    x"BDBF2981",
    x"BDBF5B8D",
    x"BDBF8D98",
    x"BDBFBFA4",
    x"BDBFF1AF",
    x"BDC023BA",
    x"BDC055C6",
    x"BDC087D1",
    x"BDC0B9DC",
    x"BDC0EBE6",
    x"BDC11DF1",
    x"BDC14FFC",
    x"BDC18206",
    x"BDC1B410",
    x"BDC1E61B",
    x"BDC21825",
    x"BDC24A2F",
    x"BDC27C39",
    x"BDC2AE42",
    x"BDC2E04C",
    x"BDC31255",
    x"BDC3445F",
    x"BDC37668",
    x"BDC3A871",
    x"BDC3DA7A",
    x"BDC40C83",
    x"BDC43E8C",
    x"BDC47095",
    x"BDC4A29D",
    x"BDC4D4A6",
    x"BDC506AE",
    x"BDC538B6",
    x"BDC56ABE",
    x"BDC59CC6",
    x"BDC5CECE",
    x"BDC600D6",
    x"BDC632DE",
    x"BDC664E5",
    x"BDC696ED",
    x"BDC6C8F4",
    x"BDC6FAFB",
    x"BDC72D02",
    x"BDC75F09",
    x"BDC79110",
    x"BDC7C316",
    x"BDC7F51D",
    x"BDC82723",
    x"BDC8592A",
    x"BDC88B30",
    x"BDC8BD36",
    x"BDC8EF3C",
    x"BDC92142",
    x"BDC95347",
    x"BDC9854D",
    x"BDC9B752",
    x"BDC9E958",
    x"BDCA1B5D",
    x"BDCA4D62",
    x"BDCA7F67",
    x"BDCAB16C",
    x"BDCAE371",
    x"BDCB1575",
    x"BDCB477A",
    x"BDCB797E",
    x"BDCBAB82",
    x"BDCBDD86",
    x"BDCC0F8A",
    x"BDCC418E",
    x"BDCC7392",
    x"BDCCA596",
    x"BDCCD799",
    x"BDCD099C",
    x"BDCD3BA0",
    x"BDCD6DA3",
    x"BDCD9FA6",
    x"BDCDD1A9",
    x"BDCE03AB",
    x"BDCE35AE",
    x"BDCE67B1",
    x"BDCE99B3",
    x"BDCECBB5",
    x"BDCEFDB7",
    x"BDCF2FB9",
    x"BDCF61BB",
    x"BDCF93BD",
    x"BDCFC5BF",
    x"BDCFF7C0",
    x"BDD029C2",
    x"BDD05BC3",
    x"BDD08DC4",
    x"BDD0BFC5",
    x"BDD0F1C6",
    x"BDD123C7",
    x"BDD155C7",
    x"BDD187C8",
    x"BDD1B9C8",
    x"BDD1EBC8",
    x"BDD21DC8",
    x"BDD24FC8",
    x"BDD281C8",
    x"BDD2B3C8",
    x"BDD2E5C8",
    x"BDD317C7",
    x"BDD349C7",
    x"BDD37BC6",
    x"BDD3ADC5",
    x"BDD3DFC4",
    x"BDD411C3",
    x"BDD443C1",
    x"BDD475C0",
    x"BDD4A7BE",
    x"BDD4D9BD",
    x"BDD50BBB",
    x"BDD53DB9",
    x"BDD56FB7",
    x"BDD5A1B5",
    x"BDD5D3B3",
    x"BDD605B0",
    x"BDD637AE",
    x"BDD669AB",
    x"BDD69BA8",
    x"BDD6CDA5",
    x"BDD6FFA2",
    x"BDD7319F",
    x"BDD7639C",
    x"BDD79598",
    x"BDD7C795",
    x"BDD7F991",
    x"BDD82B8D",
    x"BDD85D89",
    x"BDD88F85",
    x"BDD8C181",
    x"BDD8F37C",
    x"BDD92578",
    x"BDD95773",
    x"BDD9896E",
    x"BDD9BB69",
    x"BDD9ED64",
    x"BDDA1F5F",
    x"BDDA515A",
    x"BDDA8354",
    x"BDDAB54F",
    x"BDDAE749",
    x"BDDB1943",
    x"BDDB4B3D",
    x"BDDB7D37",
    x"BDDBAF31",
    x"BDDBE12B",
    x"BDDC1324",
    x"BDDC451E",
    x"BDDC7717",
    x"BDDCA910",
    x"BDDCDB09",
    x"BDDD0D02",
    x"BDDD3EFB",
    x"BDDD70F3",
    x"BDDDA2EC",
    x"BDDDD4E4",
    x"BDDE06DC",
    x"BDDE38D4",
    x"BDDE6ACC",
    x"BDDE9CC4",
    x"BDDECEBC",
    x"BDDF00B3",
    x"BDDF32AB",
    x"BDDF64A2",
    x"BDDF9699",
    x"BDDFC890",
    x"BDDFFA87",
    x"BDE02C7D",
    x"BDE05E74",
    x"BDE0906A",
    x"BDE0C261",
    x"BDE0F457",
    x"BDE1264D",
    x"BDE15843",
    x"BDE18A39",
    x"BDE1BC2E",
    x"BDE1EE24",
    x"BDE22019",
    x"BDE2520E",
    x"BDE28403",
    x"BDE2B5F8",
    x"BDE2E7ED",
    x"BDE319E2",
    x"BDE34BD6",
    x"BDE37DCB",
    x"BDE3AFBF",
    x"BDE3E1B3",
    x"BDE413A7",
    x"BDE4459B",
    x"BDE4778F",
    x"BDE4A982",
    x"BDE4DB76",
    x"BDE50D69",
    x"BDE53F5C",
    x"BDE5714F",
    x"BDE5A342",
    x"BDE5D535",
    x"BDE60727",
    x"BDE6391A",
    x"BDE66B0C",
    x"BDE69CFE",
    x"BDE6CEF0",
    x"BDE700E2",
    x"BDE732D4",
    x"BDE764C6",
    x"BDE796B7",
    x"BDE7C8A9",
    x"BDE7FA9A",
    x"BDE82C8B",
    x"BDE85E7C",
    x"BDE8906D",
    x"BDE8C25D",
    x"BDE8F44E",
    x"BDE9263E",
    x"BDE9582E",
    x"BDE98A1F",
    x"BDE9BC0E",
    x"BDE9EDFE",
    x"BDEA1FEE",
    x"BDEA51DE",
    x"BDEA83CD",
    x"BDEAB5BC",
    x"BDEAE7AB",
    x"BDEB199A",
    x"BDEB4B89",
    x"BDEB7D78",
    x"BDEBAF66",
    x"BDEBE155",
    x"BDEC1343",
    x"BDEC4531",
    x"BDEC771F",
    x"BDECA90D",
    x"BDECDAFB",
    x"BDED0CE8",
    x"BDED3ED5",
    x"BDED70C3",
    x"BDEDA2B0",
    x"BDEDD49D",
    x"BDEE068A",
    x"BDEE3876",
    x"BDEE6A63",
    x"BDEE9C4F",
    x"BDEECE3C",
    x"BDEF0028",
    x"BDEF3214",
    x"BDEF63FF",
    x"BDEF95EB",
    x"BDEFC7D7",
    x"BDEFF9C2",
    x"BDF02BAD",
    x"BDF05D98",
    x"BDF08F83",
    x"BDF0C16E",
    x"BDF0F359",
    x"BDF12543",
    x"BDF1572E",
    x"BDF18918",
    x"BDF1BB02",
    x"BDF1ECEC",
    x"BDF21ED6",
    x"BDF250BF",
    x"BDF282A9",
    x"BDF2B492",
    x"BDF2E67C",
    x"BDF31865",
    x"BDF34A4E",
    x"BDF37C36",
    x"BDF3AE1F",
    x"BDF3E007",
    x"BDF411F0",
    x"BDF443D8",
    x"BDF475C0",
    x"BDF4A7A8",
    x"BDF4D990",
    x"BDF50B77",
    x"BDF53D5F",
    x"BDF56F46",
    x"BDF5A12D",
    x"BDF5D314",
    x"BDF604FB",
    x"BDF636E2",
    x"BDF668C8",
    x"BDF69AAF",
    x"BDF6CC95",
    x"BDF6FE7B",
    x"BDF73061",
    x"BDF76247",
    x"BDF7942C",
    x"BDF7C612",
    x"BDF7F7F7",
    x"BDF829DD",
    x"BDF85BC2",
    x"BDF88DA7",
    x"BDF8BF8B",
    x"BDF8F170",
    x"BDF92354",
    x"BDF95539",
    x"BDF9871D",
    x"BDF9B901",
    x"BDF9EAE5",
    x"BDFA1CC8",
    x"BDFA4EAC",
    x"BDFA808F",
    x"BDFAB273",
    x"BDFAE456",
    x"BDFB1639",
    x"BDFB481C",
    x"BDFB79FE",
    x"BDFBABE1",
    x"BDFBDDC3",
    x"BDFC0FA5",
    x"BDFC4187",
    x"BDFC7369",
    x"BDFCA54B",
    x"BDFCD72D",
    x"BDFD090E",
    x"BDFD3AEF",
    x"BDFD6CD1",
    x"BDFD9EB2",
    x"BDFDD092",
    x"BDFE0273",
    x"BDFE3454",
    x"BDFE6634",
    x"BDFE9814",
    x"BDFEC9F4",
    x"BDFEFBD4",
    x"BDFF2DB4",
    x"BDFF5F94",
    x"BDFF9173",
    x"BDFFC352",
    x"BDFFF531",
    x"BE001388",
    x"BE002C78",
    x"BE004567",
    x"BE005E56",
    x"BE007745",
    x"BE009035",
    x"BE00A924",
    x"BE00C213",
    x"BE00DB01",
    x"BE00F3F0",
    x"BE010CDF",
    x"BE0125CE",
    x"BE013EBC",
    x"BE0157AB",
    x"BE017099",
    x"BE018987",
    x"BE01A276",
    x"BE01BB64",
    x"BE01D452",
    x"BE01ED40",
    x"BE02062E",
    x"BE021F1C",
    x"BE02380A",
    x"BE0250F7",
    x"BE0269E5",
    x"BE0282D2",
    x"BE029BC0",
    x"BE02B4AD",
    x"BE02CD9B",
    x"BE02E688",
    x"BE02FF75",
    x"BE031862",
    x"BE03314F",
    x"BE034A3C",
    x"BE036329",
    x"BE037C16",
    x"BE039502",
    x"BE03ADEF",
    x"BE03C6DB",
    x"BE03DFC8",
    x"BE03F8B4",
    x"BE0411A0",
    x"BE042A8D",
    x"BE044379",
    x"BE045C65",
    x"BE047551",
    x"BE048E3D",
    x"BE04A729",
    x"BE04C014",
    x"BE04D900",
    x"BE04F1EB",
    x"BE050AD7",
    x"BE0523C2",
    x"BE053CAE",
    x"BE055599",
    x"BE056E84",
    x"BE05876F",
    x"BE05A05A",
    x"BE05B945",
    x"BE05D230",
    x"BE05EB1B",
    x"BE060405",
    x"BE061CF0",
    x"BE0635DB",
    x"BE064EC5",
    x"BE0667AF",
    x"BE06809A",
    x"BE069984",
    x"BE06B26E",
    x"BE06CB58",
    x"BE06E442",
    x"BE06FD2C",
    x"BE071616",
    x"BE072EFF",
    x"BE0747E9",
    x"BE0760D2",
    x"BE0779BC",
    x"BE0792A5",
    x"BE07AB8F",
    x"BE07C478",
    x"BE07DD61",
    x"BE07F64A",
    x"BE080F33",
    x"BE08281C",
    x"BE084105",
    x"BE0859ED",
    x"BE0872D6",
    x"BE088BBF",
    x"BE08A4A7",
    x"BE08BD90",
    x"BE08D678",
    x"BE08EF60",
    x"BE090848",
    x"BE092130",
    x"BE093A18",
    x"BE095300",
    x"BE096BE8",
    x"BE0984D0",
    x"BE099DB7",
    x"BE09B69F",
    x"BE09CF86",
    x"BE09E86E",
    x"BE0A0155",
    x"BE0A1A3C",
    x"BE0A3324",
    x"BE0A4C0B",
    x"BE0A64F2",
    x"BE0A7DD9",
    x"BE0A96BF",
    x"BE0AAFA6",
    x"BE0AC88D",
    x"BE0AE173",
    x"BE0AFA5A",
    x"BE0B1340",
    x"BE0B2C27",
    x"BE0B450D",
    x"BE0B5DF3",
    x"BE0B76D9",
    x"BE0B8FBF",
    x"BE0BA8A5",
    x"BE0BC18B",
    x"BE0BDA71",
    x"BE0BF356",
    x"BE0C0C3C",
    x"BE0C2521",
    x"BE0C3E07",
    x"BE0C56EC",
    x"BE0C6FD1",
    x"BE0C88B6",
    x"BE0CA19B",
    x"BE0CBA80",
    x"BE0CD365",
    x"BE0CEC4A",
    x"BE0D052F",
    x"BE0D1E13",
    x"BE0D36F8",
    x"BE0D4FDC",
    x"BE0D68C1",
    x"BE0D81A5",
    x"BE0D9A89",
    x"BE0DB36D",
    x"BE0DCC51",
    x"BE0DE535",
    x"BE0DFE19",
    x"BE0E16FD",
    x"BE0E2FE1",
    x"BE0E48C4",
    x"BE0E61A8",
    x"BE0E7A8B",
    x"BE0E936F",
    x"BE0EAC52",
    x"BE0EC535",
    x"BE0EDE18",
    x"BE0EF6FB",
    x"BE0F0FDE",
    x"BE0F28C1",
    x"BE0F41A4",
    x"BE0F5A86",
    x"BE0F7369",
    x"BE0F8C4B",
    x"BE0FA52E",
    x"BE0FBE10",
    x"BE0FD6F2",
    x"BE0FEFD5",
    x"BE1008B7",
    x"BE102199",
    x"BE103A7B",
    x"BE10535C",
    x"BE106C3E",
    x"BE108520",
    x"BE109E01",
    x"BE10B6E3",
    x"BE10CFC4",
    x"BE10E8A5",
    x"BE110186",
    x"BE111A68",
    x"BE113349",
    x"BE114C2A",
    x"BE11650A",
    x"BE117DEB",
    x"BE1196CC",
    x"BE11AFAC",
    x"BE11C88D",
    x"BE11E16D",
    x"BE11FA4E",
    x"BE12132E",
    x"BE122C0E",
    x"BE1244EE",
    x"BE125DCE",
    x"BE1276AE",
    x"BE128F8E",
    x"BE12A86D",
    x"BE12C14D",
    x"BE12DA2C",
    x"BE12F30C",
    x"BE130BEB",
    x"BE1324CA",
    x"BE133DAA",
    x"BE135689",
    x"BE136F68",
    x"BE138847",
    x"BE13A125",
    x"BE13BA04",
    x"BE13D2E3",
    x"BE13EBC1",
    x"BE1404A0",
    x"BE141D7E",
    x"BE14365C",
    x"BE144F3B",
    x"BE146819",
    x"BE1480F7",
    x"BE1499D5",
    x"BE14B2B2",
    x"BE14CB90",
    x"BE14E46E",
    x"BE14FD4B",
    x"BE151629",
    x"BE152F06",
    x"BE1547E4",
    x"BE1560C1",
    x"BE15799E",
    x"BE15927B",
    x"BE15AB58",
    x"BE15C435",
    x"BE15DD11",
    x"BE15F5EE",
    x"BE160ECB",
    x"BE1627A7",
    x"BE164083",
    x"BE165960",
    x"BE16723C",
    x"BE168B18",
    x"BE16A3F4",
    x"BE16BCD0",
    x"BE16D5AC",
    x"BE16EE88",
    x"BE170763",
    x"BE17203F",
    x"BE17391A",
    x"BE1751F6",
    x"BE176AD1",
    x"BE1783AC",
    x"BE179C87",
    x"BE17B562",
    x"BE17CE3D",
    x"BE17E718",
    x"BE17FFF3",
    x"BE1818CE",
    x"BE1831A8",
    x"BE184A83",
    x"BE18635D",
    x"BE187C37",
    x"BE189511",
    x"BE18ADEC",
    x"BE18C6C6",
    x"BE18DFA0",
    x"BE18F879",
    x"BE191153",
    x"BE192A2D",
    x"BE194306",
    x"BE195BE0",
    x"BE1974B9",
    x"BE198D92",
    x"BE19A66C",
    x"BE19BF45",
    x"BE19D81E",
    x"BE19F0F7",
    x"BE1A09CF",
    x"BE1A22A8",
    x"BE1A3B81",
    x"BE1A5459",
    x"BE1A6D32",
    x"BE1A860A",
    x"BE1A9EE2",
    x"BE1AB7BB",
    x"BE1AD093",
    x"BE1AE96B",
    x"BE1B0242",
    x"BE1B1B1A",
    x"BE1B33F2",
    x"BE1B4CCA",
    x"BE1B65A1",
    x"BE1B7E79",
    x"BE1B9750",
    x"BE1BB027",
    x"BE1BC8FE",
    x"BE1BE1D5",
    x"BE1BFAAC",
    x"BE1C1383",
    x"BE1C2C5A",
    x"BE1C4530",
    x"BE1C5E07",
    x"BE1C76DE",
    x"BE1C8FB4",
    x"BE1CA88A",
    x"BE1CC160",
    x"BE1CDA36",
    x"BE1CF30D",
    x"BE1D0BE2",
    x"BE1D24B8",
    x"BE1D3D8E",
    x"BE1D5664",
    x"BE1D6F39",
    x"BE1D880F",
    x"BE1DA0E4",
    x"BE1DB9B9",
    x"BE1DD28E",
    x"BE1DEB63",
    x"BE1E0438",
    x"BE1E1D0D",
    x"BE1E35E2",
    x"BE1E4EB7",
    x"BE1E678B",
    x"BE1E8060",
    x"BE1E9934",
    x"BE1EB208",
    x"BE1ECADD",
    x"BE1EE3B1",
    x"BE1EFC85",
    x"BE1F1559",
    x"BE1F2E2C",
    x"BE1F4700",
    x"BE1F5FD4",
    x"BE1F78A7",
    x"BE1F917B",
    x"BE1FAA4E",
    x"BE1FC321",
    x"BE1FDBF4",
    x"BE1FF4C8",
    x"BE200D9A",
    x"BE20266D",
    x"BE203F40",
    x"BE205813",
    x"BE2070E5",
    x"BE2089B8",
    x"BE20A28A",
    x"BE20BB5C",
    x"BE20D42F",
    x"BE20ED01",
    x"BE2105D3",
    x"BE211EA5",
    x"BE213776",
    x"BE215048",
    x"BE21691A",
    x"BE2181EB",
    x"BE219ABD",
    x"BE21B38E",
    x"BE21CC5F",
    x"BE21E530",
    x"BE21FE01",
    x"BE2216D2",
    x"BE222FA3",
    x"BE224874",
    x"BE226144",
    x"BE227A15",
    x"BE2292E5",
    x"BE22ABB6",
    x"BE22C486",
    x"BE22DD56",
    x"BE22F626",
    x"BE230EF6",
    x"BE2327C6",
    x"BE234095",
    x"BE235965",
    x"BE237235",
    x"BE238B04",
    x"BE23A3D3",
    x"BE23BCA3",
    x"BE23D572",
    x"BE23EE41",
    x"BE240710",
    x"BE241FDF",
    x"BE2438AD",
    x"BE24517C",
    x"BE246A4B",
    x"BE248319",
    x"BE249BE7",
    x"BE24B4B6",
    x"BE24CD84",
    x"BE24E652",
    x"BE24FF20",
    x"BE2517EE",
    x"BE2530BC",
    x"BE254989",
    x"BE256257",
    x"BE257B24",
    x"BE2593F2",
    x"BE25ACBF",
    x"BE25C58C",
    x"BE25DE59",
    x"BE25F726",
    x"BE260FF3",
    x"BE2628C0",
    x"BE26418C",
    x"BE265A59",
    x"BE267325",
    x"BE268BF2",
    x"BE26A4BE",
    x"BE26BD8A",
    x"BE26D656",
    x"BE26EF22",
    x"BE2707EE",
    x"BE2720BA",
    x"BE273985",
    x"BE275251",
    x"BE276B1C",
    x"BE2783E8",
    x"BE279CB3",
    x"BE27B57E",
    x"BE27CE49",
    x"BE27E714",
    x"BE27FFDF",
    x"BE2818AA",
    x"BE283174",
    x"BE284A3F",
    x"BE286309",
    x"BE287BD4",
    x"BE28949E",
    x"BE28AD68",
    x"BE28C632",
    x"BE28DEFC",
    x"BE28F7C6",
    x"BE291090",
    x"BE292959",
    x"BE294223",
    x"BE295AEC",
    x"BE2973B6",
    x"BE298C7F",
    x"BE29A548",
    x"BE29BE11",
    x"BE29D6DA",
    x"BE29EFA3",
    x"BE2A086B",
    x"BE2A2134",
    x"BE2A39FD",
    x"BE2A52C5",
    x"BE2A6B8D",
    x"BE2A8456",
    x"BE2A9D1E",
    x"BE2AB5E6",
    x"BE2ACEAE",
    x"BE2AE775",
    x"BE2B003D",
    x"BE2B1905",
    x"BE2B31CC",
    x"BE2B4A93",
    x"BE2B635B",
    x"BE2B7C22",
    x"BE2B94E9",
    x"BE2BADB0",
    x"BE2BC677",
    x"BE2BDF3E",
    x"BE2BF804",
    x"BE2C10CB",
    x"BE2C2991",
    x"BE2C4258",
    x"BE2C5B1E",
    x"BE2C73E4",
    x"BE2C8CAA",
    x"BE2CA570",
    x"BE2CBE36",
    x"BE2CD6FB",
    x"BE2CEFC1",
    x"BE2D0887",
    x"BE2D214C",
    x"BE2D3A11",
    x"BE2D52D6",
    x"BE2D6B9C",
    x"BE2D8461",
    x"BE2D9D25",
    x"BE2DB5EA",
    x"BE2DCEAF",
    x"BE2DE773",
    x"BE2E0038",
    x"BE2E18FC",
    x"BE2E31C1",
    x"BE2E4A85",
    x"BE2E6349",
    x"BE2E7C0D",
    x"BE2E94D1",
    x"BE2EAD94",
    x"BE2EC658",
    x"BE2EDF1B",
    x"BE2EF7DF",
    x"BE2F10A2",
    x"BE2F2965",
    x"BE2F4228",
    x"BE2F5AEB",
    x"BE2F73AE",
    x"BE2F8C71",
    x"BE2FA534",
    x"BE2FBDF6",
    x"BE2FD6B9",
    x"BE2FEF7B",
    x"BE30083D",
    x"BE302100",
    x"BE3039C2",
    x"BE305284",
    x"BE306B45",
    x"BE308407",
    x"BE309CC9",
    x"BE30B58A",
    x"BE30CE4C",
    x"BE30E70D",
    x"BE30FFCE",
    x"BE31188F",
    x"BE313150",
    x"BE314A11",
    x"BE3162D2",
    x"BE317B92",
    x"BE319453",
    x"BE31AD13",
    x"BE31C5D4",
    x"BE31DE94",
    x"BE31F754",
    x"BE321014",
    x"BE3228D4",
    x"BE324194",
    x"BE325A54",
    x"BE327313",
    x"BE328BD3",
    x"BE32A492",
    x"BE32BD51",
    x"BE32D610",
    x"BE32EECF",
    x"BE33078E",
    x"BE33204D",
    x"BE33390C",
    x"BE3351CB",
    x"BE336A89",
    x"BE338348",
    x"BE339C06",
    x"BE33B4C4",
    x"BE33CD82",
    x"BE33E640",
    x"BE33FEFE",
    x"BE3417BC",
    x"BE343079",
    x"BE344937",
    x"BE3461F4",
    x"BE347AB2",
    x"BE34936F",
    x"BE34AC2C",
    x"BE34C4E9",
    x"BE34DDA6",
    x"BE34F662",
    x"BE350F1F",
    x"BE3527DC",
    x"BE354098",
    x"BE355954",
    x"BE357211",
    x"BE358ACD",
    x"BE35A389",
    x"BE35BC45",
    x"BE35D501",
    x"BE35EDBC",
    x"BE360678",
    x"BE361F33",
    x"BE3637EF",
    x"BE3650AA",
    x"BE366965",
    x"BE368220",
    x"BE369ADB",
    x"BE36B396",
    x"BE36CC50",
    x"BE36E50B",
    x"BE36FDC5",
    x"BE371680",
    x"BE372F3A",
    x"BE3747F4",
    x"BE3760AE",
    x"BE377968",
    x"BE379222",
    x"BE37AADC",
    x"BE37C395",
    x"BE37DC4F",
    x"BE37F508",
    x"BE380DC1",
    x"BE38267A",
    x"BE383F33",
    x"BE3857EC",
    x"BE3870A5",
    x"BE38895E",
    x"BE38A217",
    x"BE38BACF",
    x"BE38D387",
    x"BE38EC40",
    x"BE3904F8",
    x"BE391DB0",
    x"BE393668",
    x"BE394F20",
    x"BE3967D7",
    x"BE39808F",
    x"BE399946",
    x"BE39B1FE",
    x"BE39CAB5",
    x"BE39E36C",
    x"BE39FC23",
    x"BE3A14DA",
    x"BE3A2D91",
    x"BE3A4647",
    x"BE3A5EFE",
    x"BE3A77B4",
    x"BE3A906B",
    x"BE3AA921",
    x"BE3AC1D7",
    x"BE3ADA8D",
    x"BE3AF343",
    x"BE3B0BF9",
    x"BE3B24AF",
    x"BE3B3D64",
    x"BE3B561A",
    x"BE3B6ECF",
    x"BE3B8784",
    x"BE3BA039",
    x"BE3BB8EE",
    x"BE3BD1A3",
    x"BE3BEA58",
    x"BE3C030D",
    x"BE3C1BC1",
    x"BE3C3476",
    x"BE3C4D2A",
    x"BE3C65DE",
    x"BE3C7E92",
    x"BE3C9746",
    x"BE3CAFFA",
    x"BE3CC8AE",
    x"BE3CE161",
    x"BE3CFA15",
    x"BE3D12C8",
    x"BE3D2B7C",
    x"BE3D442F",
    x"BE3D5CE2",
    x"BE3D7595",
    x"BE3D8E48",
    x"BE3DA6FA",
    x"BE3DBFAD",
    x"BE3DD860",
    x"BE3DF112",
    x"BE3E09C4",
    x"BE3E2276",
    x"BE3E3B28",
    x"BE3E53DA",
    x"BE3E6C8C",
    x"BE3E853E",
    x"BE3E9DEF",
    x"BE3EB6A1",
    x"BE3ECF52",
    x"BE3EE804",
    x"BE3F00B5",
    x"BE3F1966",
    x"BE3F3217",
    x"BE3F4AC7",
    x"BE3F6378",
    x"BE3F7C29",
    x"BE3F94D9",
    x"BE3FAD89",
    x"BE3FC639",
    x"BE3FDEEA",
    x"BE3FF79A",
    x"BE401049",
    x"BE4028F9",
    x"BE4041A9",
    x"BE405A58",
    x"BE407308",
    x"BE408BB7",
    x"BE40A466",
    x"BE40BD15",
    x"BE40D5C4",
    x"BE40EE73",
    x"BE410722",
    x"BE411FD0",
    x"BE41387F",
    x"BE41512D",
    x"BE4169DB",
    x"BE418289",
    x"BE419B37",
    x"BE41B3E5",
    x"BE41CC93",
    x"BE41E541",
    x"BE41FDEE",
    x"BE42169B",
    x"BE422F49",
    x"BE4247F6",
    x"BE4260A3",
    x"BE427950",
    x"BE4291FD",
    x"BE42AAAA",
    x"BE42C356",
    x"BE42DC03",
    x"BE42F4AF",
    x"BE430D5B",
    x"BE432607",
    x"BE433EB3",
    x"BE43575F",
    x"BE43700B",
    x"BE4388B7",
    x"BE43A162",
    x"BE43BA0E",
    x"BE43D2B9",
    x"BE43EB64",
    x"BE44040F",
    x"BE441CBA",
    x"BE443565",
    x"BE444E10",
    x"BE4466BA",
    x"BE447F65",
    x"BE44980F",
    x"BE44B0B9",
    x"BE44C963",
    x"BE44E20D",
    x"BE44FAB7",
    x"BE451361",
    x"BE452C0B",
    x"BE4544B4",
    x"BE455D5E",
    x"BE457607",
    x"BE458EB0",
    x"BE45A759",
    x"BE45C002",
    x"BE45D8AB",
    x"BE45F153",
    x"BE4609FC",
    x"BE4622A5",
    x"BE463B4D",
    x"BE4653F5",
    x"BE466C9D",
    x"BE468545",
    x"BE469DED",
    x"BE46B695",
    x"BE46CF3C",
    x"BE46E7E4",
    x"BE47008B",
    x"BE471932",
    x"BE4731DA",
    x"BE474A81",
    x"BE476328",
    x"BE477BCE",
    x"BE479475",
    x"BE47AD1B",
    x"BE47C5C2",
    x"BE47DE68",
    x"BE47F70E",
    x"BE480FB4",
    x"BE48285A",
    x"BE484100",
    x"BE4859A6",
    x"BE48724B",
    x"BE488AF1",
    x"BE48A396",
    x"BE48BC3B",
    x"BE48D4E0",
    x"BE48ED85",
    x"BE49062A",
    x"BE491ECF",
    x"BE493774",
    x"BE495018",
    x"BE4968BC",
    x"BE498161",
    x"BE499A05",
    x"BE49B2A9",
    x"BE49CB4D",
    x"BE49E3F0",
    x"BE49FC94",
    x"BE4A1538",
    x"BE4A2DDB",
    x"BE4A467E",
    x"BE4A5F21",
    x"BE4A77C4",
    x"BE4A9067",
    x"BE4AA90A",
    x"BE4AC1AD",
    x"BE4ADA4F",
    x"BE4AF2F2",
    x"BE4B0B94",
    x"BE4B2436",
    x"BE4B3CD8",
    x"BE4B557A",
    x"BE4B6E1C",
    x"BE4B86BE",
    x"BE4B9F5F",
    x"BE4BB801",
    x"BE4BD0A2",
    x"BE4BE943",
    x"BE4C01E4",
    x"BE4C1A85",
    x"BE4C3326",
    x"BE4C4BC7",
    x"BE4C6467",
    x"BE4C7D08",
    x"BE4C95A8",
    x"BE4CAE48",
    x"BE4CC6E8",
    x"BE4CDF88",
    x"BE4CF828",
    x"BE4D10C8",
    x"BE4D2967",
    x"BE4D4207",
    x"BE4D5AA6",
    x"BE4D7345",
    x"BE4D8BE4",
    x"BE4DA483",
    x"BE4DBD22",
    x"BE4DD5C1",
    x"BE4DEE60",
    x"BE4E06FE",
    x"BE4E1F9C",
    x"BE4E383B",
    x"BE4E50D9",
    x"BE4E6977",
    x"BE4E8215",
    x"BE4E9AB2",
    x"BE4EB350",
    x"BE4ECBED",
    x"BE4EE48B",
    x"BE4EFD28",
    x"BE4F15C5",
    x"BE4F2E62",
    x"BE4F46FF",
    x"BE4F5F9C",
    x"BE4F7838",
    x"BE4F90D5",
    x"BE4FA971",
    x"BE4FC20D",
    x"BE4FDAA9",
    x"BE4FF345",
    x"BE500BE1",
    x"BE50247D",
    x"BE503D19",
    x"BE5055B4",
    x"BE506E4F",
    x"BE5086EB",
    x"BE509F86",
    x"BE50B821",
    x"BE50D0BC",
    x"BE50E956",
    x"BE5101F1",
    x"BE511A8B",
    x"BE513326",
    x"BE514BC0",
    x"BE51645A",
    x"BE517CF4",
    x"BE51958E",
    x"BE51AE28",
    x"BE51C6C1",
    x"BE51DF5B",
    x"BE51F7F4",
    x"BE52108D",
    x"BE522926",
    x"BE5241BF",
    x"BE525A58",
    x"BE5272F1",
    x"BE528B89",
    x"BE52A422",
    x"BE52BCBA",
    x"BE52D552",
    x"BE52EDEA",
    x"BE530682",
    x"BE531F1A",
    x"BE5337B2",
    x"BE535049",
    x"BE5368E1",
    x"BE538178",
    x"BE539A0F",
    x"BE53B2A6",
    x"BE53CB3D",
    x"BE53E3D4",
    x"BE53FC6B",
    x"BE541501",
    x"BE542D98",
    x"BE54462E",
    x"BE545EC4",
    x"BE54775A",
    x"BE548FF0",
    x"BE54A886",
    x"BE54C11B",
    x"BE54D9B1",
    x"BE54F246",
    x"BE550ADC",
    x"BE552371",
    x"BE553C06",
    x"BE55549B",
    x"BE556D2F",
    x"BE5585C4",
    x"BE559E58",
    x"BE55B6ED",
    x"BE55CF81",
    x"BE55E815",
    x"BE5600A9",
    x"BE56193D",
    x"BE5631D1",
    x"BE564A64",
    x"BE5662F8",
    x"BE567B8B",
    x"BE56941E",
    x"BE56ACB1",
    x"BE56C544",
    x"BE56DDD7",
    x"BE56F66A",
    x"BE570EFC",
    x"BE57278F",
    x"BE574021",
    x"BE5758B3",
    x"BE577145",
    x"BE5789D7",
    x"BE57A269",
    x"BE57BAFB",
    x"BE57D38C",
    x"BE57EC1D",
    x"BE5804AF",
    x"BE581D40",
    x"BE5835D1",
    x"BE584E62",
    x"BE5866F2",
    x"BE587F83",
    x"BE589813",
    x"BE58B0A4",
    x"BE58C934",
    x"BE58E1C4",
    x"BE58FA54",
    x"BE5912E4",
    x"BE592B74",
    x"BE594403",
    x"BE595C93",
    x"BE597522",
    x"BE598DB1",
    x"BE59A640",
    x"BE59BECF",
    x"BE59D75E",
    x"BE59EFEC",
    x"BE5A087B",
    x"BE5A2109",
    x"BE5A3997",
    x"BE5A5226",
    x"BE5A6AB4",
    x"BE5A8341",
    x"BE5A9BCF",
    x"BE5AB45D",
    x"BE5ACCEA",
    x"BE5AE578",
    x"BE5AFE05",
    x"BE5B1692",
    x"BE5B2F1F",
    x"BE5B47AC",
    x"BE5B6038",
    x"BE5B78C5",
    x"BE5B9151",
    x"BE5BA9DD",
    x"BE5BC26A",
    x"BE5BDAF6",
    x"BE5BF381",
    x"BE5C0C0D",
    x"BE5C2499",
    x"BE5C3D24",
    x"BE5C55B0",
    x"BE5C6E3B",
    x"BE5C86C6",
    x"BE5C9F51",
    x"BE5CB7DC",
    x"BE5CD066",
    x"BE5CE8F1",
    x"BE5D017B",
    x"BE5D1A05",
    x"BE5D3290",
    x"BE5D4B1A",
    x"BE5D63A4",
    x"BE5D7C2D",
    x"BE5D94B7",
    x"BE5DAD40",
    x"BE5DC5CA",
    x"BE5DDE53",
    x"BE5DF6DC",
    x"BE5E0F65",
    x"BE5E27EE",
    x"BE5E4076",
    x"BE5E58FF",
    x"BE5E7187",
    x"BE5E8A10",
    x"BE5EA298",
    x"BE5EBB20",
    x"BE5ED3A8",
    x"BE5EEC2F",
    x"BE5F04B7",
    x"BE5F1D3E",
    x"BE5F35C6",
    x"BE5F4E4D",
    x"BE5F66D4",
    x"BE5F7F5B",
    x"BE5F97E2",
    x"BE5FB068",
    x"BE5FC8EF",
    x"BE5FE175",
    x"BE5FF9FC",
    x"BE601282",
    x"BE602B08",
    x"BE60438E",
    x"BE605C13",
    x"BE607499",
    x"BE608D1E",
    x"BE60A5A4",
    x"BE60BE29",
    x"BE60D6AE",
    x"BE60EF33",
    x"BE6107B8",
    x"BE61203C",
    x"BE6138C1",
    x"BE615145",
    x"BE6169C9",
    x"BE61824D",
    x"BE619AD1",
    x"BE61B355",
    x"BE61CBD9",
    x"BE61E45C",
    x"BE61FCE0",
    x"BE621563",
    x"BE622DE6",
    x"BE624669",
    x"BE625EEC",
    x"BE62776F",
    x"BE628FF1",
    x"BE62A874",
    x"BE62C0F6",
    x"BE62D978",
    x"BE62F1FA",
    x"BE630A7C",
    x"BE6322FE",
    x"BE633B80",
    x"BE635401",
    x"BE636C83",
    x"BE638504",
    x"BE639D85",
    x"BE63B606",
    x"BE63CE87",
    x"BE63E707",
    x"BE63FF88",
    x"BE641808",
    x"BE643089",
    x"BE644909",
    x"BE646189",
    x"BE647A09",
    x"BE649288",
    x"BE64AB08",
    x"BE64C387",
    x"BE64DC07",
    x"BE64F486",
    x"BE650D05",
    x"BE652584",
    x"BE653E02",
    x"BE655681",
    x"BE656F00",
    x"BE65877E",
    x"BE659FFC",
    x"BE65B87A",
    x"BE65D0F8",
    x"BE65E976",
    x"BE6601F3",
    x"BE661A71",
    x"BE6632EE",
    x"BE664B6C",
    x"BE6663E9",
    x"BE667C66",
    x"BE6694E2",
    x"BE66AD5F",
    x"BE66C5DC",
    x"BE66DE58",
    x"BE66F6D4",
    x"BE670F50",
    x"BE6727CC",
    x"BE674048",
    x"BE6758C4",
    x"BE67713F",
    x"BE6789BB",
    x"BE67A236",
    x"BE67BAB1",
    x"BE67D32C",
    x"BE67EBA7",
    x"BE680422",
    x"BE681C9C",
    x"BE683517",
    x"BE684D91",
    x"BE68660B",
    x"BE687E85",
    x"BE6896FF",
    x"BE68AF79",
    x"BE68C7F3",
    x"BE68E06C",
    x"BE68F8E5",
    x"BE69115F",
    x"BE6929D8",
    x"BE694251",
    x"BE695AC9",
    x"BE697342",
    x"BE698BBA",
    x"BE69A433",
    x"BE69BCAB",
    x"BE69D523",
    x"BE69ED9B",
    x"BE6A0613",
    x"BE6A1E8A",
    x"BE6A3702",
    x"BE6A4F79",
    x"BE6A67F0",
    x"BE6A8067",
    x"BE6A98DE",
    x"BE6AB155",
    x"BE6AC9CC",
    x"BE6AE242",
    x"BE6AFAB9",
    x"BE6B132F",
    x"BE6B2BA5",
    x"BE6B441B",
    x"BE6B5C91",
    x"BE6B7506",
    x"BE6B8D7C",
    x"BE6BA5F1",
    x"BE6BBE66",
    x"BE6BD6DC",
    x"BE6BEF51",
    x"BE6C07C5",
    x"BE6C203A",
    x"BE6C38AF",
    x"BE6C5123",
    x"BE6C6997",
    x"BE6C820B",
    x"BE6C9A7F",
    x"BE6CB2F3",
    x"BE6CCB67",
    x"BE6CE3DA",
    x"BE6CFC4E",
    x"BE6D14C1",
    x"BE6D2D34",
    x"BE6D45A7",
    x"BE6D5E1A",
    x"BE6D768C",
    x"BE6D8EFF",
    x"BE6DA771",
    x"BE6DBFE3",
    x"BE6DD856",
    x"BE6DF0C7",
    x"BE6E0939",
    x"BE6E21AB",
    x"BE6E3A1C",
    x"BE6E528E",
    x"BE6E6AFF",
    x"BE6E8370",
    x"BE6E9BE1",
    x"BE6EB452",
    x"BE6ECCC3",
    x"BE6EE533",
    x"BE6EFDA3",
    x"BE6F1614",
    x"BE6F2E84",
    x"BE6F46F4",
    x"BE6F5F63",
    x"BE6F77D3",
    x"BE6F9043",
    x"BE6FA8B2",
    x"BE6FC121",
    x"BE6FD990",
    x"BE6FF1FF",
    x"BE700A6E",
    x"BE7022DD",
    x"BE703B4B",
    x"BE7053B9",
    x"BE706C28",
    x"BE708496",
    x"BE709D04",
    x"BE70B571",
    x"BE70CDDF",
    x"BE70E64C",
    x"BE70FEBA",
    x"BE711727",
    x"BE712F94",
    x"BE714801",
    x"BE71606E",
    x"BE7178DA",
    x"BE719147",
    x"BE71A9B3",
    x"BE71C21F",
    x"BE71DA8B",
    x"BE71F2F7",
    x"BE720B63",
    x"BE7223CE",
    x"BE723C3A",
    x"BE7254A5",
    x"BE726D10",
    x"BE72857B",
    x"BE729DE6",
    x"BE72B651",
    x"BE72CEBC",
    x"BE72E726",
    x"BE72FF90",
    x"BE7317FA",
    x"BE733064",
    x"BE7348CE",
    x"BE736138",
    x"BE7379A1",
    x"BE73920B",
    x"BE73AA74",
    x"BE73C2DD",
    x"BE73DB46",
    x"BE73F3AF",
    x"BE740C18",
    x"BE742480",
    x"BE743CE8",
    x"BE745551",
    x"BE746DB9",
    x"BE748621",
    x"BE749E88",
    x"BE74B6F0",
    x"BE74CF57",
    x"BE74E7BF",
    x"BE750026",
    x"BE75188D",
    x"BE7530F4",
    x"BE75495B",
    x"BE7561C1",
    x"BE757A28",
    x"BE75928E",
    x"BE75AAF4",
    x"BE75C35A",
    x"BE75DBC0",
    x"BE75F426",
    x"BE760C8B",
    x"BE7624F1",
    x"BE763D56",
    x"BE7655BB",
    x"BE766E20",
    x"BE768685",
    x"BE769EEA",
    x"BE76B74E",
    x"BE76CFB2",
    x"BE76E817",
    x"BE77007B",
    x"BE7718DF",
    x"BE773142",
    x"BE7749A6",
    x"BE77620A",
    x"BE777A6D",
    x"BE7792D0",
    x"BE77AB33",
    x"BE77C396",
    x"BE77DBF9",
    x"BE77F45B",
    x"BE780CBE",
    x"BE782520",
    x"BE783D82",
    x"BE7855E4",
    x"BE786E46",
    x"BE7886A8",
    x"BE789F09",
    x"BE78B76B",
    x"BE78CFCC",
    x"BE78E82D",
    x"BE79008E",
    x"BE7918EF",
    x"BE79314F",
    x"BE7949B0",
    x"BE796210",
    x"BE797A70",
    x"BE7992D0",
    x"BE79AB30",
    x"BE79C390",
    x"BE79DBF0",
    x"BE79F44F",
    x"BE7A0CAE",
    x"BE7A250D",
    x"BE7A3D6C",
    x"BE7A55CB",
    x"BE7A6E2A",
    x"BE7A8688",
    x"BE7A9EE7",
    x"BE7AB745",
    x"BE7ACFA3",
    x"BE7AE801",
    x"BE7B005F",
    x"BE7B18BC",
    x"BE7B311A",
    x"BE7B4977",
    x"BE7B61D4",
    x"BE7B7A31",
    x"BE7B928E",
    x"BE7BAAEB",
    x"BE7BC348",
    x"BE7BDBA4",
    x"BE7BF400",
    x"BE7C0C5C",
    x"BE7C24B8",
    x"BE7C3D14",
    x"BE7C5570",
    x"BE7C6DCB",
    x"BE7C8627",
    x"BE7C9E82",
    x"BE7CB6DD",
    x"BE7CCF38",
    x"BE7CE793",
    x"BE7CFFED",
    x"BE7D1848",
    x"BE7D30A2",
    x"BE7D48FC",
    x"BE7D6156",
    x"BE7D79B0",
    x"BE7D9209",
    x"BE7DAA63",
    x"BE7DC2BC",
    x"BE7DDB16",
    x"BE7DF36F",
    x"BE7E0BC8",
    x"BE7E2420",
    x"BE7E3C79",
    x"BE7E54D1",
    x"BE7E6D2A",
    x"BE7E8582",
    x"BE7E9DDA",
    x"BE7EB632",
    x"BE7ECE89",
    x"BE7EE6E1",
    x"BE7EFF38",
    x"BE7F178F",
    x"BE7F2FE7",
    x"BE7F483D",
    x"BE7F6094",
    x"BE7F78EB",
    x"BE7F9141",
    x"BE7FA998",
    x"BE7FC1EE",
    x"BE7FDA44",
    x"BE7FF29A",
    x"BE800578",
    x"BE8011A2",
    x"BE801DCD",
    x"BE8029F8",
    x"BE803622",
    x"BE80424D",
    x"BE804E77",
    x"BE805AA1",
    x"BE8066CC",
    x"BE8072F6",
    x"BE807F20",
    x"BE808B4A",
    x"BE809774",
    x"BE80A39E",
    x"BE80AFC7",
    x"BE80BBF1",
    x"BE80C81B",
    x"BE80D444",
    x"BE80E06E",
    x"BE80EC97",
    x"BE80F8C0",
    x"BE8104E9",
    x"BE811113",
    x"BE811D3C",
    x"BE812965",
    x"BE81358E",
    x"BE8141B6",
    x"BE814DDF",
    x"BE815A08",
    x"BE816630",
    x"BE817259",
    x"BE817E81",
    x"BE818AAA",
    x"BE8196D2",
    x"BE81A2FA",
    x"BE81AF22",
    x"BE81BB4A",
    x"BE81C772",
    x"BE81D39A",
    x"BE81DFC2",
    x"BE81EBEA",
    x"BE81F811",
    x"BE820439",
    x"BE821060",
    x"BE821C88",
    x"BE8228AF",
    x"BE8234D7",
    x"BE8240FE",
    x"BE824D25",
    x"BE82594C",
    x"BE826573",
    x"BE82719A",
    x"BE827DC0",
    x"BE8289E7",
    x"BE82960E",
    x"BE82A234",
    x"BE82AE5B",
    x"BE82BA81",
    x"BE82C6A8",
    x"BE82D2CE",
    x"BE82DEF4",
    x"BE82EB1A",
    x"BE82F740",
    x"BE830366",
    x"BE830F8C",
    x"BE831BB2",
    x"BE8327D7",
    x"BE8333FD",
    x"BE834022",
    x"BE834C48",
    x"BE83586D",
    x"BE836493",
    x"BE8370B8",
    x"BE837CDD",
    x"BE838902",
    x"BE839527",
    x"BE83A14C",
    x"BE83AD71",
    x"BE83B995",
    x"BE83C5BA",
    x"BE83D1DF",
    x"BE83DE03",
    x"BE83EA28",
    x"BE83F64C",
    x"BE840270",
    x"BE840E94",
    x"BE841AB8",
    x"BE8426DD",
    x"BE843300",
    x"BE843F24",
    x"BE844B48",
    x"BE84576C",
    x"BE84638F",
    x"BE846FB3",
    x"BE847BD6",
    x"BE8487FA",
    x"BE84941D",
    x"BE84A040",
    x"BE84AC64",
    x"BE84B887",
    x"BE84C4AA",
    x"BE84D0CC",
    x"BE84DCEF",
    x"BE84E912",
    x"BE84F535",
    x"BE850157",
    x"BE850D7A",
    x"BE85199C",
    x"BE8525BF",
    x"BE8531E1",
    x"BE853E03",
    x"BE854A25",
    x"BE855647",
    x"BE856269",
    x"BE856E8B",
    x"BE857AAD",
    x"BE8586CE",
    x"BE8592F0",
    x"BE859F12",
    x"BE85AB33",
    x"BE85B755",
    x"BE85C376",
    x"BE85CF97",
    x"BE85DBB8",
    x"BE85E7D9",
    x"BE85F3FA",
    x"BE86001B",
    x"BE860C3C",
    x"BE86185D",
    x"BE86247D",
    x"BE86309E",
    x"BE863CBE",
    x"BE8648DF",
    x"BE8654FF",
    x"BE86611F",
    x"BE866D40",
    x"BE867960",
    x"BE868580",
    x"BE8691A0",
    x"BE869DBF",
    x"BE86A9DF",
    x"BE86B5FF",
    x"BE86C21F",
    x"BE86CE3E",
    x"BE86DA5D",
    x"BE86E67D",
    x"BE86F29C",
    x"BE86FEBB",
    x"BE870ADA",
    x"BE8716F9",
    x"BE872318",
    x"BE872F37",
    x"BE873B56",
    x"BE874775",
    x"BE875393",
    x"BE875FB2",
    x"BE876BD0",
    x"BE8777EF",
    x"BE87840D",
    x"BE87902B",
    x"BE879C49",
    x"BE87A868",
    x"BE87B486",
    x"BE87C0A3",
    x"BE87CCC1",
    x"BE87D8DF",
    x"BE87E4FD",
    x"BE87F11A",
    x"BE87FD38",
    x"BE880955",
    x"BE881572",
    x"BE882190",
    x"BE882DAD",
    x"BE8839CA",
    x"BE8845E7",
    x"BE885204",
    x"BE885E21",
    x"BE886A3D",
    x"BE88765A",
    x"BE888277",
    x"BE888E93",
    x"BE889AB0",
    x"BE88A6CC",
    x"BE88B2E8",
    x"BE88BF04",
    x"BE88CB20",
    x"BE88D73C",
    x"BE88E358",
    x"BE88EF74",
    x"BE88FB90",
    x"BE8907AC",
    x"BE8913C7",
    x"BE891FE3",
    x"BE892BFE",
    x"BE893819",
    x"BE894435",
    x"BE895050",
    x"BE895C6B",
    x"BE896886",
    x"BE8974A1",
    x"BE8980BC",
    x"BE898CD7",
    x"BE8998F1",
    x"BE89A50C",
    x"BE89B126",
    x"BE89BD41",
    x"BE89C95B",
    x"BE89D575",
    x"BE89E190",
    x"BE89EDAA",
    x"BE89F9C4",
    x"BE8A05DE",
    x"BE8A11F7",
    x"BE8A1E11",
    x"BE8A2A2B",
    x"BE8A3645",
    x"BE8A425E",
    x"BE8A4E78",
    x"BE8A5A91",
    x"BE8A66AA",
    x"BE8A72C3",
    x"BE8A7EDC",
    x"BE8A8AF5",
    x"BE8A970E",
    x"BE8AA327",
    x"BE8AAF40",
    x"BE8ABB59",
    x"BE8AC771",
    x"BE8AD38A",
    x"BE8ADFA2",
    x"BE8AEBBB",
    x"BE8AF7D3",
    x"BE8B03EB",
    x"BE8B1003",
    x"BE8B1C1B",
    x"BE8B2833",
    x"BE8B344B",
    x"BE8B4063",
    x"BE8B4C7A",
    x"BE8B5892",
    x"BE8B64AA",
    x"BE8B70C1",
    x"BE8B7CD8",
    x"BE8B88F0",
    x"BE8B9507",
    x"BE8BA11E",
    x"BE8BAD35",
    x"BE8BB94C",
    x"BE8BC563",
    x"BE8BD179",
    x"BE8BDD90",
    x"BE8BE9A7",
    x"BE8BF5BD",
    x"BE8C01D4",
    x"BE8C0DEA",
    x"BE8C1A00",
    x"BE8C2616",
    x"BE8C322C",
    x"BE8C3E42",
    x"BE8C4A58",
    x"BE8C566E",
    x"BE8C6284",
    x"BE8C6E9A",
    x"BE8C7AAF",
    x"BE8C86C5",
    x"BE8C92DA",
    x"BE8C9EEF",
    x"BE8CAB05",
    x"BE8CB71A",
    x"BE8CC32F",
    x"BE8CCF44",
    x"BE8CDB59",
    x"BE8CE76D",
    x"BE8CF382",
    x"BE8CFF97",
    x"BE8D0BAB",
    x"BE8D17C0",
    x"BE8D23D4",
    x"BE8D2FE9",
    x"BE8D3BFD",
    x"BE8D4811",
    x"BE8D5425",
    x"BE8D6039",
    x"BE8D6C4D",
    x"BE8D7861",
    x"BE8D8474",
    x"BE8D9088",
    x"BE8D9C9B",
    x"BE8DA8AF",
    x"BE8DB4C2",
    x"BE8DC0D6",
    x"BE8DCCE9",
    x"BE8DD8FC",
    x"BE8DE50F",
    x"BE8DF122",
    x"BE8DFD35",
    x"BE8E0947",
    x"BE8E155A",
    x"BE8E216D",
    x"BE8E2D7F",
    x"BE8E3992",
    x"BE8E45A4",
    x"BE8E51B6",
    x"BE8E5DC8",
    x"BE8E69DB",
    x"BE8E75ED",
    x"BE8E81FE",
    x"BE8E8E10",
    x"BE8E9A22",
    x"BE8EA634",
    x"BE8EB245",
    x"BE8EBE57",
    x"BE8ECA68",
    x"BE8ED679",
    x"BE8EE28B",
    x"BE8EEE9C",
    x"BE8EFAAD",
    x"BE8F06BE",
    x"BE8F12CF",
    x"BE8F1EDF",
    x"BE8F2AF0",
    x"BE8F3701",
    x"BE8F4311",
    x"BE8F4F22",
    x"BE8F5B32",
    x"BE8F6742",
    x"BE8F7353",
    x"BE8F7F63",
    x"BE8F8B73",
    x"BE8F9783",
    x"BE8FA392",
    x"BE8FAFA2",
    x"BE8FBBB2",
    x"BE8FC7C1",
    x"BE8FD3D1",
    x"BE8FDFE0",
    x"BE8FEBF0",
    x"BE8FF7FF",
    x"BE90040E",
    x"BE90101D",
    x"BE901C2C",
    x"BE90283B",
    x"BE90344A",
    x"BE904059",
    x"BE904C67",
    x"BE905876",
    x"BE906484",
    x"BE907093",
    x"BE907CA1",
    x"BE9088AF",
    x"BE9094BD",
    x"BE90A0CB",
    x"BE90ACD9",
    x"BE90B8E7",
    x"BE90C4F5",
    x"BE90D102",
    x"BE90DD10",
    x"BE90E91D",
    x"BE90F52B",
    x"BE910138",
    x"BE910D45",
    x"BE911953",
    x"BE912560",
    x"BE91316D",
    x"BE913D79",
    x"BE914986",
    x"BE915593",
    x"BE9161A0",
    x"BE916DAC",
    x"BE9179B9",
    x"BE9185C5",
    x"BE9191D1",
    x"BE919DDD",
    x"BE91A9E9",
    x"BE91B5F5",
    x"BE91C201",
    x"BE91CE0D",
    x"BE91DA19",
    x"BE91E625",
    x"BE91F230",
    x"BE91FE3C",
    x"BE920A47",
    x"BE921652",
    x"BE92225E",
    x"BE922E69",
    x"BE923A74",
    x"BE92467F",
    x"BE92528A",
    x"BE925E94",
    x"BE926A9F",
    x"BE9276AA",
    x"BE9282B4",
    x"BE928EBF",
    x"BE929AC9",
    x"BE92A6D3",
    x"BE92B2DD",
    x"BE92BEE7",
    x"BE92CAF1",
    x"BE92D6FB",
    x"BE92E305",
    x"BE92EF0F",
    x"BE92FB18",
    x"BE930722",
    x"BE93132B",
    x"BE931F35",
    x"BE932B3E",
    x"BE933747",
    x"BE934350",
    x"BE934F59",
    x"BE935B62",
    x"BE93676B",
    x"BE937374",
    x"BE937F7D",
    x"BE938B85",
    x"BE93978E",
    x"BE93A396",
    x"BE93AF9E",
    x"BE93BBA6",
    x"BE93C7AF",
    x"BE93D3B7",
    x"BE93DFBF",
    x"BE93EBC6",
    x"BE93F7CE",
    x"BE9403D6",
    x"BE940FDD",
    x"BE941BE5",
    x"BE9427EC",
    x"BE9433F4",
    x"BE943FFB",
    x"BE944C02",
    x"BE945809",
    x"BE946410",
    x"BE947017",
    x"BE947C1E",
    x"BE948824",
    x"BE94942B",
    x"BE94A031",
    x"BE94AC38",
    x"BE94B83E",
    x"BE94C444",
    x"BE94D04B",
    x"BE94DC51",
    x"BE94E857",
    x"BE94F45D",
    x"BE950062",
    x"BE950C68",
    x"BE95186E",
    x"BE952473",
    x"BE953079",
    x"BE953C7E",
    x"BE954883",
    x"BE955488",
    x"BE95608D",
    x"BE956C92",
    x"BE957897",
    x"BE95849C",
    x"BE9590A1",
    x"BE959CA6",
    x"BE95A8AA",
    x"BE95B4AE",
    x"BE95C0B3",
    x"BE95CCB7",
    x"BE95D8BB",
    x"BE95E4BF",
    x"BE95F0C3",
    x"BE95FCC7",
    x"BE9608CB",
    x"BE9614CF",
    x"BE9620D2",
    x"BE962CD6",
    x"BE9638D9",
    x"BE9644DD",
    x"BE9650E0",
    x"BE965CE3",
    x"BE9668E6",
    x"BE9674E9",
    x"BE9680EC",
    x"BE968CEF",
    x"BE9698F2",
    x"BE96A4F4",
    x"BE96B0F7",
    x"BE96BCF9",
    x"BE96C8FC",
    x"BE96D4FE",
    x"BE96E100",
    x"BE96ED02",
    x"BE96F904",
    x"BE970506",
    x"BE971108",
    x"BE971D0A",
    x"BE97290B",
    x"BE97350D",
    x"BE97410E",
    x"BE974D10",
    x"BE975911",
    x"BE976512",
    x"BE977113",
    x"BE977D14",
    x"BE978915",
    x"BE979516",
    x"BE97A117",
    x"BE97AD17",
    x"BE97B918",
    x"BE97C518",
    x"BE97D119",
    x"BE97DD19",
    x"BE97E919",
    x"BE97F519",
    x"BE980119",
    x"BE980D19",
    x"BE981919",
    x"BE982519",
    x"BE983118",
    x"BE983D18",
    x"BE984917",
    x"BE985517",
    x"BE986116",
    x"BE986D15",
    x"BE987914",
    x"BE988513",
    x"BE989112",
    x"BE989D11",
    x"BE98A910",
    x"BE98B50E",
    x"BE98C10D",
    x"BE98CD0B",
    x"BE98D90A",
    x"BE98E508",
    x"BE98F106",
    x"BE98FD04",
    x"BE990902",
    x"BE991500",
    x"BE9920FE",
    x"BE992CFB",
    x"BE9938F9",
    x"BE9944F7",
    x"BE9950F4",
    x"BE995CF1",
    x"BE9968EE",
    x"BE9974EC",
    x"BE9980E9",
    x"BE998CE6",
    x"BE9998E3",
    x"BE99A4DF",
    x"BE99B0DC",
    x"BE99BCD9",
    x"BE99C8D5",
    x"BE99D4D1",
    x"BE99E0CE",
    x"BE99ECCA",
    x"BE99F8C6",
    x"BE9A04C2",
    x"BE9A10BE",
    x"BE9A1CBA",
    x"BE9A28B6",
    x"BE9A34B1",
    x"BE9A40AD",
    x"BE9A4CA8",
    x"BE9A58A4",
    x"BE9A649F",
    x"BE9A709A",
    x"BE9A7C95",
    x"BE9A8890",
    x"BE9A948B",
    x"BE9AA086",
    x"BE9AAC81",
    x"BE9AB87B",
    x"BE9AC476",
    x"BE9AD070",
    x"BE9ADC6B",
    x"BE9AE865",
    x"BE9AF45F",
    x"BE9B0059",
    x"BE9B0C53",
    x"BE9B184D",
    x"BE9B2447",
    x"BE9B3041",
    x"BE9B3C3A",
    x"BE9B4834",
    x"BE9B542D",
    x"BE9B6027",
    x"BE9B6C20",
    x"BE9B7819",
    x"BE9B8412",
    x"BE9B900B",
    x"BE9B9C04",
    x"BE9BA7FD",
    x"BE9BB3F5",
    x"BE9BBFEE",
    x"BE9BCBE6",
    x"BE9BD7DF",
    x"BE9BE3D7",
    x"BE9BEFCF",
    x"BE9BFBC7",
    x"BE9C07BF",
    x"BE9C13B7",
    x"BE9C1FAF",
    x"BE9C2BA7",
    x"BE9C379E",
    x"BE9C4396",
    x"BE9C4F8D",
    x"BE9C5B85",
    x"BE9C677C",
    x"BE9C7373",
    x"BE9C7F6A",
    x"BE9C8B61",
    x"BE9C9758",
    x"BE9CA34F",
    x"BE9CAF46",
    x"BE9CBB3C",
    x"BE9CC733",
    x"BE9CD329",
    x"BE9CDF20",
    x"BE9CEB16",
    x"BE9CF70C",
    x"BE9D0302",
    x"BE9D0EF8",
    x"BE9D1AEE",
    x"BE9D26E3",
    x"BE9D32D9",
    x"BE9D3ECF",
    x"BE9D4AC4",
    x"BE9D56BA",
    x"BE9D62AF",
    x"BE9D6EA4",
    x"BE9D7A99",
    x"BE9D868E",
    x"BE9D9283",
    x"BE9D9E78",
    x"BE9DAA6D",
    x"BE9DB661",
    x"BE9DC256",
    x"BE9DCE4A",
    x"BE9DDA3E",
    x"BE9DE633",
    x"BE9DF227",
    x"BE9DFE1B",
    x"BE9E0A0F",
    x"BE9E1603",
    x"BE9E21F6",
    x"BE9E2DEA",
    x"BE9E39DE",
    x"BE9E45D1",
    x"BE9E51C4",
    x"BE9E5DB8",
    x"BE9E69AB",
    x"BE9E759E",
    x"BE9E8191",
    x"BE9E8D84",
    x"BE9E9977",
    x"BE9EA569",
    x"BE9EB15C",
    x"BE9EBD4F",
    x"BE9EC941",
    x"BE9ED533",
    x"BE9EE126",
    x"BE9EED18",
    x"BE9EF90A",
    x"BE9F04FC",
    x"BE9F10EE",
    x"BE9F1CDF",
    x"BE9F28D1",
    x"BE9F34C3",
    x"BE9F40B4",
    x"BE9F4CA5",
    x"BE9F5897",
    x"BE9F6488",
    x"BE9F7079",
    x"BE9F7C6A",
    x"BE9F885B",
    x"BE9F944C",
    x"BE9FA03C",
    x"BE9FAC2D",
    x"BE9FB81D",
    x"BE9FC40E",
    x"BE9FCFFE",
    x"BE9FDBEE",
    x"BE9FE7DE",
    x"BE9FF3CE",
    x"BE9FFFBE",
    x"BEA00BAE",
    x"BEA0179E",
    x"BEA0238E",
    x"BEA02F7D",
    x"BEA03B6D",
    x"BEA0475C",
    x"BEA0534B",
    x"BEA05F3A",
    x"BEA06B29",
    x"BEA07718",
    x"BEA08307",
    x"BEA08EF6",
    x"BEA09AE5",
    x"BEA0A6D3",
    x"BEA0B2C2",
    x"BEA0BEB0",
    x"BEA0CA9E",
    x"BEA0D68D",
    x"BEA0E27B",
    x"BEA0EE69",
    x"BEA0FA57",
    x"BEA10644",
    x"BEA11232",
    x"BEA11E20",
    x"BEA12A0D",
    x"BEA135FB",
    x"BEA141E8",
    x"BEA14DD5",
    x"BEA159C2",
    x"BEA165AF",
    x"BEA1719C",
    x"BEA17D89",
    x"BEA18976",
    x"BEA19562",
    x"BEA1A14F",
    x"BEA1AD3B",
    x"BEA1B928",
    x"BEA1C514",
    x"BEA1D100",
    x"BEA1DCEC",
    x"BEA1E8D8",
    x"BEA1F4C4",
    x"BEA200B0",
    x"BEA20C9B",
    x"BEA21887",
    x"BEA22472",
    x"BEA2305E",
    x"BEA23C49",
    x"BEA24834",
    x"BEA2541F",
    x"BEA2600A",
    x"BEA26BF5",
    x"BEA277E0",
    x"BEA283CB",
    x"BEA28FB5",
    x"BEA29BA0",
    x"BEA2A78A",
    x"BEA2B374",
    x"BEA2BF5E",
    x"BEA2CB49",
    x"BEA2D733",
    x"BEA2E31C",
    x"BEA2EF06",
    x"BEA2FAF0",
    x"BEA306DA",
    x"BEA312C3",
    x"BEA31EAD",
    x"BEA32A96",
    x"BEA3367F",
    x"BEA34268",
    x"BEA34E51",
    x"BEA35A3A",
    x"BEA36623",
    x"BEA3720C",
    x"BEA37DF4",
    x"BEA389DD",
    x"BEA395C5",
    x"BEA3A1AD",
    x"BEA3AD96",
    x"BEA3B97E",
    x"BEA3C566",
    x"BEA3D14E",
    x"BEA3DD36",
    x"BEA3E91D",
    x"BEA3F505",
    x"BEA400ED",
    x"BEA40CD4",
    x"BEA418BB",
    x"BEA424A3",
    x"BEA4308A",
    x"BEA43C71",
    x"BEA44858",
    x"BEA4543F",
    x"BEA46025",
    x"BEA46C0C",
    x"BEA477F2",
    x"BEA483D9",
    x"BEA48FBF",
    x"BEA49BA6",
    x"BEA4A78C",
    x"BEA4B372",
    x"BEA4BF58",
    x"BEA4CB3E",
    x"BEA4D723",
    x"BEA4E309",
    x"BEA4EEEE",
    x"BEA4FAD4",
    x"BEA506B9",
    x"BEA5129F",
    x"BEA51E84",
    x"BEA52A69",
    x"BEA5364E",
    x"BEA54233",
    x"BEA54E17",
    x"BEA559FC",
    x"BEA565E1",
    x"BEA571C5",
    x"BEA57DA9",
    x"BEA5898E",
    x"BEA59572",
    x"BEA5A156",
    x"BEA5AD3A",
    x"BEA5B91E",
    x"BEA5C501",
    x"BEA5D0E5",
    x"BEA5DCC9",
    x"BEA5E8AC",
    x"BEA5F48F",
    x"BEA60073",
    x"BEA60C56",
    x"BEA61839",
    x"BEA6241C",
    x"BEA62FFF",
    x"BEA63BE2",
    x"BEA647C4",
    x"BEA653A7",
    x"BEA65F89",
    x"BEA66B6C",
    x"BEA6774E",
    x"BEA68330",
    x"BEA68F12",
    x"BEA69AF4",
    x"BEA6A6D6",
    x"BEA6B2B8",
    x"BEA6BE99",
    x"BEA6CA7B",
    x"BEA6D65C",
    x"BEA6E23E",
    x"BEA6EE1F",
    x"BEA6FA00",
    x"BEA705E1",
    x"BEA711C2",
    x"BEA71DA3",
    x"BEA72984",
    x"BEA73564",
    x"BEA74145",
    x"BEA74D25",
    x"BEA75906",
    x"BEA764E6",
    x"BEA770C6",
    x"BEA77CA6",
    x"BEA78886",
    x"BEA79466",
    x"BEA7A046",
    x"BEA7AC25",
    x"BEA7B805",
    x"BEA7C3E4",
    x"BEA7CFC4",
    x"BEA7DBA3",
    x"BEA7E782",
    x"BEA7F361",
    x"BEA7FF40",
    x"BEA80B1F",
    x"BEA816FE",
    x"BEA822DC",
    x"BEA82EBB",
    x"BEA83A99",
    x"BEA84678",
    x"BEA85256",
    x"BEA85E34",
    x"BEA86A12",
    x"BEA875F0",
    x"BEA881CE",
    x"BEA88DAB",
    x"BEA89989",
    x"BEA8A567",
    x"BEA8B144",
    x"BEA8BD21",
    x"BEA8C8FE",
    x"BEA8D4DC",
    x"BEA8E0B9",
    x"BEA8EC95",
    x"BEA8F872",
    x"BEA9044F",
    x"BEA9102C",
    x"BEA91C08",
    x"BEA927E5",
    x"BEA933C1",
    x"BEA93F9D",
    x"BEA94B79",
    x"BEA95755",
    x"BEA96331",
    x"BEA96F0D",
    x"BEA97AE8",
    x"BEA986C4",
    x"BEA992A0",
    x"BEA99E7B",
    x"BEA9AA56",
    x"BEA9B631",
    x"BEA9C20C",
    x"BEA9CDE7",
    x"BEA9D9C2",
    x"BEA9E59D",
    x"BEA9F178",
    x"BEA9FD52",
    x"BEAA092D",
    x"BEAA1507",
    x"BEAA20E1",
    x"BEAA2CBB",
    x"BEAA3895",
    x"BEAA446F",
    x"BEAA5049",
    x"BEAA5C23",
    x"BEAA67FD",
    x"BEAA73D6",
    x"BEAA7FB0",
    x"BEAA8B89",
    x"BEAA9762",
    x"BEAAA33B",
    x"BEAAAF14",
    x"BEAABAED",
    x"BEAAC6C6",
    x"BEAAD29F",
    x"BEAADE77",
    x"BEAAEA50",
    x"BEAAF628",
    x"BEAB0201",
    x"BEAB0DD9",
    x"BEAB19B1",
    x"BEAB2589",
    x"BEAB3161",
    x"BEAB3D39",
    x"BEAB4910",
    x"BEAB54E8",
    x"BEAB60BF",
    x"BEAB6C97",
    x"BEAB786E",
    x"BEAB8445",
    x"BEAB901C",
    x"BEAB9BF3",
    x"BEABA7CA",
    x"BEABB3A1",
    x"BEABBF77",
    x"BEABCB4E",
    x"BEABD724",
    x"BEABE2FB",
    x"BEABEED1",
    x"BEABFAA7",
    x"BEAC067D",
    x"BEAC1253",
    x"BEAC1E29",
    x"BEAC29FF",
    x"BEAC35D4",
    x"BEAC41AA",
    x"BEAC4D7F",
    x"BEAC5954",
    x"BEAC652A",
    x"BEAC70FF",
    x"BEAC7CD4",
    x"BEAC88A9",
    x"BEAC947D",
    x"BEACA052",
    x"BEACAC27",
    x"BEACB7FB",
    x"BEACC3CF",
    x"BEACCFA4",
    x"BEACDB78",
    x"BEACE74C",
    x"BEACF320",
    x"BEACFEF4",
    x"BEAD0AC7",
    x"BEAD169B",
    x"BEAD226F",
    x"BEAD2E42",
    x"BEAD3A15",
    x"BEAD45E9",
    x"BEAD51BC",
    x"BEAD5D8F",
    x"BEAD6962",
    x"BEAD7534",
    x"BEAD8107",
    x"BEAD8CDA",
    x"BEAD98AC",
    x"BEADA47F",
    x"BEADB051",
    x"BEADBC23",
    x"BEADC7F5",
    x"BEADD3C7",
    x"BEADDF99",
    x"BEADEB6B",
    x"BEADF73C",
    x"BEAE030E",
    x"BEAE0EDF",
    x"BEAE1AB1",
    x"BEAE2682",
    x"BEAE3253",
    x"BEAE3E24",
    x"BEAE49F5",
    x"BEAE55C6",
    x"BEAE6197",
    x"BEAE6D67",
    x"BEAE7938",
    x"BEAE8508",
    x"BEAE90D8",
    x"BEAE9CA8",
    x"BEAEA879",
    x"BEAEB449",
    x"BEAEC018",
    x"BEAECBE8",
    x"BEAED7B8",
    x"BEAEE387",
    x"BEAEEF57",
    x"BEAEFB26",
    x"BEAF06F5",
    x"BEAF12C5",
    x"BEAF1E94",
    x"BEAF2A62",
    x"BEAF3631",
    x"BEAF4200",
    x"BEAF4DCF",
    x"BEAF599D",
    x"BEAF656B",
    x"BEAF713A",
    x"BEAF7D08",
    x"BEAF88D6",
    x"BEAF94A4",
    x"BEAFA072",
    x"BEAFAC40",
    x"BEAFB80D",
    x"BEAFC3DB",
    x"BEAFCFA8",
    x"BEAFDB76",
    x"BEAFE743",
    x"BEAFF310",
    x"BEAFFEDD",
    x"BEB00AAA",
    x"BEB01677",
    x"BEB02243",
    x"BEB02E10",
    x"BEB039DC",
    x"BEB045A9",
    x"BEB05175",
    x"BEB05D41",
    x"BEB0690D",
    x"BEB074D9",
    x"BEB080A5",
    x"BEB08C71",
    x"BEB0983C",
    x"BEB0A408",
    x"BEB0AFD3",
    x"BEB0BB9F",
    x"BEB0C76A",
    x"BEB0D335",
    x"BEB0DF00",
    x"BEB0EACB",
    x"BEB0F696",
    x"BEB10260",
    x"BEB10E2B",
    x"BEB119F5",
    x"BEB125C0",
    x"BEB1318A",
    x"BEB13D54",
    x"BEB1491E",
    x"BEB154E8",
    x"BEB160B2",
    x"BEB16C7C",
    x"BEB17845",
    x"BEB1840F",
    x"BEB18FD8",
    x"BEB19BA1",
    x"BEB1A76B",
    x"BEB1B334",
    x"BEB1BEFD",
    x"BEB1CAC5",
    x"BEB1D68E",
    x"BEB1E257",
    x"BEB1EE1F",
    x"BEB1F9E8",
    x"BEB205B0",
    x"BEB21178",
    x"BEB21D41",
    x"BEB22909",
    x"BEB234D0",
    x"BEB24098",
    x"BEB24C60",
    x"BEB25827",
    x"BEB263EF",
    x"BEB26FB6",
    x"BEB27B7E",
    x"BEB28745",
    x"BEB2930C",
    x"BEB29ED3",
    x"BEB2AA99",
    x"BEB2B660",
    x"BEB2C227",
    x"BEB2CDED",
    x"BEB2D9B4",
    x"BEB2E57A",
    x"BEB2F140",
    x"BEB2FD06",
    x"BEB308CC",
    x"BEB31492",
    x"BEB32058",
    x"BEB32C1D",
    x"BEB337E3",
    x"BEB343A8",
    x"BEB34F6E",
    x"BEB35B33",
    x"BEB366F8",
    x"BEB372BD",
    x"BEB37E82",
    x"BEB38A47",
    x"BEB3960B",
    x"BEB3A1D0",
    x"BEB3AD94",
    x"BEB3B959",
    x"BEB3C51D",
    x"BEB3D0E1",
    x"BEB3DCA5",
    x"BEB3E869",
    x"BEB3F42D",
    x"BEB3FFF0",
    x"BEB40BB4",
    x"BEB41777",
    x"BEB4233B",
    x"BEB42EFE",
    x"BEB43AC1",
    x"BEB44684",
    x"BEB45247",
    x"BEB45E0A",
    x"BEB469CD",
    x"BEB4758F",
    x"BEB48152",
    x"BEB48D14",
    x"BEB498D6",
    x"BEB4A499",
    x"BEB4B05B",
    x"BEB4BC1D",
    x"BEB4C7DE",
    x"BEB4D3A0",
    x"BEB4DF62",
    x"BEB4EB23",
    x"BEB4F6E5",
    x"BEB502A6",
    x"BEB50E67",
    x"BEB51A28",
    x"BEB525E9",
    x"BEB531AA",
    x"BEB53D6B",
    x"BEB5492B",
    x"BEB554EC",
    x"BEB560AC",
    x"BEB56C6D",
    x"BEB5782D",
    x"BEB583ED",
    x"BEB58FAD",
    x"BEB59B6D",
    x"BEB5A72D",
    x"BEB5B2EC",
    x"BEB5BEAC",
    x"BEB5CA6B",
    x"BEB5D62B",
    x"BEB5E1EA",
    x"BEB5EDA9",
    x"BEB5F968",
    x"BEB60527",
    x"BEB610E6",
    x"BEB61CA4",
    x"BEB62863",
    x"BEB63421",
    x"BEB63FE0",
    x"BEB64B9E",
    x"BEB6575C",
    x"BEB6631A",
    x"BEB66ED8",
    x"BEB67A96",
    x"BEB68653",
    x"BEB69211",
    x"BEB69DCE",
    x"BEB6A98C",
    x"BEB6B549",
    x"BEB6C106",
    x"BEB6CCC3",
    x"BEB6D880",
    x"BEB6E43D",
    x"BEB6EFFA",
    x"BEB6FBB6",
    x"BEB70773",
    x"BEB7132F",
    x"BEB71EEB",
    x"BEB72AA7",
    x"BEB73663",
    x"BEB7421F",
    x"BEB74DDB",
    x"BEB75997",
    x"BEB76552",
    x"BEB7710E",
    x"BEB77CC9",
    x"BEB78884",
    x"BEB79440",
    x"BEB79FFB",
    x"BEB7ABB6",
    x"BEB7B770",
    x"BEB7C32B",
    x"BEB7CEE6",
    x"BEB7DAA0",
    x"BEB7E65B",
    x"BEB7F215",
    x"BEB7FDCF",
    x"BEB80989",
    x"BEB81543",
    x"BEB820FD",
    x"BEB82CB6",
    x"BEB83870",
    x"BEB8442A",
    x"BEB84FE3",
    x"BEB85B9C",
    x"BEB86755",
    x"BEB8730E",
    x"BEB87EC7",
    x"BEB88A80",
    x"BEB89639",
    x"BEB8A1F1",
    x"BEB8ADAA",
    x"BEB8B962",
    x"BEB8C51B",
    x"BEB8D0D3",
    x"BEB8DC8B",
    x"BEB8E843",
    x"BEB8F3FA",
    x"BEB8FFB2",
    x"BEB90B6A",
    x"BEB91721",
    x"BEB922D9",
    x"BEB92E90",
    x"BEB93A47",
    x"BEB945FE",
    x"BEB951B5",
    x"BEB95D6C",
    x"BEB96923",
    x"BEB974D9",
    x"BEB98090",
    x"BEB98C46",
    x"BEB997FC",
    x"BEB9A3B2",
    x"BEB9AF68",
    x"BEB9BB1E",
    x"BEB9C6D4",
    x"BEB9D28A",
    x"BEB9DE3F",
    x"BEB9E9F5",
    x"BEB9F5AA",
    x"BEBA015F",
    x"BEBA0D15",
    x"BEBA18CA",
    x"BEBA247F",
    x"BEBA3033",
    x"BEBA3BE8",
    x"BEBA479D",
    x"BEBA5351",
    x"BEBA5F05",
    x"BEBA6ABA",
    x"BEBA766E",
    x"BEBA8222",
    x"BEBA8DD6",
    x"BEBA9989",
    x"BEBAA53D",
    x"BEBAB0F1",
    x"BEBABCA4",
    x"BEBAC857",
    x"BEBAD40B",
    x"BEBADFBE",
    x"BEBAEB71",
    x"BEBAF724",
    x"BEBB02D6",
    x"BEBB0E89",
    x"BEBB1A3C",
    x"BEBB25EE",
    x"BEBB31A0",
    x"BEBB3D53",
    x"BEBB4905",
    x"BEBB54B7",
    x"BEBB6069",
    x"BEBB6C1A",
    x"BEBB77CC",
    x"BEBB837E",
    x"BEBB8F2F",
    x"BEBB9AE0",
    x"BEBBA692",
    x"BEBBB243",
    x"BEBBBDF4",
    x"BEBBC9A4",
    x"BEBBD555",
    x"BEBBE106",
    x"BEBBECB6",
    x"BEBBF867",
    x"BEBC0417",
    x"BEBC0FC7",
    x"BEBC1B77",
    x"BEBC2727",
    x"BEBC32D7",
    x"BEBC3E87",
    x"BEBC4A36",
    x"BEBC55E6",
    x"BEBC6195",
    x"BEBC6D45",
    x"BEBC78F4",
    x"BEBC84A3",
    x"BEBC9052",
    x"BEBC9C00",
    x"BEBCA7AF",
    x"BEBCB35E",
    x"BEBCBF0C",
    x"BEBCCABB",
    x"BEBCD669",
    x"BEBCE217",
    x"BEBCEDC5",
    x"BEBCF973",
    x"BEBD0521",
    x"BEBD10CE",
    x"BEBD1C7C",
    x"BEBD2829",
    x"BEBD33D7",
    x"BEBD3F84",
    x"BEBD4B31",
    x"BEBD56DE",
    x"BEBD628B",
    x"BEBD6E38",
    x"BEBD79E4",
    x"BEBD8591",
    x"BEBD913D",
    x"BEBD9CEA",
    x"BEBDA896",
    x"BEBDB442",
    x"BEBDBFEE",
    x"BEBDCB9A",
    x"BEBDD746",
    x"BEBDE2F1",
    x"BEBDEE9D",
    x"BEBDFA48",
    x"BEBE05F3",
    x"BEBE119E",
    x"BEBE1D4A",
    x"BEBE28F4",
    x"BEBE349F",
    x"BEBE404A",
    x"BEBE4BF5",
    x"BEBE579F",
    x"BEBE6349",
    x"BEBE6EF4",
    x"BEBE7A9E",
    x"BEBE8648",
    x"BEBE91F2",
    x"BEBE9D9C",
    x"BEBEA945",
    x"BEBEB4EF",
    x"BEBEC098",
    x"BEBECC42",
    x"BEBED7EB",
    x"BEBEE394",
    x"BEBEEF3D",
    x"BEBEFAE6",
    x"BEBF068F",
    x"BEBF1237",
    x"BEBF1DE0",
    x"BEBF2988",
    x"BEBF3530",
    x"BEBF40D9",
    x"BEBF4C81",
    x"BEBF5829",
    x"BEBF63D0",
    x"BEBF6F78",
    x"BEBF7B20",
    x"BEBF86C7",
    x"BEBF926F",
    x"BEBF9E16",
    x"BEBFA9BD",
    x"BEBFB564",
    x"BEBFC10B",
    x"BEBFCCB2",
    x"BEBFD858",
    x"BEBFE3FF",
    x"BEBFEFA5",
    x"BEBFFB4C",
    x"BEC006F2",
    x"BEC01298",
    x"BEC01E3E",
    x"BEC029E4",
    x"BEC0358A",
    x"BEC0412F",
    x"BEC04CD5",
    x"BEC0587A",
    x"BEC06420",
    x"BEC06FC5",
    x"BEC07B6A",
    x"BEC0870F",
    x"BEC092B4",
    x"BEC09E58",
    x"BEC0A9FD",
    x"BEC0B5A1",
    x"BEC0C146",
    x"BEC0CCEA",
    x"BEC0D88E",
    x"BEC0E432",
    x"BEC0EFD6",
    x"BEC0FB7A",
    x"BEC1071E",
    x"BEC112C1",
    x"BEC11E64",
    x"BEC12A08",
    x"BEC135AB",
    x"BEC1414E",
    x"BEC14CF1",
    x"BEC15894",
    x"BEC16437",
    x"BEC16FD9",
    x"BEC17B7C",
    x"BEC1871E",
    x"BEC192C0",
    x"BEC19E63",
    x"BEC1AA05",
    x"BEC1B5A7",
    x"BEC1C148",
    x"BEC1CCEA",
    x"BEC1D88C",
    x"BEC1E42D",
    x"BEC1EFCE",
    x"BEC1FB70",
    x"BEC20711",
    x"BEC212B2",
    x"BEC21E53",
    x"BEC229F3",
    x"BEC23594",
    x"BEC24135",
    x"BEC24CD5",
    x"BEC25875",
    x"BEC26415",
    x"BEC26FB5",
    x"BEC27B55",
    x"BEC286F5",
    x"BEC29295",
    x"BEC29E34",
    x"BEC2A9D4",
    x"BEC2B573",
    x"BEC2C112",
    x"BEC2CCB2",
    x"BEC2D851",
    x"BEC2E3EF",
    x"BEC2EF8E",
    x"BEC2FB2D",
    x"BEC306CB",
    x"BEC3126A",
    x"BEC31E08",
    x"BEC329A6",
    x"BEC33544",
    x"BEC340E2",
    x"BEC34C80",
    x"BEC3581E",
    x"BEC363BB",
    x"BEC36F59",
    x"BEC37AF6",
    x"BEC38693",
    x"BEC39231",
    x"BEC39DCE",
    x"BEC3A96A",
    x"BEC3B507",
    x"BEC3C0A4",
    x"BEC3CC40",
    x"BEC3D7DD",
    x"BEC3E379",
    x"BEC3EF15",
    x"BEC3FAB1",
    x"BEC4064D",
    x"BEC411E9",
    x"BEC41D85",
    x"BEC42920",
    x"BEC434BC",
    x"BEC44057",
    x"BEC44BF2",
    x"BEC4578D",
    x"BEC46328",
    x"BEC46EC3",
    x"BEC47A5E",
    x"BEC485F9",
    x"BEC49193",
    x"BEC49D2E",
    x"BEC4A8C8",
    x"BEC4B462",
    x"BEC4BFFC",
    x"BEC4CB96",
    x"BEC4D730",
    x"BEC4E2C9",
    x"BEC4EE63",
    x"BEC4F9FD",
    x"BEC50596",
    x"BEC5112F",
    x"BEC51CC8",
    x"BEC52861",
    x"BEC533FA",
    x"BEC53F93",
    x"BEC54B2B",
    x"BEC556C4",
    x"BEC5625C",
    x"BEC56DF4",
    x"BEC5798D",
    x"BEC58525",
    x"BEC590BD",
    x"BEC59C54",
    x"BEC5A7EC",
    x"BEC5B384",
    x"BEC5BF1B",
    x"BEC5CAB2",
    x"BEC5D649",
    x"BEC5E1E1",
    x"BEC5ED77",
    x"BEC5F90E",
    x"BEC604A5",
    x"BEC6103C",
    x"BEC61BD2",
    x"BEC62768",
    x"BEC632FF",
    x"BEC63E95",
    x"BEC64A2B",
    x"BEC655C1",
    x"BEC66156",
    x"BEC66CEC",
    x"BEC67882",
    x"BEC68417",
    x"BEC68FAC",
    x"BEC69B41",
    x"BEC6A6D6",
    x"BEC6B26B",
    x"BEC6BE00",
    x"BEC6C995",
    x"BEC6D529",
    x"BEC6E0BE",
    x"BEC6EC52",
    x"BEC6F7E6",
    x"BEC7037B",
    x"BEC70F0E",
    x"BEC71AA2",
    x"BEC72636",
    x"BEC731CA",
    x"BEC73D5D",
    x"BEC748F0",
    x"BEC75484",
    x"BEC76017",
    x"BEC76BAA",
    x"BEC7773D",
    x"BEC782D0",
    x"BEC78E62",
    x"BEC799F5",
    x"BEC7A587",
    x"BEC7B119",
    x"BEC7BCAC",
    x"BEC7C83E",
    x"BEC7D3CF",
    x"BEC7DF61",
    x"BEC7EAF3",
    x"BEC7F685",
    x"BEC80216",
    x"BEC80DA7",
    x"BEC81938",
    x"BEC824CA",
    x"BEC8305B",
    x"BEC83BEB",
    x"BEC8477C",
    x"BEC8530D",
    x"BEC85E9D",
    x"BEC86A2D",
    x"BEC875BE",
    x"BEC8814E",
    x"BEC88CDE",
    x"BEC8986E",
    x"BEC8A3FD",
    x"BEC8AF8D",
    x"BEC8BB1D",
    x"BEC8C6AC",
    x"BEC8D23B",
    x"BEC8DDCA",
    x"BEC8E959",
    x"BEC8F4E8",
    x"BEC90077",
    x"BEC90C06",
    x"BEC91794",
    x"BEC92323",
    x"BEC92EB1",
    x"BEC93A3F",
    x"BEC945CD",
    x"BEC9515B",
    x"BEC95CE9",
    x"BEC96877",
    x"BEC97404",
    x"BEC97F92",
    x"BEC98B1F",
    x"BEC996AC",
    x"BEC9A239",
    x"BEC9ADC6",
    x"BEC9B953",
    x"BEC9C4E0",
    x"BEC9D06C",
    x"BEC9DBF9",
    x"BEC9E785",
    x"BEC9F312",
    x"BEC9FE9E",
    x"BECA0A2A",
    x"BECA15B5",
    x"BECA2141",
    x"BECA2CCD",
    x"BECA3858",
    x"BECA43E4",
    x"BECA4F6F",
    x"BECA5AFA",
    x"BECA6685",
    x"BECA7210",
    x"BECA7D9B",
    x"BECA8925",
    x"BECA94B0",
    x"BECAA03A",
    x"BECAABC5",
    x"BECAB74F",
    x"BECAC2D9",
    x"BECACE63",
    x"BECAD9ED",
    x"BECAE576",
    x"BECAF100",
    x"BECAFC89",
    x"BECB0813",
    x"BECB139C",
    x"BECB1F25",
    x"BECB2AAE",
    x"BECB3637",
    x"BECB41BF",
    x"BECB4D48",
    x"BECB58D0",
    x"BECB6459",
    x"BECB6FE1",
    x"BECB7B69",
    x"BECB86F1",
    x"BECB9279",
    x"BECB9E00",
    x"BECBA988",
    x"BECBB50F",
    x"BECBC097",
    x"BECBCC1E",
    x"BECBD7A5",
    x"BECBE32C",
    x"BECBEEB3",
    x"BECBFA3A",
    x"BECC05C0",
    x"BECC1147",
    x"BECC1CCD",
    x"BECC2853",
    x"BECC33DA",
    x"BECC3F60",
    x"BECC4AE5",
    x"BECC566B",
    x"BECC61F1",
    x"BECC6D76",
    x"BECC78FC",
    x"BECC8481",
    x"BECC9006",
    x"BECC9B8B",
    x"BECCA710",
    x"BECCB295",
    x"BECCBE19",
    x"BECCC99E",
    x"BECCD522",
    x"BECCE0A7",
    x"BECCEC2B",
    x"BECCF7AF",
    x"BECD0333",
    x"BECD0EB6",
    x"BECD1A3A",
    x"BECD25BE",
    x"BECD3141",
    x"BECD3CC4",
    x"BECD4847",
    x"BECD53CA",
    x"BECD5F4D",
    x"BECD6AD0",
    x"BECD7653",
    x"BECD81D5",
    x"BECD8D58",
    x"BECD98DA",
    x"BECDA45C",
    x"BECDAFDE",
    x"BECDBB60",
    x"BECDC6E2",
    x"BECDD264",
    x"BECDDDE5",
    x"BECDE967",
    x"BECDF4E8",
    x"BECE0069",
    x"BECE0BEA",
    x"BECE176B",
    x"BECE22EC",
    x"BECE2E6D",
    x"BECE39ED",
    x"BECE456E",
    x"BECE50EE",
    x"BECE5C6E",
    x"BECE67EE",
    x"BECE736E",
    x"BECE7EEE",
    x"BECE8A6E",
    x"BECE95ED",
    x"BECEA16D",
    x"BECEACEC",
    x"BECEB86B",
    x"BECEC3EA",
    x"BECECF69",
    x"BECEDAE8",
    x"BECEE667",
    x"BECEF1E5",
    x"BECEFD64",
    x"BECF08E2",
    x"BECF1460",
    x"BECF1FDE",
    x"BECF2B5C",
    x"BECF36DA",
    x"BECF4258",
    x"BECF4DD5",
    x"BECF5953",
    x"BECF64D0",
    x"BECF704D",
    x"BECF7BCA",
    x"BECF8747",
    x"BECF92C4",
    x"BECF9E41",
    x"BECFA9BD",
    x"BECFB53A",
    x"BECFC0B6",
    x"BECFCC32",
    x"BECFD7AE",
    x"BECFE32A",
    x"BECFEEA6",
    x"BECFFA22",
    x"BED0059D",
    x"BED01119",
    x"BED01C94",
    x"BED0280F",
    x"BED0338A",
    x"BED03F05",
    x"BED04A80",
    x"BED055FB",
    x"BED06175",
    x"BED06CF0",
    x"BED0786A",
    x"BED083E4",
    x"BED08F5E",
    x"BED09AD8",
    x"BED0A652",
    x"BED0B1CC",
    x"BED0BD45",
    x"BED0C8BF",
    x"BED0D438",
    x"BED0DFB1",
    x"BED0EB2A",
    x"BED0F6A3",
    x"BED1021C",
    x"BED10D95",
    x"BED1190D",
    x"BED12485",
    x"BED12FFE",
    x"BED13B76",
    x"BED146EE",
    x"BED15266",
    x"BED15DDE",
    x"BED16955",
    x"BED174CD",
    x"BED18044",
    x"BED18BBC",
    x"BED19733",
    x"BED1A2AA",
    x"BED1AE21",
    x"BED1B998",
    x"BED1C50E",
    x"BED1D085",
    x"BED1DBFB",
    x"BED1E771",
    x"BED1F2E8",
    x"BED1FE5E",
    x"BED209D3",
    x"BED21549",
    x"BED220BF",
    x"BED22C34",
    x"BED237AA",
    x"BED2431F",
    x"BED24E94",
    x"BED25A09",
    x"BED2657E",
    x"BED270F3",
    x"BED27C68",
    x"BED287DC",
    x"BED29350",
    x"BED29EC5",
    x"BED2AA39",
    x"BED2B5AD",
    x"BED2C121",
    x"BED2CC94",
    x"BED2D808",
    x"BED2E37C",
    x"BED2EEEF",
    x"BED2FA62",
    x"BED305D5",
    x"BED31148",
    x"BED31CBB",
    x"BED3282E",
    x"BED333A0",
    x"BED33F13",
    x"BED34A85",
    x"BED355F7",
    x"BED3616A",
    x"BED36CDB",
    x"BED3784D",
    x"BED383BF",
    x"BED38F31",
    x"BED39AA2",
    x"BED3A613",
    x"BED3B185",
    x"BED3BCF6",
    x"BED3C867",
    x"BED3D3D7",
    x"BED3DF48",
    x"BED3EAB9",
    x"BED3F629",
    x"BED40199",
    x"BED40D0A",
    x"BED4187A",
    x"BED423EA",
    x"BED42F59",
    x"BED43AC9",
    x"BED44639",
    x"BED451A8",
    x"BED45D17",
    x"BED46886",
    x"BED473F5",
    x"BED47F64",
    x"BED48AD3",
    x"BED49642",
    x"BED4A1B0",
    x"BED4AD1F",
    x"BED4B88D",
    x"BED4C3FB",
    x"BED4CF69",
    x"BED4DAD7",
    x"BED4E645",
    x"BED4F1B2",
    x"BED4FD20",
    x"BED5088D",
    x"BED513FA",
    x"BED51F68",
    x"BED52AD5",
    x"BED53641",
    x"BED541AE",
    x"BED54D1B",
    x"BED55887",
    x"BED563F3",
    x"BED56F60",
    x"BED57ACC",
    x"BED58638",
    x"BED591A4",
    x"BED59D0F",
    x"BED5A87B",
    x"BED5B3E6",
    x"BED5BF52",
    x"BED5CABD",
    x"BED5D628",
    x"BED5E193",
    x"BED5ECFD",
    x"BED5F868",
    x"BED603D3",
    x"BED60F3D",
    x"BED61AA7",
    x"BED62611",
    x"BED6317B",
    x"BED63CE5",
    x"BED6484F",
    x"BED653B9",
    x"BED65F22",
    x"BED66A8C",
    x"BED675F5",
    x"BED6815E",
    x"BED68CC7",
    x"BED69830",
    x"BED6A399",
    x"BED6AF01",
    x"BED6BA6A",
    x"BED6C5D2",
    x"BED6D13A",
    x"BED6DCA2",
    x"BED6E80A",
    x"BED6F372",
    x"BED6FEDA",
    x"BED70A41",
    x"BED715A9",
    x"BED72110",
    x"BED72C77",
    x"BED737DE",
    x"BED74345",
    x"BED74EAC",
    x"BED75A13",
    x"BED76579",
    x"BED770E0",
    x"BED77C46",
    x"BED787AC",
    x"BED79312",
    x"BED79E78",
    x"BED7A9DE",
    x"BED7B543",
    x"BED7C0A9",
    x"BED7CC0E",
    x"BED7D773",
    x"BED7E2D8",
    x"BED7EE3D",
    x"BED7F9A2",
    x"BED80507",
    x"BED8106B",
    x"BED81BD0",
    x"BED82734",
    x"BED83298",
    x"BED83DFC",
    x"BED84960",
    x"BED854C4",
    x"BED86028",
    x"BED86B8B",
    x"BED876EF",
    x"BED88252",
    x"BED88DB5",
    x"BED89918",
    x"BED8A47B",
    x"BED8AFDE",
    x"BED8BB40",
    x"BED8C6A3",
    x"BED8D205",
    x"BED8DD67",
    x"BED8E8CA",
    x"BED8F42C",
    x"BED8FF8D",
    x"BED90AEF",
    x"BED91651",
    x"BED921B2",
    x"BED92D13",
    x"BED93875",
    x"BED943D6",
    x"BED94F37",
    x"BED95A97",
    x"BED965F8",
    x"BED97159",
    x"BED97CB9",
    x"BED98819",
    x"BED99379",
    x"BED99ED9",
    x"BED9AA39",
    x"BED9B599",
    x"BED9C0F9",
    x"BED9CC58",
    x"BED9D7B7",
    x"BED9E317",
    x"BED9EE76",
    x"BED9F9D5",
    x"BEDA0533",
    x"BEDA1092",
    x"BEDA1BF1",
    x"BEDA274F",
    x"BEDA32AD",
    x"BEDA3E0C",
    x"BEDA496A",
    x"BEDA54C8",
    x"BEDA6025",
    x"BEDA6B83",
    x"BEDA76E0",
    x"BEDA823E",
    x"BEDA8D9B",
    x"BEDA98F8",
    x"BEDAA455",
    x"BEDAAFB2",
    x"BEDABB0F",
    x"BEDAC66B",
    x"BEDAD1C8",
    x"BEDADD24",
    x"BEDAE880",
    x"BEDAF3DC",
    x"BEDAFF38",
    x"BEDB0A94",
    x"BEDB15F0",
    x"BEDB214B",
    x"BEDB2CA7",
    x"BEDB3802",
    x"BEDB435D",
    x"BEDB4EB8",
    x"BEDB5A13",
    x"BEDB656E",
    x"BEDB70C8",
    x"BEDB7C23",
    x"BEDB877D",
    x"BEDB92D7",
    x"BEDB9E31",
    x"BEDBA98B",
    x"BEDBB4E5",
    x"BEDBC03F",
    x"BEDBCB98",
    x"BEDBD6F2",
    x"BEDBE24B",
    x"BEDBEDA4",
    x"BEDBF8FD",
    x"BEDC0456",
    x"BEDC0FAF",
    x"BEDC1B08",
    x"BEDC2660",
    x"BEDC31B8",
    x"BEDC3D11",
    x"BEDC4869",
    x"BEDC53C1",
    x"BEDC5F18",
    x"BEDC6A70",
    x"BEDC75C8",
    x"BEDC811F",
    x"BEDC8C76",
    x"BEDC97CE",
    x"BEDCA325",
    x"BEDCAE7C",
    x"BEDCB9D2",
    x"BEDCC529",
    x"BEDCD07F",
    x"BEDCDBD6",
    x"BEDCE72C",
    x"BEDCF282",
    x"BEDCFDD8",
    x"BEDD092E",
    x"BEDD1484",
    x"BEDD1FD9",
    x"BEDD2B2F",
    x"BEDD3684",
    x"BEDD41D9",
    x"BEDD4D2E",
    x"BEDD5883",
    x"BEDD63D8",
    x"BEDD6F2C",
    x"BEDD7A81",
    x"BEDD85D5",
    x"BEDD912A",
    x"BEDD9C7E",
    x"BEDDA7D2",
    x"BEDDB325",
    x"BEDDBE79",
    x"BEDDC9CD",
    x"BEDDD520",
    x"BEDDE073",
    x"BEDDEBC7",
    x"BEDDF71A",
    x"BEDE026C",
    x"BEDE0DBF",
    x"BEDE1912",
    x"BEDE2464",
    x"BEDE2FB7",
    x"BEDE3B09",
    x"BEDE465B",
    x"BEDE51AD",
    x"BEDE5CFF",
    x"BEDE6851",
    x"BEDE73A2",
    x"BEDE7EF3",
    x"BEDE8A45",
    x"BEDE9596",
    x"BEDEA0E7",
    x"BEDEAC38",
    x"BEDEB789",
    x"BEDEC2D9",
    x"BEDECE2A",
    x"BEDED97A",
    x"BEDEE4CA",
    x"BEDEF01A",
    x"BEDEFB6A",
    x"BEDF06BA",
    x"BEDF120A",
    x"BEDF1D59",
    x"BEDF28A9",
    x"BEDF33F8",
    x"BEDF3F47",
    x"BEDF4A96",
    x"BEDF55E5",
    x"BEDF6134",
    x"BEDF6C82",
    x"BEDF77D1",
    x"BEDF831F",
    x"BEDF8E6D",
    x"BEDF99BB",
    x"BEDFA509",
    x"BEDFB057",
    x"BEDFBBA5",
    x"BEDFC6F2",
    x"BEDFD240",
    x"BEDFDD8D",
    x"BEDFE8DA",
    x"BEDFF427",
    x"BEDFFF74",
    x"BEE00AC1",
    x"BEE0160D",
    x"BEE0215A",
    x"BEE02CA6",
    x"BEE037F2",
    x"BEE0433E",
    x"BEE04E8A",
    x"BEE059D6",
    x"BEE06522",
    x"BEE0706D",
    x"BEE07BB8",
    x"BEE08704",
    x"BEE0924F",
    x"BEE09D9A",
    x"BEE0A8E5",
    x"BEE0B42F",
    x"BEE0BF7A",
    x"BEE0CAC4",
    x"BEE0D60E",
    x"BEE0E159",
    x"BEE0ECA3",
    x"BEE0F7ED",
    x"BEE10336",
    x"BEE10E80",
    x"BEE119C9",
    x"BEE12513",
    x"BEE1305C",
    x"BEE13BA5",
    x"BEE146EE",
    x"BEE15237",
    x"BEE15D7F",
    x"BEE168C8",
    x"BEE17410",
    x"BEE17F58",
    x"BEE18AA1",
    x"BEE195E9",
    x"BEE1A130",
    x"BEE1AC78",
    x"BEE1B7C0",
    x"BEE1C307",
    x"BEE1CE4E",
    x"BEE1D996",
    x"BEE1E4DD",
    x"BEE1F023",
    x"BEE1FB6A",
    x"BEE206B1",
    x"BEE211F7",
    x"BEE21D3E",
    x"BEE22884",
    x"BEE233CA",
    x"BEE23F10",
    x"BEE24A56",
    x"BEE2559B",
    x"BEE260E1",
    x"BEE26C26",
    x"BEE2776C",
    x"BEE282B1",
    x"BEE28DF6",
    x"BEE2993A",
    x"BEE2A47F",
    x"BEE2AFC4",
    x"BEE2BB08",
    x"BEE2C64C",
    x"BEE2D191",
    x"BEE2DCD5",
    x"BEE2E819",
    x"BEE2F35C",
    x"BEE2FEA0",
    x"BEE309E3",
    x"BEE31527",
    x"BEE3206A",
    x"BEE32BAD",
    x"BEE336F0",
    x"BEE34233",
    x"BEE34D75",
    x"BEE358B8",
    x"BEE363FA",
    x"BEE36F3D",
    x"BEE37A7F",
    x"BEE385C1",
    x"BEE39102",
    x"BEE39C44",
    x"BEE3A786",
    x"BEE3B2C7",
    x"BEE3BE08",
    x"BEE3C94A",
    x"BEE3D48B",
    x"BEE3DFCB",
    x"BEE3EB0C",
    x"BEE3F64D",
    x"BEE4018D",
    x"BEE40CCE",
    x"BEE4180E",
    x"BEE4234E",
    x"BEE42E8E",
    x"BEE439CE",
    x"BEE4450D",
    x"BEE4504D",
    x"BEE45B8C",
    x"BEE466CB",
    x"BEE4720A",
    x"BEE47D49",
    x"BEE48888",
    x"BEE493C7",
    x"BEE49F05",
    x"BEE4AA44",
    x"BEE4B582",
    x"BEE4C0C0",
    x"BEE4CBFE",
    x"BEE4D73C",
    x"BEE4E27A",
    x"BEE4EDB7",
    x"BEE4F8F5",
    x"BEE50432",
    x"BEE50F6F",
    x"BEE51AAC",
    x"BEE525E9",
    x"BEE53126",
    x"BEE53C62",
    x"BEE5479F",
    x"BEE552DB",
    x"BEE55E17",
    x"BEE56953",
    x"BEE5748F",
    x"BEE57FCB",
    x"BEE58B07",
    x"BEE59642",
    x"BEE5A17E",
    x"BEE5ACB9",
    x"BEE5B7F4",
    x"BEE5C32F",
    x"BEE5CE6A",
    x"BEE5D9A4",
    x"BEE5E4DF",
    x"BEE5F019",
    x"BEE5FB54",
    x"BEE6068E",
    x"BEE611C8",
    x"BEE61D02",
    x"BEE6283B",
    x"BEE63375",
    x"BEE63EAE",
    x"BEE649E7",
    x"BEE65521",
    x"BEE6605A",
    x"BEE66B93",
    x"BEE676CB",
    x"BEE68204",
    x"BEE68D3C",
    x"BEE69875",
    x"BEE6A3AD",
    x"BEE6AEE5",
    x"BEE6BA1D",
    x"BEE6C554",
    x"BEE6D08C",
    x"BEE6DBC4",
    x"BEE6E6FB",
    x"BEE6F232",
    x"BEE6FD69",
    x"BEE708A0",
    x"BEE713D7",
    x"BEE71F0E",
    x"BEE72A44",
    x"BEE7357A",
    x"BEE740B1",
    x"BEE74BE7",
    x"BEE7571D",
    x"BEE76253",
    x"BEE76D88",
    x"BEE778BE",
    x"BEE783F3",
    x"BEE78F28",
    x"BEE79A5D",
    x"BEE7A592",
    x"BEE7B0C7",
    x"BEE7BBFC",
    x"BEE7C731",
    x"BEE7D265",
    x"BEE7DD99",
    x"BEE7E8CD",
    x"BEE7F401",
    x"BEE7FF35",
    x"BEE80A69",
    x"BEE8159C",
    x"BEE820D0",
    x"BEE82C03",
    x"BEE83736",
    x"BEE84269",
    x"BEE84D9C",
    x"BEE858CF",
    x"BEE86402",
    x"BEE86F34",
    x"BEE87A66",
    x"BEE88599",
    x"BEE890CB",
    x"BEE89BFD",
    x"BEE8A72E",
    x"BEE8B260",
    x"BEE8BD91",
    x"BEE8C8C3",
    x"BEE8D3F4",
    x"BEE8DF25",
    x"BEE8EA56",
    x"BEE8F587",
    x"BEE900B7",
    x"BEE90BE8",
    x"BEE91718",
    x"BEE92248",
    x"BEE92D78",
    x"BEE938A8",
    x"BEE943D8",
    x"BEE94F08",
    x"BEE95A37",
    x"BEE96567",
    x"BEE97096",
    x"BEE97BC5",
    x"BEE986F4",
    x"BEE99223",
    x"BEE99D51",
    x"BEE9A880",
    x"BEE9B3AE",
    x"BEE9BEDD",
    x"BEE9CA0B",
    x"BEE9D539",
    x"BEE9E066",
    x"BEE9EB94",
    x"BEE9F6C2",
    x"BEEA01EF",
    x"BEEA0D1C",
    x"BEEA1849",
    x"BEEA2376",
    x"BEEA2EA3",
    x"BEEA39D0",
    x"BEEA44FD",
    x"BEEA5029",
    x"BEEA5B55",
    x"BEEA6681",
    x"BEEA71AD",
    x"BEEA7CD9",
    x"BEEA8805",
    x"BEEA9330",
    x"BEEA9E5C",
    x"BEEAA987",
    x"BEEAB4B2",
    x"BEEABFDD",
    x"BEEACB08",
    x"BEEAD633",
    x"BEEAE15D",
    x"BEEAEC88",
    x"BEEAF7B2",
    x"BEEB02DC",
    x"BEEB0E06",
    x"BEEB1930",
    x"BEEB245A",
    x"BEEB2F84",
    x"BEEB3AAD",
    x"BEEB45D6",
    x"BEEB50FF",
    x"BEEB5C28",
    x"BEEB6751",
    x"BEEB727A",
    x"BEEB7DA3",
    x"BEEB88CB",
    x"BEEB93F3",
    x"BEEB9F1C",
    x"BEEBAA44",
    x"BEEBB56C",
    x"BEEBC093",
    x"BEEBCBBB",
    x"BEEBD6E2",
    x"BEEBE20A",
    x"BEEBED31",
    x"BEEBF858",
    x"BEEC037F",
    x"BEEC0EA5",
    x"BEEC19CC",
    x"BEEC24F3",
    x"BEEC3019",
    x"BEEC3B3F",
    x"BEEC4665",
    x"BEEC518B",
    x"BEEC5CB1",
    x"BEEC67D6",
    x"BEEC72FC",
    x"BEEC7E21",
    x"BEEC8946",
    x"BEEC946B",
    x"BEEC9F90",
    x"BEECAAB5",
    x"BEECB5DA",
    x"BEECC0FE",
    x"BEECCC22",
    x"BEECD747",
    x"BEECE26B",
    x"BEECED8F",
    x"BEECF8B2",
    x"BEED03D6",
    x"BEED0EF9",
    x"BEED1A1D",
    x"BEED2540",
    x"BEED3063",
    x"BEED3B86",
    x"BEED46A9",
    x"BEED51CB",
    x"BEED5CEE",
    x"BEED6810",
    x"BEED7332",
    x"BEED7E54",
    x"BEED8976",
    x"BEED9498",
    x"BEED9FB9",
    x"BEEDAADB",
    x"BEEDB5FC",
    x"BEEDC11D",
    x"BEEDCC3E",
    x"BEEDD75F",
    x"BEEDE280",
    x"BEEDEDA1",
    x"BEEDF8C1",
    x"BEEE03E2",
    x"BEEE0F02",
    x"BEEE1A22",
    x"BEEE2542",
    x"BEEE3061",
    x"BEEE3B81",
    x"BEEE46A0",
    x"BEEE51C0",
    x"BEEE5CDF",
    x"BEEE67FE",
    x"BEEE731D",
    x"BEEE7E3C",
    x"BEEE895A",
    x"BEEE9479",
    x"BEEE9F97",
    x"BEEEAAB5",
    x"BEEEB5D3",
    x"BEEEC0F1",
    x"BEEECC0F",
    x"BEEED72C",
    x"BEEEE24A",
    x"BEEEED67",
    x"BEEEF884",
    x"BEEF03A1",
    x"BEEF0EBE",
    x"BEEF19DB",
    x"BEEF24F7",
    x"BEEF3014",
    x"BEEF3B30",
    x"BEEF464C",
    x"BEEF5168",
    x"BEEF5C84",
    x"BEEF67A0",
    x"BEEF72BC",
    x"BEEF7DD7",
    x"BEEF88F2",
    x"BEEF940D",
    x"BEEF9F28",
    x"BEEFAA43",
    x"BEEFB55E",
    x"BEEFC079",
    x"BEEFCB93",
    x"BEEFD6AD",
    x"BEEFE1C7",
    x"BEEFECE1",
    x"BEEFF7FB",
    x"BEF00315",
    x"BEF00E2E",
    x"BEF01948",
    x"BEF02461",
    x"BEF02F7A",
    x"BEF03A93",
    x"BEF045AC",
    x"BEF050C5",
    x"BEF05BDD",
    x"BEF066F6",
    x"BEF0720E",
    x"BEF07D26",
    x"BEF0883E",
    x"BEF09356",
    x"BEF09E6E",
    x"BEF0A985",
    x"BEF0B49C",
    x"BEF0BFB4",
    x"BEF0CACB",
    x"BEF0D5E2",
    x"BEF0E0F9",
    x"BEF0EC0F",
    x"BEF0F726",
    x"BEF1023C",
    x"BEF10D52",
    x"BEF11868",
    x"BEF1237E",
    x"BEF12E94",
    x"BEF139AA",
    x"BEF144BF",
    x"BEF14FD5",
    x"BEF15AEA",
    x"BEF165FF",
    x"BEF17114",
    x"BEF17C28",
    x"BEF1873D",
    x"BEF19252",
    x"BEF19D66",
    x"BEF1A87A",
    x"BEF1B38E",
    x"BEF1BEA2",
    x"BEF1C9B6",
    x"BEF1D4C9",
    x"BEF1DFDD",
    x"BEF1EAF0",
    x"BEF1F603",
    x"BEF20116",
    x"BEF20C29",
    x"BEF2173C",
    x"BEF2224F",
    x"BEF22D61",
    x"BEF23873",
    x"BEF24385",
    x"BEF24E97",
    x"BEF259A9",
    x"BEF264BB",
    x"BEF26FCD",
    x"BEF27ADE",
    x"BEF285EF",
    x"BEF29100",
    x"BEF29C11",
    x"BEF2A722",
    x"BEF2B233",
    x"BEF2BD43",
    x"BEF2C854",
    x"BEF2D364",
    x"BEF2DE74",
    x"BEF2E984",
    x"BEF2F494",
    x"BEF2FFA4",
    x"BEF30AB3",
    x"BEF315C2",
    x"BEF320D2",
    x"BEF32BE1",
    x"BEF336F0",
    x"BEF341FE",
    x"BEF34D0D",
    x"BEF3581C",
    x"BEF3632A",
    x"BEF36E38",
    x"BEF37946",
    x"BEF38454",
    x"BEF38F62",
    x"BEF39A6F",
    x"BEF3A57D",
    x"BEF3B08A",
    x"BEF3BB97",
    x"BEF3C6A4",
    x"BEF3D1B1",
    x"BEF3DCBE",
    x"BEF3E7CB",
    x"BEF3F2D7",
    x"BEF3FDE3",
    x"BEF408F0",
    x"BEF413FB",
    x"BEF41F07",
    x"BEF42A13",
    x"BEF4351F",
    x"BEF4402A",
    x"BEF44B35",
    x"BEF45640",
    x"BEF4614B",
    x"BEF46C56",
    x"BEF47761",
    x"BEF4826B",
    x"BEF48D76",
    x"BEF49880",
    x"BEF4A38A",
    x"BEF4AE94",
    x"BEF4B99E",
    x"BEF4C4A7",
    x"BEF4CFB1",
    x"BEF4DABA",
    x"BEF4E5C3",
    x"BEF4F0CC",
    x"BEF4FBD5",
    x"BEF506DE",
    x"BEF511E7",
    x"BEF51CEF",
    x"BEF527F8",
    x"BEF53300",
    x"BEF53E08",
    x"BEF54910",
    x"BEF55417",
    x"BEF55F1F",
    x"BEF56A26",
    x"BEF5752E",
    x"BEF58035",
    x"BEF58B3C",
    x"BEF59643",
    x"BEF5A149",
    x"BEF5AC50",
    x"BEF5B756",
    x"BEF5C25C",
    x"BEF5CD62",
    x"BEF5D868",
    x"BEF5E36E",
    x"BEF5EE74",
    x"BEF5F979",
    x"BEF6047F",
    x"BEF60F84",
    x"BEF61A89",
    x"BEF6258E",
    x"BEF63093",
    x"BEF63B97",
    x"BEF6469C",
    x"BEF651A0",
    x"BEF65CA4",
    x"BEF667A8",
    x"BEF672AC",
    x"BEF67DB0",
    x"BEF688B3",
    x"BEF693B7",
    x"BEF69EBA",
    x"BEF6A9BD",
    x"BEF6B4C0",
    x"BEF6BFC3",
    x"BEF6CAC6",
    x"BEF6D5C8",
    x"BEF6E0CB",
    x"BEF6EBCD",
    x"BEF6F6CF",
    x"BEF701D1",
    x"BEF70CD3",
    x"BEF717D4",
    x"BEF722D6",
    x"BEF72DD7",
    x"BEF738D8",
    x"BEF743D9",
    x"BEF74EDA",
    x"BEF759DB",
    x"BEF764DC",
    x"BEF76FDC",
    x"BEF77ADC",
    x"BEF785DC",
    x"BEF790DC",
    x"BEF79BDC",
    x"BEF7A6DC",
    x"BEF7B1DC",
    x"BEF7BCDB",
    x"BEF7C7DA",
    x"BEF7D2D9",
    x"BEF7DDD8",
    x"BEF7E8D7",
    x"BEF7F3D6",
    x"BEF7FED4",
    x"BEF809D3",
    x"BEF814D1",
    x"BEF81FCF",
    x"BEF82ACD",
    x"BEF835CB",
    x"BEF840C8",
    x"BEF84BC6",
    x"BEF856C3",
    x"BEF861C0",
    x"BEF86CBD",
    x"BEF877BA",
    x"BEF882B7",
    x"BEF88DB3",
    x"BEF898B0",
    x"BEF8A3AC",
    x"BEF8AEA8",
    x"BEF8B9A4",
    x"BEF8C4A0",
    x"BEF8CF9C",
    x"BEF8DA97",
    x"BEF8E592",
    x"BEF8F08E",
    x"BEF8FB89",
    x"BEF90684",
    x"BEF9117E",
    x"BEF91C79",
    x"BEF92773",
    x"BEF9326E",
    x"BEF93D68",
    x"BEF94862",
    x"BEF9535C",
    x"BEF95E56",
    x"BEF9694F",
    x"BEF97449",
    x"BEF97F42",
    x"BEF98A3B",
    x"BEF99534",
    x"BEF9A02D",
    x"BEF9AB25",
    x"BEF9B61E",
    x"BEF9C116",
    x"BEF9CC0E",
    x"BEF9D707",
    x"BEF9E1FE",
    x"BEF9ECF6",
    x"BEF9F7EE",
    x"BEFA02E5",
    x"BEFA0DDD",
    x"BEFA18D4",
    x"BEFA23CB",
    x"BEFA2EC2",
    x"BEFA39B8",
    x"BEFA44AF",
    x"BEFA4FA5",
    x"BEFA5A9C",
    x"BEFA6592",
    x"BEFA7088",
    x"BEFA7B7D",
    x"BEFA8673",
    x"BEFA9169",
    x"BEFA9C5E",
    x"BEFAA753",
    x"BEFAB248",
    x"BEFABD3D",
    x"BEFAC832",
    x"BEFAD326",
    x"BEFADE1B",
    x"BEFAE90F",
    x"BEFAF403",
    x"BEFAFEF7",
    x"BEFB09EB",
    x"BEFB14DF",
    x"BEFB1FD2",
    x"BEFB2AC6",
    x"BEFB35B9",
    x"BEFB40AC",
    x"BEFB4B9F",
    x"BEFB5692",
    x"BEFB6184",
    x"BEFB6C77",
    x"BEFB7769",
    x"BEFB825B",
    x"BEFB8D4D",
    x"BEFB983F",
    x"BEFBA331",
    x"BEFBAE22",
    x"BEFBB914",
    x"BEFBC405",
    x"BEFBCEF6",
    x"BEFBD9E7",
    x"BEFBE4D8",
    x"BEFBEFC9",
    x"BEFBFAB9",
    x"BEFC05AA",
    x"BEFC109A",
    x"BEFC1B8A",
    x"BEFC267A",
    x"BEFC3169",
    x"BEFC3C59",
    x"BEFC4748",
    x"BEFC5238",
    x"BEFC5D27",
    x"BEFC6816",
    x"BEFC7305",
    x"BEFC7DF3",
    x"BEFC88E2",
    x"BEFC93D0",
    x"BEFC9EBF",
    x"BEFCA9AD",
    x"BEFCB49B",
    x"BEFCBF88",
    x"BEFCCA76",
    x"BEFCD563",
    x"BEFCE051",
    x"BEFCEB3E",
    x"BEFCF62B",
    x"BEFD0118",
    x"BEFD0C04",
    x"BEFD16F1",
    x"BEFD21DD",
    x"BEFD2CCA",
    x"BEFD37B6",
    x"BEFD42A2",
    x"BEFD4D8D",
    x"BEFD5879",
    x"BEFD6365",
    x"BEFD6E50",
    x"BEFD793B",
    x"BEFD8426",
    x"BEFD8F11",
    x"BEFD99FC",
    x"BEFDA4E6",
    x"BEFDAFD1",
    x"BEFDBABB",
    x"BEFDC5A5",
    x"BEFDD08F",
    x"BEFDDB79",
    x"BEFDE662",
    x"BEFDF14C",
    x"BEFDFC35",
    x"BEFE071E",
    x"BEFE1207",
    x"BEFE1CF0",
    x"BEFE27D9",
    x"BEFE32C2",
    x"BEFE3DAA",
    x"BEFE4892",
    x"BEFE537A",
    x"BEFE5E62",
    x"BEFE694A",
    x"BEFE7432",
    x"BEFE7F19",
    x"BEFE8A01",
    x"BEFE94E8",
    x"BEFE9FCF",
    x"BEFEAAB6",
    x"BEFEB59D",
    x"BEFEC083",
    x"BEFECB6A",
    x"BEFED650",
    x"BEFEE136",
    x"BEFEEC1C",
    x"BEFEF702",
    x"BEFF01E8",
    x"BEFF0CCD",
    x"BEFF17B2",
    x"BEFF2298",
    x"BEFF2D7D",
    x"BEFF3862",
    x"BEFF4346",
    x"BEFF4E2B",
    x"BEFF590F",
    x"BEFF63F4",
    x"BEFF6ED8",
    x"BEFF79BC",
    x"BEFF849F",
    x"BEFF8F83",
    x"BEFF9A67",
    x"BEFFA54A",
    x"BEFFB02D",
    x"BEFFBB10",
    x"BEFFC5F3",
    x"BEFFD0D6",
    x"BEFFDBB8",
    x"BEFFE69B",
    x"BEFFF17D",
    x"BEFFFC5F",
    x"BF0003A1",
    x"BF000912",
    x"BF000E82",
    x"BF0013F3",
    x"BF001964",
    x"BF001ED4",
    x"BF002445",
    x"BF0029B5",
    x"BF002F26",
    x"BF003496",
    x"BF003A06",
    x"BF003F76",
    x"BF0044E6",
    x"BF004A56",
    x"BF004FC6",
    x"BF005536",
    x"BF005AA6",
    x"BF006016",
    x"BF006585",
    x"BF006AF5",
    x"BF007064",
    x"BF0075D4",
    x"BF007B43",
    x"BF0080B2",
    x"BF008621",
    x"BF008B90",
    x"BF0090FF",
    x"BF00966E",
    x"BF009BDD",
    x"BF00A14C",
    x"BF00A6BA",
    x"BF00AC29",
    x"BF00B197",
    x"BF00B706",
    x"BF00BC74",
    x"BF00C1E2",
    x"BF00C751",
    x"BF00CCBF",
    x"BF00D22D",
    x"BF00D79B",
    x"BF00DD09",
    x"BF00E276",
    x"BF00E7E4",
    x"BF00ED52",
    x"BF00F2BF",
    x"BF00F82D",
    x"BF00FD9A",
    x"BF010308",
    x"BF010875",
    x"BF010DE2",
    x"BF01134F",
    x"BF0118BC",
    x"BF011E29",
    x"BF012396",
    x"BF012903",
    x"BF012E70",
    x"BF0133DC",
    x"BF013949",
    x"BF013EB5",
    x"BF014422",
    x"BF01498E",
    x"BF014EFA",
    x"BF015467",
    x"BF0159D3",
    x"BF015F3F",
    x"BF0164AB",
    x"BF016A17",
    x"BF016F82",
    x"BF0174EE",
    x"BF017A5A",
    x"BF017FC5",
    x"BF018531",
    x"BF018A9C",
    x"BF019007",
    x"BF019573",
    x"BF019ADE",
    x"BF01A049",
    x"BF01A5B4",
    x"BF01AB1F",
    x"BF01B08A",
    x"BF01B5F5",
    x"BF01BB5F",
    x"BF01C0CA",
    x"BF01C634",
    x"BF01CB9F",
    x"BF01D109",
    x"BF01D674",
    x"BF01DBDE",
    x"BF01E148",
    x"BF01E6B2",
    x"BF01EC1C",
    x"BF01F186",
    x"BF01F6F0",
    x"BF01FC59",
    x"BF0201C3",
    x"BF02072D",
    x"BF020C96",
    x"BF021200",
    x"BF021769",
    x"BF021CD2",
    x"BF02223C",
    x"BF0227A5",
    x"BF022D0E",
    x"BF023277",
    x"BF0237E0",
    x"BF023D48",
    x"BF0242B1",
    x"BF02481A",
    x"BF024D82",
    x"BF0252EB",
    x"BF025853",
    x"BF025DBC",
    x"BF026324",
    x"BF02688C",
    x"BF026DF4",
    x"BF02735C",
    x"BF0278C4",
    x"BF027E2C",
    x"BF028394",
    x"BF0288FC",
    x"BF028E63",
    x"BF0293CB",
    x"BF029932",
    x"BF029E9A",
    x"BF02A401",
    x"BF02A968",
    x"BF02AED0",
    x"BF02B437",
    x"BF02B99E",
    x"BF02BF05",
    x"BF02C46B",
    x"BF02C9D2",
    x"BF02CF39",
    x"BF02D49F",
    x"BF02DA06",
    x"BF02DF6C",
    x"BF02E4D3",
    x"BF02EA39",
    x"BF02EF9F",
    x"BF02F506",
    x"BF02FA6C",
    x"BF02FFD2",
    x"BF030537",
    x"BF030A9D",
    x"BF031003",
    x"BF031569",
    x"BF031ACE",
    x"BF032034",
    x"BF032599",
    x"BF032AFF",
    x"BF033064",
    x"BF0335C9",
    x"BF033B2E",
    x"BF034093",
    x"BF0345F8",
    x"BF034B5D",
    x"BF0350C2",
    x"BF035627",
    x"BF035B8B",
    x"BF0360F0",
    x"BF036654",
    x"BF036BB9",
    x"BF03711D",
    x"BF037681",
    x"BF037BE5",
    x"BF03814A",
    x"BF0386AE",
    x"BF038C11",
    x"BF039175",
    x"BF0396D9",
    x"BF039C3D",
    x"BF03A1A0",
    x"BF03A704",
    x"BF03AC67",
    x"BF03B1CB",
    x"BF03B72E",
    x"BF03BC91",
    x"BF03C1F4",
    x"BF03C757",
    x"BF03CCBA",
    x"BF03D21D",
    x"BF03D780",
    x"BF03DCE3",
    x"BF03E246",
    x"BF03E7A8",
    x"BF03ED0B",
    x"BF03F26D",
    x"BF03F7CF",
    x"BF03FD32",
    x"BF040294",
    x"BF0407F6",
    x"BF040D58",
    x"BF0412BA",
    x"BF04181C",
    x"BF041D7E",
    x"BF0422DF",
    x"BF042841",
    x"BF042DA2",
    x"BF043304",
    x"BF043865",
    x"BF043DC7",
    x"BF044328",
    x"BF044889",
    x"BF044DEA",
    x"BF04534B",
    x"BF0458AC",
    x"BF045E0D",
    x"BF04636E",
    x"BF0468CE",
    x"BF046E2F",
    x"BF04738F",
    x"BF0478F0",
    x"BF047E50",
    x"BF0483B0",
    x"BF048911",
    x"BF048E71",
    x"BF0493D1",
    x"BF049931",
    x"BF049E91",
    x"BF04A3F0",
    x"BF04A950",
    x"BF04AEB0",
    x"BF04B40F",
    x"BF04B96F",
    x"BF04BECE",
    x"BF04C42D",
    x"BF04C98D",
    x"BF04CEEC",
    x"BF04D44B",
    x"BF04D9AA",
    x"BF04DF09",
    x"BF04E468",
    x"BF04E9C6",
    x"BF04EF25",
    x"BF04F484",
    x"BF04F9E2",
    x"BF04FF41",
    x"BF05049F",
    x"BF0509FD",
    x"BF050F5B",
    x"BF0514BA",
    x"BF051A18",
    x"BF051F75",
    x"BF0524D3",
    x"BF052A31",
    x"BF052F8F",
    x"BF0534EC",
    x"BF053A4A",
    x"BF053FA8",
    x"BF054505",
    x"BF054A62",
    x"BF054FBF",
    x"BF05551D",
    x"BF055A7A",
    x"BF055FD7",
    x"BF056534",
    x"BF056A90",
    x"BF056FED",
    x"BF05754A",
    x"BF057AA6",
    x"BF058003",
    x"BF05855F",
    x"BF058ABC",
    x"BF059018",
    x"BF059574",
    x"BF059AD0",
    x"BF05A02C",
    x"BF05A588",
    x"BF05AAE4",
    x"BF05B040",
    x"BF05B59C",
    x"BF05BAF7",
    x"BF05C053",
    x"BF05C5AE",
    x"BF05CB0A",
    x"BF05D065",
    x"BF05D5C0",
    x"BF05DB1B",
    x"BF05E076",
    x"BF05E5D1",
    x"BF05EB2C",
    x"BF05F087",
    x"BF05F5E2",
    x"BF05FB3C",
    x"BF060097",
    x"BF0605F1",
    x"BF060B4C",
    x"BF0610A6",
    x"BF061600",
    x"BF061B5B",
    x"BF0620B5",
    x"BF06260F",
    x"BF062B69",
    x"BF0630C2",
    x"BF06361C",
    x"BF063B76",
    x"BF0640CF",
    x"BF064629",
    x"BF064B82",
    x"BF0650DC",
    x"BF065635",
    x"BF065B8E",
    x"BF0660E7",
    x"BF066640",
    x"BF066B99",
    x"BF0670F2",
    x"BF06764B",
    x"BF067BA4",
    x"BF0680FC",
    x"BF068655",
    x"BF068BAD",
    x"BF069106",
    x"BF06965E",
    x"BF069BB6",
    x"BF06A10E",
    x"BF06A667",
    x"BF06ABBF",
    x"BF06B116",
    x"BF06B66E",
    x"BF06BBC6",
    x"BF06C11E",
    x"BF06C675",
    x"BF06CBCD",
    x"BF06D124",
    x"BF06D67B",
    x"BF06DBD3",
    x"BF06E12A",
    x"BF06E681",
    x"BF06EBD8",
    x"BF06F12F",
    x"BF06F686",
    x"BF06FBDD",
    x"BF070133",
    x"BF07068A",
    x"BF070BE0",
    x"BF071137",
    x"BF07168D",
    x"BF071BE3",
    x"BF07213A",
    x"BF072690",
    x"BF072BE6",
    x"BF07313C",
    x"BF073692",
    x"BF073BE7",
    x"BF07413D",
    x"BF074693",
    x"BF074BE8",
    x"BF07513E",
    x"BF075693",
    x"BF075BE8",
    x"BF07613E",
    x"BF076693",
    x"BF076BE8",
    x"BF07713D",
    x"BF077692",
    x"BF077BE6",
    x"BF07813B",
    x"BF078690",
    x"BF078BE4",
    x"BF079139",
    x"BF07968D",
    x"BF079BE2",
    x"BF07A136",
    x"BF07A68A",
    x"BF07ABDE",
    x"BF07B132",
    x"BF07B686",
    x"BF07BBDA",
    x"BF07C12E",
    x"BF07C681",
    x"BF07CBD5",
    x"BF07D128",
    x"BF07D67C",
    x"BF07DBCF",
    x"BF07E122",
    x"BF07E676",
    x"BF07EBC9",
    x"BF07F11C",
    x"BF07F66F",
    x"BF07FBC1",
    x"BF080114",
    x"BF080667",
    x"BF080BB9",
    x"BF08110C",
    x"BF08165E",
    x"BF081BB1",
    x"BF082103",
    x"BF082655",
    x"BF082BA7",
    x"BF0830F9",
    x"BF08364B",
    x"BF083B9D",
    x"BF0840EF",
    x"BF084641",
    x"BF084B92",
    x"BF0850E4",
    x"BF085635",
    x"BF085B87",
    x"BF0860D8",
    x"BF086629",
    x"BF086B7A",
    x"BF0870CB",
    x"BF08761C",
    x"BF087B6D",
    x"BF0880BE",
    x"BF08860F",
    x"BF088B5F",
    x"BF0890B0",
    x"BF089600",
    x"BF089B51",
    x"BF08A0A1",
    x"BF08A5F1",
    x"BF08AB41",
    x"BF08B091",
    x"BF08B5E1",
    x"BF08BB31",
    x"BF08C081",
    x"BF08C5D1",
    x"BF08CB20",
    x"BF08D070",
    x"BF08D5BF",
    x"BF08DB0F",
    x"BF08E05E",
    x"BF08E5AD",
    x"BF08EAFD",
    x"BF08F04C",
    x"BF08F59B",
    x"BF08FAEA",
    x"BF090038",
    x"BF090587",
    x"BF090AD6",
    x"BF091024",
    x"BF091573",
    x"BF091AC1",
    x"BF092010",
    x"BF09255E",
    x"BF092AAC",
    x"BF092FFA",
    x"BF093548",
    x"BF093A96",
    x"BF093FE4",
    x"BF094531",
    x"BF094A7F",
    x"BF094FCD",
    x"BF09551A",
    x"BF095A68",
    x"BF095FB5",
    x"BF096502",
    x"BF096A4F",
    x"BF096F9C",
    x"BF0974E9",
    x"BF097A36",
    x"BF097F83",
    x"BF0984D0",
    x"BF098A1D",
    x"BF098F69",
    x"BF0994B6",
    x"BF099A02",
    x"BF099F4E",
    x"BF09A49B",
    x"BF09A9E7",
    x"BF09AF33",
    x"BF09B47F",
    x"BF09B9CB",
    x"BF09BF17",
    x"BF09C463",
    x"BF09C9AE",
    x"BF09CEFA",
    x"BF09D445",
    x"BF09D991",
    x"BF09DEDC",
    x"BF09E427",
    x"BF09E973",
    x"BF09EEBE",
    x"BF09F409",
    x"BF09F954",
    x"BF09FE9E",
    x"BF0A03E9",
    x"BF0A0934",
    x"BF0A0E7E",
    x"BF0A13C9",
    x"BF0A1913",
    x"BF0A1E5E",
    x"BF0A23A8",
    x"BF0A28F2",
    x"BF0A2E3C",
    x"BF0A3386",
    x"BF0A38D0",
    x"BF0A3E1A",
    x"BF0A4364",
    x"BF0A48AD",
    x"BF0A4DF7",
    x"BF0A5341",
    x"BF0A588A",
    x"BF0A5DD3",
    x"BF0A631D",
    x"BF0A6866",
    x"BF0A6DAF",
    x"BF0A72F8",
    x"BF0A7841",
    x"BF0A7D8A",
    x"BF0A82D2",
    x"BF0A881B",
    x"BF0A8D64",
    x"BF0A92AC",
    x"BF0A97F5",
    x"BF0A9D3D",
    x"BF0AA285",
    x"BF0AA7CD",
    x"BF0AAD16",
    x"BF0AB25E",
    x"BF0AB7A5",
    x"BF0ABCED",
    x"BF0AC235",
    x"BF0AC77D",
    x"BF0ACCC4",
    x"BF0AD20C",
    x"BF0AD753",
    x"BF0ADC9B",
    x"BF0AE1E2",
    x"BF0AE729",
    x"BF0AEC70",
    x"BF0AF1B7",
    x"BF0AF6FE",
    x"BF0AFC45",
    x"BF0B018C",
    x"BF0B06D2",
    x"BF0B0C19",
    x"BF0B115F",
    x"BF0B16A6",
    x"BF0B1BEC",
    x"BF0B2132",
    x"BF0B2679",
    x"BF0B2BBF",
    x"BF0B3105",
    x"BF0B364B",
    x"BF0B3B90",
    x"BF0B40D6",
    x"BF0B461C",
    x"BF0B4B61",
    x"BF0B50A7",
    x"BF0B55EC",
    x"BF0B5B32",
    x"BF0B6077",
    x"BF0B65BC",
    x"BF0B6B01",
    x"BF0B7046",
    x"BF0B758B",
    x"BF0B7AD0",
    x"BF0B8015",
    x"BF0B8559",
    x"BF0B8A9E",
    x"BF0B8FE2",
    x"BF0B9527",
    x"BF0B9A6B",
    x"BF0B9FAF",
    x"BF0BA4F4",
    x"BF0BAA38",
    x"BF0BAF7C",
    x"BF0BB4BF",
    x"BF0BBA03",
    x"BF0BBF47",
    x"BF0BC48B",
    x"BF0BC9CE",
    x"BF0BCF12",
    x"BF0BD455",
    x"BF0BD998",
    x"BF0BDEDC",
    x"BF0BE41F",
    x"BF0BE962",
    x"BF0BEEA5",
    x"BF0BF3E8",
    x"BF0BF92B",
    x"BF0BFE6D",
    x"BF0C03B0",
    x"BF0C08F2",
    x"BF0C0E35",
    x"BF0C1377",
    x"BF0C18BA",
    x"BF0C1DFC",
    x"BF0C233E",
    x"BF0C2880",
    x"BF0C2DC2",
    x"BF0C3304",
    x"BF0C3846",
    x"BF0C3D87",
    x"BF0C42C9",
    x"BF0C480B",
    x"BF0C4D4C",
    x"BF0C528D",
    x"BF0C57CF",
    x"BF0C5D10",
    x"BF0C6251",
    x"BF0C6792",
    x"BF0C6CD3",
    x"BF0C7214",
    x"BF0C7755",
    x"BF0C7C95",
    x"BF0C81D6",
    x"BF0C8716",
    x"BF0C8C57",
    x"BF0C9197",
    x"BF0C96D7",
    x"BF0C9C18",
    x"BF0CA158",
    x"BF0CA698",
    x"BF0CABD8",
    x"BF0CB118",
    x"BF0CB657",
    x"BF0CBB97",
    x"BF0CC0D7",
    x"BF0CC616",
    x"BF0CCB56",
    x"BF0CD095",
    x"BF0CD5D4",
    x"BF0CDB13",
    x"BF0CE052",
    x"BF0CE591",
    x"BF0CEAD0",
    x"BF0CF00F",
    x"BF0CF54E",
    x"BF0CFA8D",
    x"BF0CFFCB",
    x"BF0D050A",
    x"BF0D0A48",
    x"BF0D0F86",
    x"BF0D14C5",
    x"BF0D1A03",
    x"BF0D1F41",
    x"BF0D247F",
    x"BF0D29BD",
    x"BF0D2EFA",
    x"BF0D3438",
    x"BF0D3976",
    x"BF0D3EB3",
    x"BF0D43F1",
    x"BF0D492E",
    x"BF0D4E6C",
    x"BF0D53A9",
    x"BF0D58E6",
    x"BF0D5E23",
    x"BF0D6360",
    x"BF0D689D",
    x"BF0D6DDA",
    x"BF0D7316",
    x"BF0D7853",
    x"BF0D7D8F",
    x"BF0D82CC",
    x"BF0D8808",
    x"BF0D8D45",
    x"BF0D9281",
    x"BF0D97BD",
    x"BF0D9CF9",
    x"BF0DA235",
    x"BF0DA771",
    x"BF0DACAC",
    x"BF0DB1E8",
    x"BF0DB724",
    x"BF0DBC5F",
    x"BF0DC19B",
    x"BF0DC6D6",
    x"BF0DCC11",
    x"BF0DD14C",
    x"BF0DD687",
    x"BF0DDBC2",
    x"BF0DE0FD",
    x"BF0DE638",
    x"BF0DEB73",
    x"BF0DF0AE",
    x"BF0DF5E8",
    x"BF0DFB23",
    x"BF0E005D",
    x"BF0E0597",
    x"BF0E0AD2",
    x"BF0E100C",
    x"BF0E1546",
    x"BF0E1A80",
    x"BF0E1FBA",
    x"BF0E24F3",
    x"BF0E2A2D",
    x"BF0E2F67",
    x"BF0E34A0",
    x"BF0E39DA",
    x"BF0E3F13",
    x"BF0E444C",
    x"BF0E4986",
    x"BF0E4EBF",
    x"BF0E53F8",
    x"BF0E5931",
    x"BF0E5E6A",
    x"BF0E63A2",
    x"BF0E68DB",
    x"BF0E6E14",
    x"BF0E734C",
    x"BF0E7885",
    x"BF0E7DBD",
    x"BF0E82F5",
    x"BF0E882D",
    x"BF0E8D65",
    x"BF0E929D",
    x"BF0E97D5",
    x"BF0E9D0D",
    x"BF0EA245",
    x"BF0EA77D",
    x"BF0EACB4",
    x"BF0EB1EC",
    x"BF0EB723",
    x"BF0EBC5A",
    x"BF0EC192",
    x"BF0EC6C9",
    x"BF0ECC00",
    x"BF0ED137",
    x"BF0ED66E",
    x"BF0EDBA4",
    x"BF0EE0DB",
    x"BF0EE612",
    x"BF0EEB48",
    x"BF0EF07F",
    x"BF0EF5B5",
    x"BF0EFAEB",
    x"BF0F0022",
    x"BF0F0558",
    x"BF0F0A8E",
    x"BF0F0FC4",
    x"BF0F14FA",
    x"BF0F1A2F",
    x"BF0F1F65",
    x"BF0F249B",
    x"BF0F29D0",
    x"BF0F2F05",
    x"BF0F343B",
    x"BF0F3970",
    x"BF0F3EA5",
    x"BF0F43DA",
    x"BF0F490F",
    x"BF0F4E44",
    x"BF0F5379",
    x"BF0F58AE",
    x"BF0F5DE2",
    x"BF0F6317",
    x"BF0F684B",
    x"BF0F6D80",
    x"BF0F72B4",
    x"BF0F77E8",
    x"BF0F7D1C",
    x"BF0F8250",
    x"BF0F8784",
    x"BF0F8CB8",
    x"BF0F91EC",
    x"BF0F9720",
    x"BF0F9C53",
    x"BF0FA187",
    x"BF0FA6BA",
    x"BF0FABEE",
    x"BF0FB121",
    x"BF0FB654",
    x"BF0FBB87",
    x"BF0FC0BA",
    x"BF0FC5ED",
    x"BF0FCB20",
    x"BF0FD053",
    x"BF0FD585",
    x"BF0FDAB8",
    x"BF0FDFEA",
    x"BF0FE51D",
    x"BF0FEA4F",
    x"BF0FEF81",
    x"BF0FF4B3",
    x"BF0FF9E5",
    x"BF0FFF17",
    x"BF100449",
    x"BF10097B",
    x"BF100EAD",
    x"BF1013DE",
    x"BF101910",
    x"BF101E41",
    x"BF102373",
    x"BF1028A4",
    x"BF102DD5",
    x"BF103306",
    x"BF103837",
    x"BF103D68",
    x"BF104299",
    x"BF1047CA",
    x"BF104CFA",
    x"BF10522B",
    x"BF10575B",
    x"BF105C8C",
    x"BF1061BC",
    x"BF1066EC",
    x"BF106C1C",
    x"BF10714C",
    x"BF10767C",
    x"BF107BAC",
    x"BF1080DC",
    x"BF10860C",
    x"BF108B3B",
    x"BF10906B",
    x"BF10959A",
    x"BF109ACA",
    x"BF109FF9",
    x"BF10A528",
    x"BF10AA57",
    x"BF10AF86",
    x"BF10B4B5",
    x"BF10B9E4",
    x"BF10BF13",
    x"BF10C441",
    x"BF10C970",
    x"BF10CE9E",
    x"BF10D3CD",
    x"BF10D8FB",
    x"BF10DE29",
    x"BF10E357",
    x"BF10E885",
    x"BF10EDB3",
    x"BF10F2E1",
    x"BF10F80F",
    x"BF10FD3D",
    x"BF11026A",
    x"BF110798",
    x"BF110CC5",
    x"BF1111F3",
    x"BF111720",
    x"BF111C4D",
    x"BF11217A",
    x"BF1126A7",
    x"BF112BD4",
    x"BF113101",
    x"BF11362E",
    x"BF113B5A",
    x"BF114087",
    x"BF1145B3",
    x"BF114AE0",
    x"BF11500C",
    x"BF115538",
    x"BF115A64",
    x"BF115F90",
    x"BF1164BC",
    x"BF1169E8",
    x"BF116F14",
    x"BF117440",
    x"BF11796B",
    x"BF117E97",
    x"BF1183C2",
    x"BF1188ED",
    x"BF118E19",
    x"BF119344",
    x"BF11986F",
    x"BF119D9A",
    x"BF11A2C5",
    x"BF11A7F0",
    x"BF11AD1A",
    x"BF11B245",
    x"BF11B76F",
    x"BF11BC9A",
    x"BF11C1C4",
    x"BF11C6EF",
    x"BF11CC19",
    x"BF11D143",
    x"BF11D66D",
    x"BF11DB97",
    x"BF11E0C1",
    x"BF11E5EA",
    x"BF11EB14",
    x"BF11F03E",
    x"BF11F567",
    x"BF11FA91",
    x"BF11FFBA",
    x"BF1204E3",
    x"BF120A0C",
    x"BF120F35",
    x"BF12145E",
    x"BF121987",
    x"BF121EB0",
    x"BF1223D9",
    x"BF122901",
    x"BF122E2A",
    x"BF123352",
    x"BF12387A",
    x"BF123DA3",
    x"BF1242CB",
    x"BF1247F3",
    x"BF124D1B",
    x"BF125243",
    x"BF12576B",
    x"BF125C92",
    x"BF1261BA",
    x"BF1266E2",
    x"BF126C09",
    x"BF127130",
    x"BF127658",
    x"BF127B7F",
    x"BF1280A6",
    x"BF1285CD",
    x"BF128AF4",
    x"BF12901B",
    x"BF129542",
    x"BF129A68",
    x"BF129F8F",
    x"BF12A4B5",
    x"BF12A9DC",
    x"BF12AF02",
    x"BF12B428",
    x"BF12B94E",
    x"BF12BE74",
    x"BF12C39A",
    x"BF12C8C0",
    x"BF12CDE6",
    x"BF12D30C",
    x"BF12D831",
    x"BF12DD57",
    x"BF12E27C",
    x"BF12E7A2",
    x"BF12ECC7",
    x"BF12F1EC",
    x"BF12F711",
    x"BF12FC36",
    x"BF13015B",
    x"BF130680",
    x"BF130BA5",
    x"BF1310C9",
    x"BF1315EE",
    x"BF131B12",
    x"BF132037",
    x"BF13255B",
    x"BF132A7F",
    x"BF132FA3",
    x"BF1334C7",
    x"BF1339EB",
    x"BF133F0F",
    x"BF134433",
    x"BF134956",
    x"BF134E7A",
    x"BF13539D",
    x"BF1358C1",
    x"BF135DE4",
    x"BF136307",
    x"BF13682A",
    x"BF136D4D",
    x"BF137270",
    x"BF137793",
    x"BF137CB6",
    x"BF1381D9",
    x"BF1386FB",
    x"BF138C1E",
    x"BF139140",
    x"BF139663",
    x"BF139B85",
    x"BF13A0A7",
    x"BF13A5C9",
    x"BF13AAEB",
    x"BF13B00D",
    x"BF13B52F",
    x"BF13BA50",
    x"BF13BF72",
    x"BF13C493",
    x"BF13C9B5",
    x"BF13CED6",
    x"BF13D3F8",
    x"BF13D919",
    x"BF13DE3A",
    x"BF13E35B",
    x"BF13E87C",
    x"BF13ED9C",
    x"BF13F2BD",
    x"BF13F7DE",
    x"BF13FCFE",
    x"BF14021F",
    x"BF14073F",
    x"BF140C5F",
    x"BF141180",
    x"BF1416A0",
    x"BF141BC0",
    x"BF1420E0",
    x"BF142600",
    x"BF142B1F",
    x"BF14303F",
    x"BF14355E",
    x"BF143A7E",
    x"BF143F9D",
    x"BF1444BD",
    x"BF1449DC",
    x"BF144EFB",
    x"BF14541A",
    x"BF145939",
    x"BF145E58",
    x"BF146377",
    x"BF146895",
    x"BF146DB4",
    x"BF1472D2",
    x"BF1477F1",
    x"BF147D0F",
    x"BF14822D",
    x"BF14874B",
    x"BF148C69",
    x"BF149187",
    x"BF1496A5",
    x"BF149BC3",
    x"BF14A0E1",
    x"BF14A5FE",
    x"BF14AB1C",
    x"BF14B039",
    x"BF14B557",
    x"BF14BA74",
    x"BF14BF91",
    x"BF14C4AE",
    x"BF14C9CB",
    x"BF14CEE8",
    x"BF14D405",
    x"BF14D921",
    x"BF14DE3E",
    x"BF14E35A",
    x"BF14E877",
    x"BF14ED93",
    x"BF14F2B0",
    x"BF14F7CC",
    x"BF14FCE8",
    x"BF150204",
    x"BF150720",
    x"BF150C3B",
    x"BF151157",
    x"BF151673",
    x"BF151B8E",
    x"BF1520AA",
    x"BF1525C5",
    x"BF152AE0",
    x"BF152FFC",
    x"BF153517",
    x"BF153A32",
    x"BF153F4D",
    x"BF154467",
    x"BF154982",
    x"BF154E9D",
    x"BF1553B7",
    x"BF1558D2",
    x"BF155DEC",
    x"BF156306",
    x"BF156821",
    x"BF156D3B",
    x"BF157255",
    x"BF15776F",
    x"BF157C88",
    x"BF1581A2",
    x"BF1586BC",
    x"BF158BD5",
    x"BF1590EF",
    x"BF159608",
    x"BF159B21",
    x"BF15A03B",
    x"BF15A554",
    x"BF15AA6D",
    x"BF15AF86",
    x"BF15B49F",
    x"BF15B9B7",
    x"BF15BED0",
    x"BF15C3E9",
    x"BF15C901",
    x"BF15CE19",
    x"BF15D332",
    x"BF15D84A",
    x"BF15DD62",
    x"BF15E27A",
    x"BF15E792",
    x"BF15ECAA",
    x"BF15F1C2",
    x"BF15F6D9",
    x"BF15FBF1",
    x"BF160108",
    x"BF160620",
    x"BF160B37",
    x"BF16104E",
    x"BF161565",
    x"BF161A7C",
    x"BF161F93",
    x"BF1624AA",
    x"BF1629C1",
    x"BF162ED8",
    x"BF1633EE",
    x"BF163905",
    x"BF163E1B",
    x"BF164331",
    x"BF164847",
    x"BF164D5E",
    x"BF165274",
    x"BF16578A",
    x"BF165C9F",
    x"BF1661B5",
    x"BF1666CB",
    x"BF166BE0",
    x"BF1670F6",
    x"BF16760B",
    x"BF167B21",
    x"BF168036",
    x"BF16854B",
    x"BF168A60",
    x"BF168F75",
    x"BF16948A",
    x"BF16999F",
    x"BF169EB3",
    x"BF16A3C8",
    x"BF16A8DC",
    x"BF16ADF1",
    x"BF16B305",
    x"BF16B819",
    x"BF16BD2D",
    x"BF16C241",
    x"BF16C755",
    x"BF16CC69",
    x"BF16D17D",
    x"BF16D691",
    x"BF16DBA4",
    x"BF16E0B8",
    x"BF16E5CB",
    x"BF16EADE",
    x"BF16EFF2",
    x"BF16F505",
    x"BF16FA18",
    x"BF16FF2B",
    x"BF17043E",
    x"BF170950",
    x"BF170E63",
    x"BF171376",
    x"BF171888",
    x"BF171D9B",
    x"BF1722AD",
    x"BF1727BF",
    x"BF172CD1",
    x"BF1731E3",
    x"BF1736F5",
    x"BF173C07",
    x"BF174119",
    x"BF17462B",
    x"BF174B3C",
    x"BF17504E",
    x"BF17555F",
    x"BF175A70",
    x"BF175F82",
    x"BF176493",
    x"BF1769A4",
    x"BF176EB5",
    x"BF1773C6",
    x"BF1778D6",
    x"BF177DE7",
    x"BF1782F8",
    x"BF178808",
    x"BF178D18",
    x"BF179229",
    x"BF179739",
    x"BF179C49",
    x"BF17A159",
    x"BF17A669",
    x"BF17AB79",
    x"BF17B089",
    x"BF17B598",
    x"BF17BAA8",
    x"BF17BFB7",
    x"BF17C4C7",
    x"BF17C9D6",
    x"BF17CEE5",
    x"BF17D3F4",
    x"BF17D903",
    x"BF17DE12",
    x"BF17E321",
    x"BF17E830",
    x"BF17ED3F",
    x"BF17F24D",
    x"BF17F75C",
    x"BF17FC6A",
    x"BF180178",
    x"BF180687",
    x"BF180B95",
    x"BF1810A3",
    x"BF1815B1",
    x"BF181ABE",
    x"BF181FCC",
    x"BF1824DA",
    x"BF1829E7",
    x"BF182EF5",
    x"BF183402",
    x"BF183910",
    x"BF183E1D",
    x"BF18432A",
    x"BF184837",
    x"BF184D44",
    x"BF185251",
    x"BF18575D",
    x"BF185C6A",
    x"BF186177",
    x"BF186683",
    x"BF186B8F",
    x"BF18709C",
    x"BF1875A8",
    x"BF187AB4",
    x"BF187FC0",
    x"BF1884CC",
    x"BF1889D8",
    x"BF188EE3",
    x"BF1893EF",
    x"BF1898FB",
    x"BF189E06",
    x"BF18A311",
    x"BF18A81D",
    x"BF18AD28",
    x"BF18B233",
    x"BF18B73E",
    x"BF18BC49",
    x"BF18C154",
    x"BF18C65E",
    x"BF18CB69",
    x"BF18D073",
    x"BF18D57E",
    x"BF18DA88",
    x"BF18DF92",
    x"BF18E49D",
    x"BF18E9A7",
    x"BF18EEB1",
    x"BF18F3BB",
    x"BF18F8C4",
    x"BF18FDCE",
    x"BF1902D8",
    x"BF1907E1",
    x"BF190CEB",
    x"BF1911F4",
    x"BF1916FD",
    x"BF191C06",
    x"BF19210F",
    x"BF192618",
    x"BF192B21",
    x"BF19302A",
    x"BF193533",
    x"BF193A3B",
    x"BF193F44",
    x"BF19444C",
    x"BF194955",
    x"BF194E5D",
    x"BF195365",
    x"BF19586D",
    x"BF195D75",
    x"BF19627D",
    x"BF196784",
    x"BF196C8C",
    x"BF197194",
    x"BF19769B",
    x"BF197BA3",
    x"BF1980AA",
    x"BF1985B1",
    x"BF198AB8",
    x"BF198FBF",
    x"BF1994C6",
    x"BF1999CD",
    x"BF199ED4",
    x"BF19A3DA",
    x"BF19A8E1",
    x"BF19ADE7",
    x"BF19B2EE",
    x"BF19B7F4",
    x"BF19BCFA",
    x"BF19C200",
    x"BF19C706",
    x"BF19CC0C",
    x"BF19D112",
    x"BF19D618",
    x"BF19DB1E",
    x"BF19E023",
    x"BF19E529",
    x"BF19EA2E",
    x"BF19EF33",
    x"BF19F438",
    x"BF19F93D",
    x"BF19FE42",
    x"BF1A0347",
    x"BF1A084C",
    x"BF1A0D51",
    x"BF1A1255",
    x"BF1A175A",
    x"BF1A1C5E",
    x"BF1A2163",
    x"BF1A2667",
    x"BF1A2B6B",
    x"BF1A306F",
    x"BF1A3573",
    x"BF1A3A77",
    x"BF1A3F7B",
    x"BF1A447E",
    x"BF1A4982",
    x"BF1A4E86",
    x"BF1A5389",
    x"BF1A588C",
    x"BF1A5D8F",
    x"BF1A6293",
    x"BF1A6796",
    x"BF1A6C99",
    x"BF1A719B",
    x"BF1A769E",
    x"BF1A7BA1",
    x"BF1A80A3",
    x"BF1A85A6",
    x"BF1A8AA8",
    x"BF1A8FAB",
    x"BF1A94AD",
    x"BF1A99AF",
    x"BF1A9EB1",
    x"BF1AA3B3",
    x"BF1AA8B5",
    x"BF1AADB6",
    x"BF1AB2B8",
    x"BF1AB7BA",
    x"BF1ABCBB",
    x"BF1AC1BC",
    x"BF1AC6BE",
    x"BF1ACBBF",
    x"BF1AD0C0",
    x"BF1AD5C1",
    x"BF1ADAC2",
    x"BF1ADFC3",
    x"BF1AE4C3",
    x"BF1AE9C4",
    x"BF1AEEC4",
    x"BF1AF3C5",
    x"BF1AF8C5",
    x"BF1AFDC5",
    x"BF1B02C6",
    x"BF1B07C6",
    x"BF1B0CC6",
    x"BF1B11C5",
    x"BF1B16C5",
    x"BF1B1BC5",
    x"BF1B20C4",
    x"BF1B25C4",
    x"BF1B2AC3",
    x"BF1B2FC3",
    x"BF1B34C2",
    x"BF1B39C1",
    x"BF1B3EC0",
    x"BF1B43BF",
    x"BF1B48BE",
    x"BF1B4DBD",
    x"BF1B52BB",
    x"BF1B57BA",
    x"BF1B5CB8",
    x"BF1B61B7",
    x"BF1B66B5",
    x"BF1B6BB3",
    x"BF1B70B1",
    x"BF1B75AF",
    x"BF1B7AAD",
    x"BF1B7FAB",
    x"BF1B84A9",
    x"BF1B89A6",
    x"BF1B8EA4",
    x"BF1B93A1",
    x"BF1B989E",
    x"BF1B9D9C",
    x"BF1BA299",
    x"BF1BA796",
    x"BF1BAC93",
    x"BF1BB190",
    x"BF1BB68D",
    x"BF1BBB89",
    x"BF1BC086",
    x"BF1BC582",
    x"BF1BCA7F",
    x"BF1BCF7B",
    x"BF1BD477",
    x"BF1BD973",
    x"BF1BDE6F",
    x"BF1BE36B",
    x"BF1BE867",
    x"BF1BED63",
    x"BF1BF25F",
    x"BF1BF75A",
    x"BF1BFC56",
    x"BF1C0151",
    x"BF1C064C",
    x"BF1C0B47",
    x"BF1C1042",
    x"BF1C153D",
    x"BF1C1A38",
    x"BF1C1F33",
    x"BF1C242E",
    x"BF1C2929",
    x"BF1C2E23",
    x"BF1C331D",
    x"BF1C3818",
    x"BF1C3D12",
    x"BF1C420C",
    x"BF1C4706",
    x"BF1C4C00",
    x"BF1C50FA",
    x"BF1C55F4",
    x"BF1C5AEE",
    x"BF1C5FE7",
    x"BF1C64E1",
    x"BF1C69DA",
    x"BF1C6ED3",
    x"BF1C73CC",
    x"BF1C78C6",
    x"BF1C7DBF",
    x"BF1C82B8",
    x"BF1C87B0",
    x"BF1C8CA9",
    x"BF1C91A2",
    x"BF1C969A",
    x"BF1C9B93",
    x"BF1CA08B",
    x"BF1CA583",
    x"BF1CAA7C",
    x"BF1CAF74",
    x"BF1CB46C",
    x"BF1CB963",
    x"BF1CBE5B",
    x"BF1CC353",
    x"BF1CC84B",
    x"BF1CCD42",
    x"BF1CD239",
    x"BF1CD731",
    x"BF1CDC28",
    x"BF1CE11F",
    x"BF1CE616",
    x"BF1CEB0D",
    x"BF1CF004",
    x"BF1CF4FB",
    x"BF1CF9F1",
    x"BF1CFEE8",
    x"BF1D03DE",
    x"BF1D08D5",
    x"BF1D0DCB",
    x"BF1D12C1",
    x"BF1D17B7",
    x"BF1D1CAD",
    x"BF1D21A3",
    x"BF1D2699",
    x"BF1D2B8F",
    x"BF1D3084",
    x"BF1D357A",
    x"BF1D3A6F",
    x"BF1D3F65",
    x"BF1D445A",
    x"BF1D494F",
    x"BF1D4E44",
    x"BF1D5339",
    x"BF1D582E",
    x"BF1D5D23",
    x"BF1D6217",
    x"BF1D670C",
    x"BF1D6C00",
    x"BF1D70F5",
    x"BF1D75E9",
    x"BF1D7ADD",
    x"BF1D7FD1",
    x"BF1D84C5",
    x"BF1D89B9",
    x"BF1D8EAD",
    x"BF1D93A1",
    x"BF1D9894",
    x"BF1D9D88",
    x"BF1DA27B",
    x"BF1DA76F",
    x"BF1DAC62",
    x"BF1DB155",
    x"BF1DB648",
    x"BF1DBB3B",
    x"BF1DC02E",
    x"BF1DC521",
    x"BF1DCA13",
    x"BF1DCF06",
    x"BF1DD3F8",
    x"BF1DD8EB",
    x"BF1DDDDD",
    x"BF1DE2CF",
    x"BF1DE7C1",
    x"BF1DECB3",
    x"BF1DF1A5",
    x"BF1DF697",
    x"BF1DFB89",
    x"BF1E007B",
    x"BF1E056C",
    x"BF1E0A5D",
    x"BF1E0F4F",
    x"BF1E1440",
    x"BF1E1931",
    x"BF1E1E22",
    x"BF1E2313",
    x"BF1E2804",
    x"BF1E2CF5",
    x"BF1E31E6",
    x"BF1E36D6",
    x"BF1E3BC7",
    x"BF1E40B7",
    x"BF1E45A7",
    x"BF1E4A98",
    x"BF1E4F88",
    x"BF1E5478",
    x"BF1E5968",
    x"BF1E5E57",
    x"BF1E6347",
    x"BF1E6837",
    x"BF1E6D26",
    x"BF1E7216",
    x"BF1E7705",
    x"BF1E7BF4",
    x"BF1E80E3",
    x"BF1E85D2",
    x"BF1E8AC1",
    x"BF1E8FB0",
    x"BF1E949F",
    x"BF1E998E",
    x"BF1E9E7C",
    x"BF1EA36B",
    x"BF1EA859",
    x"BF1EAD47",
    x"BF1EB236",
    x"BF1EB724",
    x"BF1EBC12",
    x"BF1EC100",
    x"BF1EC5ED",
    x"BF1ECADB",
    x"BF1ECFC9",
    x"BF1ED4B6",
    x"BF1ED9A4",
    x"BF1EDE91",
    x"BF1EE37E",
    x"BF1EE86C",
    x"BF1EED59",
    x"BF1EF245",
    x"BF1EF732",
    x"BF1EFC1F",
    x"BF1F010C",
    x"BF1F05F8",
    x"BF1F0AE5",
    x"BF1F0FD1",
    x"BF1F14BD",
    x"BF1F19AA",
    x"BF1F1E96",
    x"BF1F2382",
    x"BF1F286E",
    x"BF1F2D59",
    x"BF1F3245",
    x"BF1F3731",
    x"BF1F3C1C",
    x"BF1F4108",
    x"BF1F45F3",
    x"BF1F4ADE",
    x"BF1F4FC9",
    x"BF1F54B4",
    x"BF1F599F",
    x"BF1F5E8A",
    x"BF1F6375",
    x"BF1F6860",
    x"BF1F6D4A",
    x"BF1F7235",
    x"BF1F771F",
    x"BF1F7C09",
    x"BF1F80F3",
    x"BF1F85DD",
    x"BF1F8AC7",
    x"BF1F8FB1",
    x"BF1F949B",
    x"BF1F9985",
    x"BF1F9E6E",
    x"BF1FA358",
    x"BF1FA841",
    x"BF1FAD2B",
    x"BF1FB214",
    x"BF1FB6FD",
    x"BF1FBBE6",
    x"BF1FC0CF",
    x"BF1FC5B8",
    x"BF1FCAA0",
    x"BF1FCF89",
    x"BF1FD472",
    x"BF1FD95A",
    x"BF1FDE42",
    x"BF1FE32B",
    x"BF1FE813",
    x"BF1FECFB",
    x"BF1FF1E3",
    x"BF1FF6CB",
    x"BF1FFBB2",
    x"BF20009A",
    x"BF200582",
    x"BF200A69",
    x"BF200F50",
    x"BF201438",
    x"BF20191F",
    x"BF201E06",
    x"BF2022ED",
    x"BF2027D4",
    x"BF202CBB",
    x"BF2031A1",
    x"BF203688",
    x"BF203B6F",
    x"BF204055",
    x"BF20453B",
    x"BF204A21",
    x"BF204F08",
    x"BF2053EE",
    x"BF2058D4",
    x"BF205DB9",
    x"BF20629F",
    x"BF206785",
    x"BF206C6A",
    x"BF207150",
    x"BF207635",
    x"BF207B1A",
    x"BF208000",
    x"BF2084E5",
    x"BF2089CA",
    x"BF208EAE",
    x"BF209393",
    x"BF209878",
    x"BF209D5C",
    x"BF20A241",
    x"BF20A725",
    x"BF20AC0A",
    x"BF20B0EE",
    x"BF20B5D2",
    x"BF20BAB6",
    x"BF20BF9A",
    x"BF20C47E",
    x"BF20C961",
    x"BF20CE45",
    x"BF20D328",
    x"BF20D80C",
    x"BF20DCEF",
    x"BF20E1D2",
    x"BF20E6B5",
    x"BF20EB99",
    x"BF20F07B",
    x"BF20F55E",
    x"BF20FA41",
    x"BF20FF24",
    x"BF210406",
    x"BF2108E9",
    x"BF210DCB",
    x"BF2112AD",
    x"BF21178F",
    x"BF211C71",
    x"BF212153",
    x"BF212635",
    x"BF212B17",
    x"BF212FF9",
    x"BF2134DA",
    x"BF2139BC",
    x"BF213E9D",
    x"BF21437E",
    x"BF214860",
    x"BF214D41",
    x"BF215222",
    x"BF215703",
    x"BF215BE3",
    x"BF2160C4",
    x"BF2165A5",
    x"BF216A85",
    x"BF216F66",
    x"BF217446",
    x"BF217926",
    x"BF217E06",
    x"BF2182E6",
    x"BF2187C6",
    x"BF218CA6",
    x"BF219186",
    x"BF219665",
    x"BF219B45",
    x"BF21A024",
    x"BF21A504",
    x"BF21A9E3",
    x"BF21AEC2",
    x"BF21B3A1",
    x"BF21B880",
    x"BF21BD5F",
    x"BF21C23E",
    x"BF21C71C",
    x"BF21CBFB",
    x"BF21D0D9",
    x"BF21D5B8",
    x"BF21DA96",
    x"BF21DF74",
    x"BF21E452",
    x"BF21E930",
    x"BF21EE0E",
    x"BF21F2EC",
    x"BF21F7C9",
    x"BF21FCA7",
    x"BF220185",
    x"BF220662",
    x"BF220B3F",
    x"BF22101C",
    x"BF2214FA",
    x"BF2219D7",
    x"BF221EB3",
    x"BF222390",
    x"BF22286D",
    x"BF222D4A",
    x"BF223226",
    x"BF223702",
    x"BF223BDF",
    x"BF2240BB",
    x"BF224597",
    x"BF224A73",
    x"BF224F4F",
    x"BF22542B",
    x"BF225907",
    x"BF225DE2",
    x"BF2262BE",
    x"BF226799",
    x"BF226C74",
    x"BF227150",
    x"BF22762B",
    x"BF227B06",
    x"BF227FE1",
    x"BF2284BC",
    x"BF228996",
    x"BF228E71",
    x"BF22934C",
    x"BF229826",
    x"BF229D00",
    x"BF22A1DB",
    x"BF22A6B5",
    x"BF22AB8F",
    x"BF22B069",
    x"BF22B543",
    x"BF22BA1D",
    x"BF22BEF6",
    x"BF22C3D0",
    x"BF22C8A9",
    x"BF22CD83",
    x"BF22D25C",
    x"BF22D735",
    x"BF22DC0E",
    x"BF22E0E7",
    x"BF22E5C0",
    x"BF22EA99",
    x"BF22EF72",
    x"BF22F44A",
    x"BF22F923",
    x"BF22FDFB",
    x"BF2302D3",
    x"BF2307AB",
    x"BF230C84",
    x"BF23115C",
    x"BF231633",
    x"BF231B0B",
    x"BF231FE3",
    x"BF2324BB",
    x"BF232992",
    x"BF232E6A",
    x"BF233341",
    x"BF233818",
    x"BF233CEF",
    x"BF2341C6",
    x"BF23469D",
    x"BF234B74",
    x"BF23504B",
    x"BF235521",
    x"BF2359F8",
    x"BF235ECE",
    x"BF2363A5",
    x"BF23687B",
    x"BF236D51",
    x"BF237227",
    x"BF2376FD",
    x"BF237BD3",
    x"BF2380A8",
    x"BF23857E",
    x"BF238A54",
    x"BF238F29",
    x"BF2393FE",
    x"BF2398D4",
    x"BF239DA9",
    x"BF23A27E",
    x"BF23A753",
    x"BF23AC28",
    x"BF23B0FC",
    x"BF23B5D1",
    x"BF23BAA6",
    x"BF23BF7A",
    x"BF23C44F",
    x"BF23C923",
    x"BF23CDF7",
    x"BF23D2CB",
    x"BF23D79F",
    x"BF23DC73",
    x"BF23E147",
    x"BF23E61A",
    x"BF23EAEE",
    x"BF23EFC1",
    x"BF23F495",
    x"BF23F968",
    x"BF23FE3B",
    x"BF24030E",
    x"BF2407E1",
    x"BF240CB4",
    x"BF241187",
    x"BF24165A",
    x"BF241B2C",
    x"BF241FFF",
    x"BF2424D1",
    x"BF2429A3",
    x"BF242E75",
    x"BF243348",
    x"BF24381A",
    x"BF243CEB",
    x"BF2441BD",
    x"BF24468F",
    x"BF244B60",
    x"BF245032",
    x"BF245503",
    x"BF2459D5",
    x"BF245EA6",
    x"BF246377",
    x"BF246848",
    x"BF246D19",
    x"BF2471EA",
    x"BF2476BA",
    x"BF247B8B",
    x"BF24805B",
    x"BF24852C",
    x"BF2489FC",
    x"BF248ECC",
    x"BF24939C",
    x"BF24986D",
    x"BF249D3C",
    x"BF24A20C",
    x"BF24A6DC",
    x"BF24ABAC",
    x"BF24B07B",
    x"BF24B54A",
    x"BF24BA1A",
    x"BF24BEE9",
    x"BF24C3B8",
    x"BF24C887",
    x"BF24CD56",
    x"BF24D225",
    x"BF24D6F4",
    x"BF24DBC2",
    x"BF24E091",
    x"BF24E55F",
    x"BF24EA2D",
    x"BF24EEFC",
    x"BF24F3CA",
    x"BF24F898",
    x"BF24FD66",
    x"BF250234",
    x"BF250701",
    x"BF250BCF",
    x"BF25109C",
    x"BF25156A",
    x"BF251A37",
    x"BF251F04",
    x"BF2523D2",
    x"BF25289F",
    x"BF252D6C",
    x"BF253238",
    x"BF253705",
    x"BF253BD2",
    x"BF25409E",
    x"BF25456B",
    x"BF254A37",
    x"BF254F03",
    x"BF2553CF",
    x"BF25589B",
    x"BF255D67",
    x"BF256233",
    x"BF2566FF",
    x"BF256BCB",
    x"BF257096",
    x"BF257562",
    x"BF257A2D",
    x"BF257EF8",
    x"BF2583C3",
    x"BF25888E",
    x"BF258D59",
    x"BF259224",
    x"BF2596EF",
    x"BF259BB9",
    x"BF25A084",
    x"BF25A54E",
    x"BF25AA19",
    x"BF25AEE3",
    x"BF25B3AD",
    x"BF25B877",
    x"BF25BD41",
    x"BF25C20B",
    x"BF25C6D5",
    x"BF25CB9E",
    x"BF25D068",
    x"BF25D531",
    x"BF25D9FB",
    x"BF25DEC4",
    x"BF25E38D",
    x"BF25E856",
    x"BF25ED1F",
    x"BF25F1E8",
    x"BF25F6B1",
    x"BF25FB79",
    x"BF260042",
    x"BF26050A",
    x"BF2609D3",
    x"BF260E9B",
    x"BF261363",
    x"BF26182B",
    x"BF261CF3",
    x"BF2621BB",
    x"BF262682",
    x"BF262B4A",
    x"BF263012",
    x"BF2634D9",
    x"BF2639A0",
    x"BF263E68",
    x"BF26432F",
    x"BF2647F6",
    x"BF264CBD",
    x"BF265184",
    x"BF26564A",
    x"BF265B11",
    x"BF265FD8",
    x"BF26649E",
    x"BF266964",
    x"BF266E2B",
    x"BF2672F1",
    x"BF2677B7",
    x"BF267C7D",
    x"BF268143",
    x"BF268608",
    x"BF268ACE",
    x"BF268F93",
    x"BF269459",
    x"BF26991E",
    x"BF269DE3",
    x"BF26A2A9",
    x"BF26A76E",
    x"BF26AC33",
    x"BF26B0F7",
    x"BF26B5BC",
    x"BF26BA81",
    x"BF26BF45",
    x"BF26C40A",
    x"BF26C8CE",
    x"BF26CD92",
    x"BF26D256",
    x"BF26D71A",
    x"BF26DBDE",
    x"BF26E0A2",
    x"BF26E566",
    x"BF26EA2A",
    x"BF26EEED",
    x"BF26F3B0",
    x"BF26F874",
    x"BF26FD37",
    x"BF2701FA",
    x"BF2706BD",
    x"BF270B80",
    x"BF271043",
    x"BF271506",
    x"BF2719C8",
    x"BF271E8B",
    x"BF27234D",
    x"BF272810",
    x"BF272CD2",
    x"BF273194",
    x"BF273656",
    x"BF273B18",
    x"BF273FDA",
    x"BF27449B",
    x"BF27495D",
    x"BF274E1E",
    x"BF2752E0",
    x"BF2757A1",
    x"BF275C62",
    x"BF276123",
    x"BF2765E5",
    x"BF276AA5",
    x"BF276F66",
    x"BF277427",
    x"BF2778E8",
    x"BF277DA8",
    x"BF278268",
    x"BF278729",
    x"BF278BE9",
    x"BF2790A9",
    x"BF279569",
    x"BF279A29",
    x"BF279EE9",
    x"BF27A3A8",
    x"BF27A868",
    x"BF27AD28",
    x"BF27B1E7",
    x"BF27B6A6",
    x"BF27BB65",
    x"BF27C025",
    x"BF27C4E4",
    x"BF27C9A2",
    x"BF27CE61",
    x"BF27D320",
    x"BF27D7DE",
    x"BF27DC9D",
    x"BF27E15B",
    x"BF27E61A",
    x"BF27EAD8",
    x"BF27EF96",
    x"BF27F454",
    x"BF27F912",
    x"BF27FDD0",
    x"BF28028D",
    x"BF28074B",
    x"BF280C08",
    x"BF2810C6",
    x"BF281583",
    x"BF281A40",
    x"BF281EFD",
    x"BF2823BA",
    x"BF282877",
    x"BF282D34",
    x"BF2831F0",
    x"BF2836AD",
    x"BF283B69",
    x"BF284026",
    x"BF2844E2",
    x"BF28499E",
    x"BF284E5A",
    x"BF285316",
    x"BF2857D2",
    x"BF285C8E",
    x"BF286149",
    x"BF286605",
    x"BF286AC0",
    x"BF286F7C",
    x"BF287437",
    x"BF2878F2",
    x"BF287DAD",
    x"BF288268",
    x"BF288723",
    x"BF288BDE",
    x"BF289098",
    x"BF289553",
    x"BF289A0D",
    x"BF289EC8",
    x"BF28A382",
    x"BF28A83C",
    x"BF28ACF6",
    x"BF28B1B0",
    x"BF28B66A",
    x"BF28BB23",
    x"BF28BFDD",
    x"BF28C497",
    x"BF28C950",
    x"BF28CE09",
    x"BF28D2C3",
    x"BF28D77C",
    x"BF28DC35",
    x"BF28E0EE",
    x"BF28E5A6",
    x"BF28EA5F",
    x"BF28EF18",
    x"BF28F3D0",
    x"BF28F889",
    x"BF28FD41",
    x"BF2901F9",
    x"BF2906B1",
    x"BF290B69",
    x"BF291021",
    x"BF2914D9",
    x"BF291991",
    x"BF291E48",
    x"BF292300",
    x"BF2927B7",
    x"BF292C6E",
    x"BF293125",
    x"BF2935DD",
    x"BF293A93",
    x"BF293F4A",
    x"BF294401",
    x"BF2948B8",
    x"BF294D6E",
    x"BF295225",
    x"BF2956DB",
    x"BF295B91",
    x"BF296048",
    x"BF2964FE",
    x"BF2969B4",
    x"BF296E69",
    x"BF29731F",
    x"BF2977D5",
    x"BF297C8A",
    x"BF298140",
    x"BF2985F5",
    x"BF298AAA",
    x"BF298F60",
    x"BF299415",
    x"BF2998CA",
    x"BF299D7E",
    x"BF29A233",
    x"BF29A6E8",
    x"BF29AB9C",
    x"BF29B051",
    x"BF29B505",
    x"BF29B9B9",
    x"BF29BE6D",
    x"BF29C321",
    x"BF29C7D5",
    x"BF29CC89",
    x"BF29D13D",
    x"BF29D5F0",
    x"BF29DAA4",
    x"BF29DF57",
    x"BF29E40B",
    x"BF29E8BE",
    x"BF29ED71",
    x"BF29F224",
    x"BF29F6D7",
    x"BF29FB89",
    x"BF2A003C",
    x"BF2A04EF",
    x"BF2A09A1",
    x"BF2A0E54",
    x"BF2A1306",
    x"BF2A17B8",
    x"BF2A1C6A",
    x"BF2A211C",
    x"BF2A25CE",
    x"BF2A2A80",
    x"BF2A2F31",
    x"BF2A33E3",
    x"BF2A3894",
    x"BF2A3D46",
    x"BF2A41F7",
    x"BF2A46A8",
    x"BF2A4B59",
    x"BF2A500A",
    x"BF2A54BB",
    x"BF2A596C",
    x"BF2A5E1C",
    x"BF2A62CD",
    x"BF2A677D",
    x"BF2A6C2E",
    x"BF2A70DE",
    x"BF2A758E",
    x"BF2A7A3E",
    x"BF2A7EEE",
    x"BF2A839E",
    x"BF2A884D",
    x"BF2A8CFD",
    x"BF2A91AC",
    x"BF2A965C",
    x"BF2A9B0B",
    x"BF2A9FBA",
    x"BF2AA469",
    x"BF2AA918",
    x"BF2AADC7",
    x"BF2AB276",
    x"BF2AB725",
    x"BF2ABBD3",
    x"BF2AC082",
    x"BF2AC530",
    x"BF2AC9DE",
    x"BF2ACE8D",
    x"BF2AD33B",
    x"BF2AD7E9",
    x"BF2ADC96",
    x"BF2AE144",
    x"BF2AE5F2",
    x"BF2AEA9F",
    x"BF2AEF4D",
    x"BF2AF3FA",
    x"BF2AF8A7",
    x"BF2AFD55",
    x"BF2B0202",
    x"BF2B06AF",
    x"BF2B0B5B",
    x"BF2B1008",
    x"BF2B14B5",
    x"BF2B1961",
    x"BF2B1E0E",
    x"BF2B22BA",
    x"BF2B2766",
    x"BF2B2C12",
    x"BF2B30BE",
    x"BF2B356A",
    x"BF2B3A16",
    x"BF2B3EC2",
    x"BF2B436D",
    x"BF2B4819",
    x"BF2B4CC4",
    x"BF2B516F",
    x"BF2B561B",
    x"BF2B5AC6",
    x"BF2B5F71",
    x"BF2B641B",
    x"BF2B68C6",
    x"BF2B6D71",
    x"BF2B721B",
    x"BF2B76C6",
    x"BF2B7B70",
    x"BF2B801A",
    x"BF2B84C5",
    x"BF2B896F",
    x"BF2B8E19",
    x"BF2B92C2",
    x"BF2B976C",
    x"BF2B9C16",
    x"BF2BA0BF",
    x"BF2BA569",
    x"BF2BAA12",
    x"BF2BAEBB",
    x"BF2BB364",
    x"BF2BB80D",
    x"BF2BBCB6",
    x"BF2BC15F",
    x"BF2BC608",
    x"BF2BCAB0",
    x"BF2BCF59",
    x"BF2BD401",
    x"BF2BD8AA",
    x"BF2BDD52",
    x"BF2BE1FA",
    x"BF2BE6A2",
    x"BF2BEB4A",
    x"BF2BEFF1",
    x"BF2BF499",
    x"BF2BF941",
    x"BF2BFDE8",
    x"BF2C028F",
    x"BF2C0737",
    x"BF2C0BDE",
    x"BF2C1085",
    x"BF2C152C",
    x"BF2C19D3",
    x"BF2C1E79",
    x"BF2C2320",
    x"BF2C27C7",
    x"BF2C2C6D",
    x"BF2C3113",
    x"BF2C35B9",
    x"BF2C3A60",
    x"BF2C3F06",
    x"BF2C43AB",
    x"BF2C4851",
    x"BF2C4CF7",
    x"BF2C519D",
    x"BF2C5642",
    x"BF2C5AE7",
    x"BF2C5F8D",
    x"BF2C6432",
    x"BF2C68D7",
    x"BF2C6D7C",
    x"BF2C7221",
    x"BF2C76C5",
    x"BF2C7B6A",
    x"BF2C800F",
    x"BF2C84B3",
    x"BF2C8957",
    x"BF2C8DFC",
    x"BF2C92A0",
    x"BF2C9744",
    x"BF2C9BE8",
    x"BF2CA08C",
    x"BF2CA52F",
    x"BF2CA9D3",
    x"BF2CAE76",
    x"BF2CB31A",
    x"BF2CB7BD",
    x"BF2CBC60",
    x"BF2CC103",
    x"BF2CC5A6",
    x"BF2CCA49",
    x"BF2CCEEC",
    x"BF2CD38F",
    x"BF2CD831",
    x"BF2CDCD4",
    x"BF2CE176",
    x"BF2CE618",
    x"BF2CEABB",
    x"BF2CEF5D",
    x"BF2CF3FF",
    x"BF2CF8A0",
    x"BF2CFD42",
    x"BF2D01E4",
    x"BF2D0685",
    x"BF2D0B27",
    x"BF2D0FC8",
    x"BF2D1469",
    x"BF2D190A",
    x"BF2D1DAB",
    x"BF2D224C",
    x"BF2D26ED",
    x"BF2D2B8E",
    x"BF2D302E",
    x"BF2D34CF",
    x"BF2D396F",
    x"BF2D3E10",
    x"BF2D42B0",
    x"BF2D4750",
    x"BF2D4BF0",
    x"BF2D5090",
    x"BF2D552F",
    x"BF2D59CF",
    x"BF2D5E6F",
    x"BF2D630E",
    x"BF2D67AD",
    x"BF2D6C4D",
    x"BF2D70EC",
    x"BF2D758B",
    x"BF2D7A2A",
    x"BF2D7EC9",
    x"BF2D8367",
    x"BF2D8806",
    x"BF2D8CA4",
    x"BF2D9143",
    x"BF2D95E1",
    x"BF2D9A7F",
    x"BF2D9F1D",
    x"BF2DA3BB",
    x"BF2DA859",
    x"BF2DACF7",
    x"BF2DB195",
    x"BF2DB632",
    x"BF2DBAD0",
    x"BF2DBF6D",
    x"BF2DC40A",
    x"BF2DC8A7",
    x"BF2DCD44",
    x"BF2DD1E1",
    x"BF2DD67E",
    x"BF2DDB1B",
    x"BF2DDFB8",
    x"BF2DE454",
    x"BF2DE8F0",
    x"BF2DED8D",
    x"BF2DF229",
    x"BF2DF6C5",
    x"BF2DFB61",
    x"BF2DFFFD",
    x"BF2E0499",
    x"BF2E0934",
    x"BF2E0DD0",
    x"BF2E126B",
    x"BF2E1707",
    x"BF2E1BA2",
    x"BF2E203D",
    x"BF2E24D8",
    x"BF2E2973",
    x"BF2E2E0E",
    x"BF2E32A9",
    x"BF2E3743",
    x"BF2E3BDE",
    x"BF2E4078",
    x"BF2E4513",
    x"BF2E49AD",
    x"BF2E4E47",
    x"BF2E52E1",
    x"BF2E577B",
    x"BF2E5C15",
    x"BF2E60AE",
    x"BF2E6548",
    x"BF2E69E1",
    x"BF2E6E7B",
    x"BF2E7314",
    x"BF2E77AD",
    x"BF2E7C46",
    x"BF2E80DF",
    x"BF2E8578",
    x"BF2E8A11",
    x"BF2E8EA9",
    x"BF2E9342",
    x"BF2E97DA",
    x"BF2E9C73",
    x"BF2EA10B",
    x"BF2EA5A3",
    x"BF2EAA3B",
    x"BF2EAED3",
    x"BF2EB36B",
    x"BF2EB802",
    x"BF2EBC9A",
    x"BF2EC131",
    x"BF2EC5C9",
    x"BF2ECA60",
    x"BF2ECEF7",
    x"BF2ED38E",
    x"BF2ED825",
    x"BF2EDCBC",
    x"BF2EE153",
    x"BF2EE5E9",
    x"BF2EEA80",
    x"BF2EEF16",
    x"BF2EF3AD",
    x"BF2EF843",
    x"BF2EFCD9",
    x"BF2F016F",
    x"BF2F0605",
    x"BF2F0A9B",
    x"BF2F0F30",
    x"BF2F13C6",
    x"BF2F185B",
    x"BF2F1CF1",
    x"BF2F2186",
    x"BF2F261B",
    x"BF2F2AB0",
    x"BF2F2F45",
    x"BF2F33DA",
    x"BF2F386F",
    x"BF2F3D03",
    x"BF2F4198",
    x"BF2F462C",
    x"BF2F4AC1",
    x"BF2F4F55",
    x"BF2F53E9",
    x"BF2F587D",
    x"BF2F5D11",
    x"BF2F61A5",
    x"BF2F6638",
    x"BF2F6ACC",
    x"BF2F6F5F",
    x"BF2F73F3",
    x"BF2F7886",
    x"BF2F7D19",
    x"BF2F81AC",
    x"BF2F863F",
    x"BF2F8AD2",
    x"BF2F8F65",
    x"BF2F93F7",
    x"BF2F988A",
    x"BF2F9D1C",
    x"BF2FA1AF",
    x"BF2FA641",
    x"BF2FAAD3",
    x"BF2FAF65",
    x"BF2FB3F7",
    x"BF2FB888",
    x"BF2FBD1A",
    x"BF2FC1AC",
    x"BF2FC63D",
    x"BF2FCACF",
    x"BF2FCF60",
    x"BF2FD3F1",
    x"BF2FD882",
    x"BF2FDD13",
    x"BF2FE1A4",
    x"BF2FE634",
    x"BF2FEAC5",
    x"BF2FEF56",
    x"BF2FF3E6",
    x"BF2FF876",
    x"BF2FFD06",
    x"BF300196",
    x"BF300626",
    x"BF300AB6",
    x"BF300F46",
    x"BF3013D6",
    x"BF301865",
    x"BF301CF5",
    x"BF302184",
    x"BF302613",
    x"BF302AA2",
    x"BF302F31",
    x"BF3033C0",
    x"BF30384F",
    x"BF303CDE",
    x"BF30416C",
    x"BF3045FB",
    x"BF304A89",
    x"BF304F18",
    x"BF3053A6",
    x"BF305834",
    x"BF305CC2",
    x"BF306150",
    x"BF3065DD",
    x"BF306A6B",
    x"BF306EF9",
    x"BF307386",
    x"BF307813",
    x"BF307CA1",
    x"BF30812E",
    x"BF3085BB",
    x"BF308A48",
    x"BF308ED4",
    x"BF309361",
    x"BF3097EE",
    x"BF309C7A",
    x"BF30A106",
    x"BF30A593",
    x"BF30AA1F",
    x"BF30AEAB",
    x"BF30B337",
    x"BF30B7C3",
    x"BF30BC4E",
    x"BF30C0DA",
    x"BF30C566",
    x"BF30C9F1",
    x"BF30CE7C",
    x"BF30D307",
    x"BF30D792",
    x"BF30DC1D",
    x"BF30E0A8",
    x"BF30E533",
    x"BF30E9BE",
    x"BF30EE48",
    x"BF30F2D3",
    x"BF30F75D",
    x"BF30FBE7",
    x"BF310071",
    x"BF3104FB",
    x"BF310985",
    x"BF310E0F",
    x"BF311299",
    x"BF311722",
    x"BF311BAC",
    x"BF312035",
    x"BF3124BF",
    x"BF312948",
    x"BF312DD1",
    x"BF31325A",
    x"BF3136E3",
    x"BF313B6B",
    x"BF313FF4",
    x"BF31447D",
    x"BF314905",
    x"BF314D8D",
    x"BF315215",
    x"BF31569E",
    x"BF315B26",
    x"BF315FAD",
    x"BF316435",
    x"BF3168BD",
    x"BF316D44",
    x"BF3171CC",
    x"BF317653",
    x"BF317ADB",
    x"BF317F62",
    x"BF3183E9",
    x"BF318870",
    x"BF318CF6",
    x"BF31917D",
    x"BF319604",
    x"BF319A8A",
    x"BF319F11",
    x"BF31A397",
    x"BF31A81D",
    x"BF31ACA3",
    x"BF31B129",
    x"BF31B5AF",
    x"BF31BA35",
    x"BF31BEBA",
    x"BF31C340",
    x"BF31C7C5",
    x"BF31CC4B",
    x"BF31D0D0",
    x"BF31D555",
    x"BF31D9DA",
    x"BF31DE5F",
    x"BF31E2E4",
    x"BF31E768",
    x"BF31EBED",
    x"BF31F071",
    x"BF31F4F6",
    x"BF31F97A",
    x"BF31FDFE",
    x"BF320282",
    x"BF320706",
    x"BF320B8A",
    x"BF32100E",
    x"BF321491",
    x"BF321915",
    x"BF321D98",
    x"BF32221B",
    x"BF32269E",
    x"BF322B22",
    x"BF322FA5",
    x"BF323427",
    x"BF3238AA",
    x"BF323D2D",
    x"BF3241AF",
    x"BF324632",
    x"BF324AB4",
    x"BF324F36",
    x"BF3253B8",
    x"BF32583A",
    x"BF325CBC",
    x"BF32613E",
    x"BF3265C0",
    x"BF326A41",
    x"BF326EC3",
    x"BF327344",
    x"BF3277C5",
    x"BF327C46",
    x"BF3280C7",
    x"BF328548",
    x"BF3289C9",
    x"BF328E4A",
    x"BF3292CA",
    x"BF32974B",
    x"BF329BCB",
    x"BF32A04C",
    x"BF32A4CC",
    x"BF32A94C",
    x"BF32ADCC",
    x"BF32B24C",
    x"BF32B6CB",
    x"BF32BB4B",
    x"BF32BFCA",
    x"BF32C44A",
    x"BF32C8C9",
    x"BF32CD48",
    x"BF32D1C7",
    x"BF32D646",
    x"BF32DAC5",
    x"BF32DF44",
    x"BF32E3C3",
    x"BF32E841",
    x"BF32ECC0",
    x"BF32F13E",
    x"BF32F5BC",
    x"BF32FA3A",
    x"BF32FEB8",
    x"BF330336",
    x"BF3307B4",
    x"BF330C32",
    x"BF3310AF",
    x"BF33152D",
    x"BF3319AA",
    x"BF331E27",
    x"BF3322A5",
    x"BF332722",
    x"BF332B9F",
    x"BF33301B",
    x"BF333498",
    x"BF333915",
    x"BF333D91",
    x"BF33420E",
    x"BF33468A",
    x"BF334B06",
    x"BF334F82",
    x"BF3353FE",
    x"BF33587A",
    x"BF335CF6",
    x"BF336171",
    x"BF3365ED",
    x"BF336A68",
    x"BF336EE4",
    x"BF33735F",
    x"BF3377DA",
    x"BF337C55",
    x"BF3380D0",
    x"BF33854B",
    x"BF3389C5",
    x"BF338E40",
    x"BF3392BA",
    x"BF339735",
    x"BF339BAF",
    x"BF33A029",
    x"BF33A4A3",
    x"BF33A91D",
    x"BF33AD97",
    x"BF33B210",
    x"BF33B68A",
    x"BF33BB03",
    x"BF33BF7D",
    x"BF33C3F6",
    x"BF33C86F",
    x"BF33CCE8",
    x"BF33D161",
    x"BF33D5DA",
    x"BF33DA53",
    x"BF33DECB",
    x"BF33E344",
    x"BF33E7BC",
    x"BF33EC34",
    x"BF33F0AD",
    x"BF33F525",
    x"BF33F99D",
    x"BF33FE14",
    x"BF34028C",
    x"BF340704",
    x"BF340B7B",
    x"BF340FF3",
    x"BF34146A",
    x"BF3418E1",
    x"BF341D58",
    x"BF3421CF",
    x"BF342646",
    x"BF342ABD",
    x"BF342F34",
    x"BF3433AA",
    x"BF343821",
    x"BF343C97",
    x"BF34410D",
    x"BF344583",
    x"BF3449F9",
    x"BF344E6F",
    x"BF3452E5",
    x"BF34575B",
    x"BF345BD0",
    x"BF346046",
    x"BF3464BB",
    x"BF346930",
    x"BF346DA5",
    x"BF34721A",
    x"BF34768F",
    x"BF347B04",
    x"BF347F79",
    x"BF3483ED",
    x"BF348862",
    x"BF348CD6",
    x"BF34914B",
    x"BF3495BF",
    x"BF349A33",
    x"BF349EA7",
    x"BF34A31B",
    x"BF34A78E",
    x"BF34AC02",
    x"BF34B075",
    x"BF34B4E9",
    x"BF34B95C",
    x"BF34BDCF",
    x"BF34C242",
    x"BF34C6B5",
    x"BF34CB28",
    x"BF34CF9B",
    x"BF34D40D",
    x"BF34D880",
    x"BF34DCF2",
    x"BF34E165",
    x"BF34E5D7",
    x"BF34EA49",
    x"BF34EEBB",
    x"BF34F32D",
    x"BF34F79F",
    x"BF34FC10",
    x"BF350082",
    x"BF3504F3",
    x"BF350965",
    x"BF350DD6",
    x"BF351247",
    x"BF3516B8",
    x"BF351B29",
    x"BF351F9A",
    x"BF35240A",
    x"BF35287B",
    x"BF352CEB",
    x"BF35315C",
    x"BF3535CC",
    x"BF353A3C",
    x"BF353EAC",
    x"BF35431C",
    x"BF35478C",
    x"BF354BFB",
    x"BF35506B",
    x"BF3554DA",
    x"BF35594A",
    x"BF355DB9",
    x"BF356228",
    x"BF356697",
    x"BF356B06",
    x"BF356F75",
    x"BF3573E4",
    x"BF357852",
    x"BF357CC1",
    x"BF35812F",
    x"BF35859D",
    x"BF358A0B",
    x"BF358E79",
    x"BF3592E7",
    x"BF359755",
    x"BF359BC3",
    x"BF35A031",
    x"BF35A49E",
    x"BF35A90B",
    x"BF35AD79",
    x"BF35B1E6",
    x"BF35B653",
    x"BF35BAC0",
    x"BF35BF2D",
    x"BF35C39A",
    x"BF35C806",
    x"BF35CC73",
    x"BF35D0DF",
    x"BF35D54B",
    x"BF35D9B8",
    x"BF35DE24",
    x"BF35E290",
    x"BF35E6FB",
    x"BF35EB67",
    x"BF35EFD3",
    x"BF35F43E",
    x"BF35F8AA",
    x"BF35FD15",
    x"BF360180",
    x"BF3605EB",
    x"BF360A56",
    x"BF360EC1",
    x"BF36132C",
    x"BF361797",
    x"BF361C01",
    x"BF36206C",
    x"BF3624D6",
    x"BF362940",
    x"BF362DAA",
    x"BF363214",
    x"BF36367E",
    x"BF363AE8",
    x"BF363F52",
    x"BF3643BB",
    x"BF364825",
    x"BF364C8E",
    x"BF3650F7",
    x"BF365560",
    x"BF3659C9",
    x"BF365E32",
    x"BF36629B",
    x"BF366704",
    x"BF366B6C",
    x"BF366FD5",
    x"BF36743D",
    x"BF3678A5",
    x"BF367D0D",
    x"BF368175",
    x"BF3685DD",
    x"BF368A45",
    x"BF368EAD",
    x"BF369314",
    x"BF36977C",
    x"BF369BE3",
    x"BF36A04A",
    x"BF36A4B2",
    x"BF36A919",
    x"BF36AD7F",
    x"BF36B1E6",
    x"BF36B64D",
    x"BF36BAB4",
    x"BF36BF1A",
    x"BF36C380",
    x"BF36C7E7",
    x"BF36CC4D",
    x"BF36D0B3",
    x"BF36D519",
    x"BF36D97F",
    x"BF36DDE4",
    x"BF36E24A",
    x"BF36E6AF",
    x"BF36EB15",
    x"BF36EF7A",
    x"BF36F3DF",
    x"BF36F844",
    x"BF36FCA9",
    x"BF37010E",
    x"BF370573",
    x"BF3709D7",
    x"BF370E3C",
    x"BF3712A0",
    x"BF371704",
    x"BF371B69",
    x"BF371FCD",
    x"BF372431",
    x"BF372894",
    x"BF372CF8",
    x"BF37315C",
    x"BF3735BF",
    x"BF373A23",
    x"BF373E86",
    x"BF3742E9",
    x"BF37474C",
    x"BF374BAF",
    x"BF375012",
    x"BF375475",
    x"BF3758D7",
    x"BF375D3A",
    x"BF37619C",
    x"BF3765FE",
    x"BF376A61",
    x"BF376EC3",
    x"BF377325",
    x"BF377787",
    x"BF377BE8",
    x"BF37804A",
    x"BF3784AB",
    x"BF37890D",
    x"BF378D6E",
    x"BF3791CF",
    x"BF379630",
    x"BF379A91",
    x"BF379EF2",
    x"BF37A353",
    x"BF37A7B4",
    x"BF37AC14",
    x"BF37B074",
    x"BF37B4D5",
    x"BF37B935",
    x"BF37BD95",
    x"BF37C1F5",
    x"BF37C655",
    x"BF37CAB5",
    x"BF37CF14",
    x"BF37D374",
    x"BF37D7D3",
    x"BF37DC32",
    x"BF37E092",
    x"BF37E4F1",
    x"BF37E950",
    x"BF37EDAF",
    x"BF37F20D",
    x"BF37F66C",
    x"BF37FACA",
    x"BF37FF29",
    x"BF380387",
    x"BF3807E5",
    x"BF380C43",
    x"BF3810A1",
    x"BF3814FF",
    x"BF38195D",
    x"BF381DBB",
    x"BF382218",
    x"BF382676",
    x"BF382AD3",
    x"BF382F30",
    x"BF38338D",
    x"BF3837EA",
    x"BF383C47",
    x"BF3840A4",
    x"BF384500",
    x"BF38495D",
    x"BF384DB9",
    x"BF385216",
    x"BF385672",
    x"BF385ACE",
    x"BF385F2A",
    x"BF386386",
    x"BF3867E1",
    x"BF386C3D",
    x"BF387099",
    x"BF3874F4",
    x"BF38794F",
    x"BF387DAB",
    x"BF388206",
    x"BF388661",
    x"BF388ABB",
    x"BF388F16",
    x"BF389371",
    x"BF3897CB",
    x"BF389C26",
    x"BF38A080",
    x"BF38A4DA",
    x"BF38A934",
    x"BF38AD8E",
    x"BF38B1E8",
    x"BF38B642",
    x"BF38BA9C",
    x"BF38BEF5",
    x"BF38C34F",
    x"BF38C7A8",
    x"BF38CC01",
    x"BF38D05A",
    x"BF38D4B3",
    x"BF38D90C",
    x"BF38DD65",
    x"BF38E1BD",
    x"BF38E616",
    x"BF38EA6E",
    x"BF38EEC7",
    x"BF38F31F",
    x"BF38F777",
    x"BF38FBCF",
    x"BF390027",
    x"BF39047E",
    x"BF3908D6",
    x"BF390D2E",
    x"BF391185",
    x"BF3915DC",
    x"BF391A33",
    x"BF391E8B",
    x"BF3922E1",
    x"BF392738",
    x"BF392B8F",
    x"BF392FE6",
    x"BF39343C",
    x"BF393893",
    x"BF393CE9",
    x"BF39413F",
    x"BF394595",
    x"BF3949EB",
    x"BF394E41",
    x"BF395297",
    x"BF3956EC",
    x"BF395B42",
    x"BF395F97",
    x"BF3963ED",
    x"BF396842",
    x"BF396C97",
    x"BF3970EC",
    x"BF397541",
    x"BF397995",
    x"BF397DEA",
    x"BF39823E",
    x"BF398693",
    x"BF398AE7",
    x"BF398F3B",
    x"BF39938F",
    x"BF3997E3",
    x"BF399C37",
    x"BF39A08B",
    x"BF39A4DF",
    x"BF39A932",
    x"BF39AD85",
    x"BF39B1D9",
    x"BF39B62C",
    x"BF39BA7F",
    x"BF39BED2",
    x"BF39C325",
    x"BF39C777",
    x"BF39CBCA",
    x"BF39D01D",
    x"BF39D46F",
    x"BF39D8C1",
    x"BF39DD13",
    x"BF39E165",
    x"BF39E5B7",
    x"BF39EA09",
    x"BF39EE5B",
    x"BF39F2AC",
    x"BF39F6FE",
    x"BF39FB4F",
    x"BF39FFA1",
    x"BF3A03F2",
    x"BF3A0843",
    x"BF3A0C94",
    x"BF3A10E4",
    x"BF3A1535",
    x"BF3A1986",
    x"BF3A1DD6",
    x"BF3A2227",
    x"BF3A2677",
    x"BF3A2AC7",
    x"BF3A2F17",
    x"BF3A3367",
    x"BF3A37B7",
    x"BF3A3C06",
    x"BF3A4056",
    x"BF3A44A6",
    x"BF3A48F5",
    x"BF3A4D44",
    x"BF3A5193",
    x"BF3A55E2",
    x"BF3A5A31",
    x"BF3A5E80",
    x"BF3A62CF",
    x"BF3A671D",
    x"BF3A6B6C",
    x"BF3A6FBA",
    x"BF3A7408",
    x"BF3A7856",
    x"BF3A7CA4",
    x"BF3A80F2",
    x"BF3A8540",
    x"BF3A898E",
    x"BF3A8DDB",
    x"BF3A9229",
    x"BF3A9676",
    x"BF3A9AC3",
    x"BF3A9F10",
    x"BF3AA35D",
    x"BF3AA7AA",
    x"BF3AABF7",
    x"BF3AB044",
    x"BF3AB490",
    x"BF3AB8DD",
    x"BF3ABD29",
    x"BF3AC175",
    x"BF3AC5C1",
    x"BF3ACA0D",
    x"BF3ACE59",
    x"BF3AD2A5",
    x"BF3AD6F1",
    x"BF3ADB3C",
    x"BF3ADF88",
    x"BF3AE3D3",
    x"BF3AE81E",
    x"BF3AEC69",
    x"BF3AF0B4",
    x"BF3AF4FF",
    x"BF3AF94A",
    x"BF3AFD94",
    x"BF3B01DF",
    x"BF3B0629",
    x"BF3B0A74",
    x"BF3B0EBE",
    x"BF3B1308",
    x"BF3B1752",
    x"BF3B1B9C",
    x"BF3B1FE5",
    x"BF3B242F",
    x"BF3B2879",
    x"BF3B2CC2",
    x"BF3B310B",
    x"BF3B3554",
    x"BF3B399E",
    x"BF3B3DE6",
    x"BF3B422F",
    x"BF3B4678",
    x"BF3B4AC1",
    x"BF3B4F09",
    x"BF3B5351",
    x"BF3B579A",
    x"BF3B5BE2",
    x"BF3B602A",
    x"BF3B6472",
    x"BF3B68BA",
    x"BF3B6D01",
    x"BF3B7149",
    x"BF3B7590",
    x"BF3B79D8",
    x"BF3B7E1F",
    x"BF3B8266",
    x"BF3B86AD",
    x"BF3B8AF4",
    x"BF3B8F3B",
    x"BF3B9382",
    x"BF3B97C8",
    x"BF3B9C0F",
    x"BF3BA055",
    x"BF3BA49B",
    x"BF3BA8E1",
    x"BF3BAD27",
    x"BF3BB16D",
    x"BF3BB5B3",
    x"BF3BB9F9",
    x"BF3BBE3E",
    x"BF3BC284",
    x"BF3BC6C9",
    x"BF3BCB0E",
    x"BF3BCF53",
    x"BF3BD398",
    x"BF3BD7DD",
    x"BF3BDC22",
    x"BF3BE067",
    x"BF3BE4AB",
    x"BF3BE8F0",
    x"BF3BED34",
    x"BF3BF178",
    x"BF3BF5BC",
    x"BF3BFA00",
    x"BF3BFE44",
    x"BF3C0288",
    x"BF3C06CB",
    x"BF3C0B0F",
    x"BF3C0F52",
    x"BF3C1396",
    x"BF3C17D9",
    x"BF3C1C1C",
    x"BF3C205F",
    x"BF3C24A2",
    x"BF3C28E4",
    x"BF3C2D27",
    x"BF3C316A",
    x"BF3C35AC",
    x"BF3C39EE",
    x"BF3C3E30",
    x"BF3C4272",
    x"BF3C46B4",
    x"BF3C4AF6",
    x"BF3C4F38",
    x"BF3C5379",
    x"BF3C57BB",
    x"BF3C5BFC",
    x"BF3C603E",
    x"BF3C647F",
    x"BF3C68C0",
    x"BF3C6D01",
    x"BF3C7141",
    x"BF3C7582",
    x"BF3C79C3",
    x"BF3C7E03",
    x"BF3C8244",
    x"BF3C8684",
    x"BF3C8AC4",
    x"BF3C8F04",
    x"BF3C9344",
    x"BF3C9784",
    x"BF3C9BC3",
    x"BF3CA003",
    x"BF3CA442",
    x"BF3CA881",
    x"BF3CACC1",
    x"BF3CB100",
    x"BF3CB53F",
    x"BF3CB97E",
    x"BF3CBDBC",
    x"BF3CC1FB",
    x"BF3CC63A",
    x"BF3CCA78",
    x"BF3CCEB6",
    x"BF3CD2F4",
    x"BF3CD733",
    x"BF3CDB70",
    x"BF3CDFAE",
    x"BF3CE3EC",
    x"BF3CE82A",
    x"BF3CEC67",
    x"BF3CF0A5",
    x"BF3CF4E2",
    x"BF3CF91F",
    x"BF3CFD5C",
    x"BF3D0199",
    x"BF3D05D6",
    x"BF3D0A12",
    x"BF3D0E4F",
    x"BF3D128C",
    x"BF3D16C8",
    x"BF3D1B04",
    x"BF3D1F40",
    x"BF3D237C",
    x"BF3D27B8",
    x"BF3D2BF4",
    x"BF3D3030",
    x"BF3D346B",
    x"BF3D38A7",
    x"BF3D3CE2",
    x"BF3D411D",
    x"BF3D4558",
    x"BF3D4993",
    x"BF3D4DCE",
    x"BF3D5209",
    x"BF3D5644",
    x"BF3D5A7E",
    x"BF3D5EB9",
    x"BF3D62F3",
    x"BF3D672D",
    x"BF3D6B67",
    x"BF3D6FA1",
    x"BF3D73DB",
    x"BF3D7815",
    x"BF3D7C4E",
    x"BF3D8088",
    x"BF3D84C1",
    x"BF3D88FB",
    x"BF3D8D34",
    x"BF3D916D",
    x"BF3D95A6",
    x"BF3D99DF",
    x"BF3D9E17",
    x"BF3DA250",
    x"BF3DA688",
    x"BF3DAAC1",
    x"BF3DAEF9",
    x"BF3DB331",
    x"BF3DB769",
    x"BF3DBBA1",
    x"BF3DBFD9",
    x"BF3DC411",
    x"BF3DC848",
    x"BF3DCC80",
    x"BF3DD0B7",
    x"BF3DD4EE",
    x"BF3DD925",
    x"BF3DDD5C",
    x"BF3DE193",
    x"BF3DE5CA",
    x"BF3DEA01",
    x"BF3DEE37",
    x"BF3DF26E",
    x"BF3DF6A4",
    x"BF3DFADA",
    x"BF3DFF10",
    x"BF3E0346",
    x"BF3E077C",
    x"BF3E0BB2",
    x"BF3E0FE7",
    x"BF3E141D",
    x"BF3E1852",
    x"BF3E1C88",
    x"BF3E20BD",
    x"BF3E24F2",
    x"BF3E2927",
    x"BF3E2D5C",
    x"BF3E3190",
    x"BF3E35C5",
    x"BF3E39F9",
    x"BF3E3E2E",
    x"BF3E4262",
    x"BF3E4696",
    x"BF3E4ACA",
    x"BF3E4EFE",
    x"BF3E5332",
    x"BF3E5766",
    x"BF3E5B99",
    x"BF3E5FCD",
    x"BF3E6400",
    x"BF3E6833",
    x"BF3E6C66",
    x"BF3E7099",
    x"BF3E74CC",
    x"BF3E78FF",
    x"BF3E7D31",
    x"BF3E8164",
    x"BF3E8596",
    x"BF3E89C9",
    x"BF3E8DFB",
    x"BF3E922D",
    x"BF3E965F",
    x"BF3E9A91",
    x"BF3E9EC3",
    x"BF3EA2F4",
    x"BF3EA726",
    x"BF3EAB57",
    x"BF3EAF88",
    x"BF3EB3B9",
    x"BF3EB7EA",
    x"BF3EBC1B",
    x"BF3EC04C",
    x"BF3EC47D",
    x"BF3EC8AD",
    x"BF3ECCDE",
    x"BF3ED10E",
    x"BF3ED53F",
    x"BF3ED96F",
    x"BF3EDD9F",
    x"BF3EE1CF",
    x"BF3EE5FE",
    x"BF3EEA2E",
    x"BF3EEE5E",
    x"BF3EF28D",
    x"BF3EF6BC",
    x"BF3EFAEB",
    x"BF3EFF1B",
    x"BF3F034A",
    x"BF3F0778",
    x"BF3F0BA7",
    x"BF3F0FD6",
    x"BF3F1404",
    x"BF3F1833",
    x"BF3F1C61",
    x"BF3F208F",
    x"BF3F24BD",
    x"BF3F28EB",
    x"BF3F2D19",
    x"BF3F3147",
    x"BF3F3574",
    x"BF3F39A2",
    x"BF3F3DCF",
    x"BF3F41FC",
    x"BF3F4629",
    x"BF3F4A56",
    x"BF3F4E83",
    x"BF3F52B0",
    x"BF3F56DD",
    x"BF3F5B09",
    x"BF3F5F36",
    x"BF3F6362",
    x"BF3F678E",
    x"BF3F6BBA",
    x"BF3F6FE6",
    x"BF3F7412",
    x"BF3F783E",
    x"BF3F7C6A",
    x"BF3F8095",
    x"BF3F84C0",
    x"BF3F88EC",
    x"BF3F8D17",
    x"BF3F9142",
    x"BF3F956D",
    x"BF3F9998",
    x"BF3F9DC2",
    x"BF3FA1ED",
    x"BF3FA617",
    x"BF3FAA42",
    x"BF3FAE6C",
    x"BF3FB296",
    x"BF3FB6C0",
    x"BF3FBAEA",
    x"BF3FBF14",
    x"BF3FC33E",
    x"BF3FC767",
    x"BF3FCB91",
    x"BF3FCFBA",
    x"BF3FD3E3",
    x"BF3FD80C",
    x"BF3FDC35",
    x"BF3FE05E",
    x"BF3FE487",
    x"BF3FE8AF",
    x"BF3FECD8",
    x"BF3FF100",
    x"BF3FF529",
    x"BF3FF951",
    x"BF3FFD79",
    x"BF4001A1",
    x"BF4005C8",
    x"BF4009F0",
    x"BF400E18",
    x"BF40123F",
    x"BF401667",
    x"BF401A8E",
    x"BF401EB5",
    x"BF4022DC",
    x"BF402703",
    x"BF402B2A",
    x"BF402F50",
    x"BF403377",
    x"BF40379D",
    x"BF403BC4",
    x"BF403FEA",
    x"BF404410",
    x"BF404836",
    x"BF404C5C",
    x"BF405081",
    x"BF4054A7",
    x"BF4058CD",
    x"BF405CF2",
    x"BF406117",
    x"BF40653C",
    x"BF406961",
    x"BF406D86",
    x"BF4071AB",
    x"BF4075D0",
    x"BF4079F4",
    x"BF407E19",
    x"BF40823D",
    x"BF408661",
    x"BF408A85",
    x"BF408EA9",
    x"BF4092CD",
    x"BF4096F1",
    x"BF409B15",
    x"BF409F38",
    x"BF40A35C",
    x"BF40A77F",
    x"BF40ABA2",
    x"BF40AFC5",
    x"BF40B3E8",
    x"BF40B80B",
    x"BF40BC2E",
    x"BF40C050",
    x"BF40C473",
    x"BF40C895",
    x"BF40CCB7",
    x"BF40D0DA",
    x"BF40D4FC",
    x"BF40D91E",
    x"BF40DD3F",
    x"BF40E161",
    x"BF40E583",
    x"BF40E9A4",
    x"BF40EDC5",
    x"BF40F1E7",
    x"BF40F608",
    x"BF40FA29",
    x"BF40FE49",
    x"BF41026A",
    x"BF41068B",
    x"BF410AAB",
    x"BF410ECC",
    x"BF4112EC",
    x"BF41170C",
    x"BF411B2C",
    x"BF411F4C",
    x"BF41236C",
    x"BF41278C",
    x"BF412BAB",
    x"BF412FCB",
    x"BF4133EA",
    x"BF413809",
    x"BF413C28",
    x"BF414047",
    x"BF414466",
    x"BF414885",
    x"BF414CA4",
    x"BF4150C2",
    x"BF4154E1",
    x"BF4158FF",
    x"BF415D1D",
    x"BF41613B",
    x"BF416559",
    x"BF416977",
    x"BF416D95",
    x"BF4171B2",
    x"BF4175D0",
    x"BF4179ED",
    x"BF417E0A",
    x"BF418228",
    x"BF418645",
    x"BF418A61",
    x"BF418E7E",
    x"BF41929B",
    x"BF4196B7",
    x"BF419AD4",
    x"BF419EF0",
    x"BF41A30C",
    x"BF41A728",
    x"BF41AB44",
    x"BF41AF60",
    x"BF41B37C",
    x"BF41B798",
    x"BF41BBB3",
    x"BF41BFCF",
    x"BF41C3EA",
    x"BF41C805",
    x"BF41CC20",
    x"BF41D03B",
    x"BF41D456",
    x"BF41D870",
    x"BF41DC8B",
    x"BF41E0A5",
    x"BF41E4C0",
    x"BF41E8DA",
    x"BF41ECF4",
    x"BF41F10E",
    x"BF41F528",
    x"BF41F942",
    x"BF41FD5B",
    x"BF420175",
    x"BF42058E",
    x"BF4209A7",
    x"BF420DC1",
    x"BF4211DA",
    x"BF4215F3",
    x"BF421A0B",
    x"BF421E24",
    x"BF42223D",
    x"BF422655",
    x"BF422A6E",
    x"BF422E86",
    x"BF42329E",
    x"BF4236B6",
    x"BF423ACE",
    x"BF423EE5",
    x"BF4242FD",
    x"BF424715",
    x"BF424B2C",
    x"BF424F43",
    x"BF42535B",
    x"BF425772",
    x"BF425B89",
    x"BF425F9F",
    x"BF4263B6",
    x"BF4267CD",
    x"BF426BE3",
    x"BF426FFA",
    x"BF427410",
    x"BF427826",
    x"BF427C3C",
    x"BF428052",
    x"BF428468",
    x"BF42887D",
    x"BF428C93",
    x"BF4290A8",
    x"BF4294BD",
    x"BF4298D3",
    x"BF429CE8",
    x"BF42A0FD",
    x"BF42A511",
    x"BF42A926",
    x"BF42AD3B",
    x"BF42B14F",
    x"BF42B564",
    x"BF42B978",
    x"BF42BD8C",
    x"BF42C1A0",
    x"BF42C5B4",
    x"BF42C9C8",
    x"BF42CDDB",
    x"BF42D1EF",
    x"BF42D602",
    x"BF42DA16",
    x"BF42DE29",
    x"BF42E23C",
    x"BF42E64F",
    x"BF42EA62",
    x"BF42EE74",
    x"BF42F287",
    x"BF42F69A",
    x"BF42FAAC",
    x"BF42FEBE",
    x"BF4302D0",
    x"BF4306E2",
    x"BF430AF4",
    x"BF430F06",
    x"BF431318",
    x"BF431729",
    x"BF431B3B",
    x"BF431F4C",
    x"BF43235D",
    x"BF43276E",
    x"BF432B7F",
    x"BF432F90",
    x"BF4333A1",
    x"BF4337B1",
    x"BF433BC2",
    x"BF433FD2",
    x"BF4343E2",
    x"BF4347F3",
    x"BF434C03",
    x"BF435012",
    x"BF435422",
    x"BF435832",
    x"BF435C41",
    x"BF436051",
    x"BF436460",
    x"BF43686F",
    x"BF436C7F",
    x"BF43708D",
    x"BF43749C",
    x"BF4378AB",
    x"BF437CBA",
    x"BF4380C8",
    x"BF4384D6",
    x"BF4388E5",
    x"BF438CF3",
    x"BF439101",
    x"BF43950F",
    x"BF43991D",
    x"BF439D2A",
    x"BF43A138",
    x"BF43A545",
    x"BF43A953",
    x"BF43AD60",
    x"BF43B16D",
    x"BF43B57A",
    x"BF43B987",
    x"BF43BD93",
    x"BF43C1A0",
    x"BF43C5AC",
    x"BF43C9B9",
    x"BF43CDC5",
    x"BF43D1D1",
    x"BF43D5DD",
    x"BF43D9E9",
    x"BF43DDF5",
    x"BF43E200",
    x"BF43E60C",
    x"BF43EA17",
    x"BF43EE23",
    x"BF43F22E",
    x"BF43F639",
    x"BF43FA44",
    x"BF43FE4F",
    x"BF44025A",
    x"BF440664",
    x"BF440A6F",
    x"BF440E79",
    x"BF441283",
    x"BF44168D",
    x"BF441A97",
    x"BF441EA1",
    x"BF4422AB",
    x"BF4426B5",
    x"BF442ABE",
    x"BF442EC8",
    x"BF4432D1",
    x"BF4436DA",
    x"BF443AE3",
    x"BF443EEC",
    x"BF4442F5",
    x"BF4446FE",
    x"BF444B06",
    x"BF444F0F",
    x"BF445317",
    x"BF44571F",
    x"BF445B27",
    x"BF445F2F",
    x"BF446337",
    x"BF44673F",
    x"BF446B47",
    x"BF446F4E",
    x"BF447356",
    x"BF44775D",
    x"BF447B64",
    x"BF447F6B",
    x"BF448372",
    x"BF448779",
    x"BF448B80",
    x"BF448F86",
    x"BF44938D",
    x"BF449793",
    x"BF449B99",
    x"BF449F9F",
    x"BF44A3A5",
    x"BF44A7AB",
    x"BF44ABB1",
    x"BF44AFB6",
    x"BF44B3BC",
    x"BF44B7C1",
    x"BF44BBC7",
    x"BF44BFCC",
    x"BF44C3D1",
    x"BF44C7D6",
    x"BF44CBDB",
    x"BF44CFDF",
    x"BF44D3E4",
    x"BF44D7E8",
    x"BF44DBED",
    x"BF44DFF1",
    x"BF44E3F5",
    x"BF44E7F9",
    x"BF44EBFD",
    x"BF44F000",
    x"BF44F404",
    x"BF44F807",
    x"BF44FC0B",
    x"BF45000E",
    x"BF450411",
    x"BF450814",
    x"BF450C17",
    x"BF45101A",
    x"BF45141D",
    x"BF45181F",
    x"BF451C22",
    x"BF452024",
    x"BF452426",
    x"BF452828",
    x"BF452C2A",
    x"BF45302C",
    x"BF45342E",
    x"BF45382F",
    x"BF453C31",
    x"BF454032",
    x"BF454433",
    x"BF454834",
    x"BF454C35",
    x"BF455036",
    x"BF455437",
    x"BF455838",
    x"BF455C38",
    x"BF456039",
    x"BF456439",
    x"BF456839",
    x"BF456C39",
    x"BF457039",
    x"BF457439",
    x"BF457839",
    x"BF457C38",
    x"BF458038",
    x"BF458437",
    x"BF458836",
    x"BF458C35",
    x"BF459034",
    x"BF459433",
    x"BF459832",
    x"BF459C31",
    x"BF45A02F",
    x"BF45A42D",
    x"BF45A82C",
    x"BF45AC2A",
    x"BF45B028",
    x"BF45B426",
    x"BF45B824",
    x"BF45BC21",
    x"BF45C01F",
    x"BF45C41C",
    x"BF45C819",
    x"BF45CC17",
    x"BF45D014",
    x"BF45D411",
    x"BF45D80E",
    x"BF45DC0A",
    x"BF45E007",
    x"BF45E403",
    x"BF45E800",
    x"BF45EBFC",
    x"BF45EFF8",
    x"BF45F3F4",
    x"BF45F7F0",
    x"BF45FBEC",
    x"BF45FFE7",
    x"BF4603E3",
    x"BF4607DE",
    x"BF460BDA",
    x"BF460FD5",
    x"BF4613D0",
    x"BF4617CB",
    x"BF461BC6",
    x"BF461FC0",
    x"BF4623BB",
    x"BF4627B5",
    x"BF462BB0",
    x"BF462FAA",
    x"BF4633A4",
    x"BF46379E",
    x"BF463B98",
    x"BF463F91",
    x"BF46438B",
    x"BF464785",
    x"BF464B7E",
    x"BF464F77",
    x"BF465370",
    x"BF465769",
    x"BF465B62",
    x"BF465F5B",
    x"BF466354",
    x"BF46674C",
    x"BF466B45",
    x"BF466F3D",
    x"BF467335",
    x"BF46772D",
    x"BF467B25",
    x"BF467F1D",
    x"BF468315",
    x"BF46870C",
    x"BF468B04",
    x"BF468EFB",
    x"BF4692F2",
    x"BF4696E9",
    x"BF469AE0",
    x"BF469ED7",
    x"BF46A2CE",
    x"BF46A6C5",
    x"BF46AABB",
    x"BF46AEB1",
    x"BF46B2A8",
    x"BF46B69E",
    x"BF46BA94",
    x"BF46BE8A",
    x"BF46C280",
    x"BF46C675",
    x"BF46CA6B",
    x"BF46CE60",
    x"BF46D256",
    x"BF46D64B",
    x"BF46DA40",
    x"BF46DE35",
    x"BF46E22A",
    x"BF46E61E",
    x"BF46EA13",
    x"BF46EE07",
    x"BF46F1FC",
    x"BF46F5F0",
    x"BF46F9E4",
    x"BF46FDD8",
    x"BF4701CC",
    x"BF4705C0",
    x"BF4709B3",
    x"BF470DA7",
    x"BF47119A",
    x"BF47158D",
    x"BF471981",
    x"BF471D74",
    x"BF472167",
    x"BF472559",
    x"BF47294C",
    x"BF472D3F",
    x"BF473131",
    x"BF473523",
    x"BF473916",
    x"BF473D08",
    x"BF4740FA",
    x"BF4744EB",
    x"BF4748DD",
    x"BF474CCF",
    x"BF4750C0",
    x"BF4754B2",
    x"BF4758A3",
    x"BF475C94",
    x"BF476085",
    x"BF476476",
    x"BF476866",
    x"BF476C57",
    x"BF477048",
    x"BF477438",
    x"BF477828",
    x"BF477C18",
    x"BF478008",
    x"BF4783F8",
    x"BF4787E8",
    x"BF478BD8",
    x"BF478FC7",
    x"BF4793B7",
    x"BF4797A6",
    x"BF479B95",
    x"BF479F84",
    x"BF47A373",
    x"BF47A762",
    x"BF47AB51",
    x"BF47AF3F",
    x"BF47B32E",
    x"BF47B71C",
    x"BF47BB0A",
    x"BF47BEF9",
    x"BF47C2E7",
    x"BF47C6D4",
    x"BF47CAC2",
    x"BF47CEB0",
    x"BF47D29D",
    x"BF47D68B",
    x"BF47DA78",
    x"BF47DE65",
    x"BF47E252",
    x"BF47E63F",
    x"BF47EA2C",
    x"BF47EE18",
    x"BF47F205",
    x"BF47F5F1",
    x"BF47F9DE",
    x"BF47FDCA",
    x"BF4801B6",
    x"BF4805A2",
    x"BF48098E",
    x"BF480D79",
    x"BF481165",
    x"BF481550",
    x"BF48193C",
    x"BF481D27",
    x"BF482112",
    x"BF4824FD",
    x"BF4828E8",
    x"BF482CD3",
    x"BF4830BD",
    x"BF4834A8",
    x"BF483892",
    x"BF483C7C",
    x"BF484067",
    x"BF484451",
    x"BF48483A",
    x"BF484C24",
    x"BF48500E",
    x"BF4853F7",
    x"BF4857E1",
    x"BF485BCA",
    x"BF485FB3",
    x"BF48639C",
    x"BF486785",
    x"BF486B6E",
    x"BF486F57",
    x"BF48733F",
    x"BF487728",
    x"BF487B10",
    x"BF487EF8",
    x"BF4882E0",
    x"BF4886C8",
    x"BF488AB0",
    x"BF488E98",
    x"BF48927F",
    x"BF489667",
    x"BF489A4E",
    x"BF489E36",
    x"BF48A21D",
    x"BF48A604",
    x"BF48A9EA",
    x"BF48ADD1",
    x"BF48B1B8",
    x"BF48B59E",
    x"BF48B985",
    x"BF48BD6B",
    x"BF48C151",
    x"BF48C537",
    x"BF48C91D",
    x"BF48CD03",
    x"BF48D0E9",
    x"BF48D4CE",
    x"BF48D8B3",
    x"BF48DC99",
    x"BF48E07E",
    x"BF48E463",
    x"BF48E848",
    x"BF48EC2D",
    x"BF48F011",
    x"BF48F3F6",
    x"BF48F7DA",
    x"BF48FBBF",
    x"BF48FFA3",
    x"BF490387",
    x"BF49076B",
    x"BF490B4F",
    x"BF490F33",
    x"BF491316",
    x"BF4916FA",
    x"BF491ADD",
    x"BF491EC0",
    x"BF4922A3",
    x"BF492686",
    x"BF492A69",
    x"BF492E4C",
    x"BF49322F",
    x"BF493611",
    x"BF4939F4",
    x"BF493DD6",
    x"BF4941B8",
    x"BF49459A",
    x"BF49497C",
    x"BF494D5E",
    x"BF49513F",
    x"BF495521",
    x"BF495902",
    x"BF495CE4",
    x"BF4960C5",
    x"BF4964A6",
    x"BF496887",
    x"BF496C68",
    x"BF497048",
    x"BF497429",
    x"BF497809",
    x"BF497BEA",
    x"BF497FCA",
    x"BF4983AA",
    x"BF49878A",
    x"BF498B6A",
    x"BF498F4A",
    x"BF499329",
    x"BF499709",
    x"BF499AE8",
    x"BF499EC7",
    x"BF49A2A6",
    x"BF49A685",
    x"BF49AA64",
    x"BF49AE43",
    x"BF49B222",
    x"BF49B600",
    x"BF49B9DF",
    x"BF49BDBD",
    x"BF49C19B",
    x"BF49C579",
    x"BF49C957",
    x"BF49CD35",
    x"BF49D112",
    x"BF49D4F0",
    x"BF49D8CD",
    x"BF49DCAB",
    x"BF49E088",
    x"BF49E465",
    x"BF49E842",
    x"BF49EC1F",
    x"BF49EFFB",
    x"BF49F3D8",
    x"BF49F7B4",
    x"BF49FB91",
    x"BF49FF6D",
    x"BF4A0349",
    x"BF4A0725",
    x"BF4A0B01",
    x"BF4A0EDC",
    x"BF4A12B8",
    x"BF4A1693",
    x"BF4A1A6F",
    x"BF4A1E4A",
    x"BF4A2225",
    x"BF4A2600",
    x"BF4A29DB",
    x"BF4A2DB6",
    x"BF4A3190",
    x"BF4A356B",
    x"BF4A3945",
    x"BF4A3D1F",
    x"BF4A40F9",
    x"BF4A44D3",
    x"BF4A48AD",
    x"BF4A4C87",
    x"BF4A5061",
    x"BF4A543A",
    x"BF4A5814",
    x"BF4A5BED",
    x"BF4A5FC6",
    x"BF4A639F",
    x"BF4A6778",
    x"BF4A6B51",
    x"BF4A6F29",
    x"BF4A7302",
    x"BF4A76DA",
    x"BF4A7AB3",
    x"BF4A7E8B",
    x"BF4A8263",
    x"BF4A863B",
    x"BF4A8A13",
    x"BF4A8DEA",
    x"BF4A91C2",
    x"BF4A9599",
    x"BF4A9971",
    x"BF4A9D48",
    x"BF4AA11F",
    x"BF4AA4F6",
    x"BF4AA8CD",
    x"BF4AACA4",
    x"BF4AB07A",
    x"BF4AB451",
    x"BF4AB827",
    x"BF4ABBFD",
    x"BF4ABFD3",
    x"BF4AC3A9",
    x"BF4AC77F",
    x"BF4ACB55",
    x"BF4ACF2A",
    x"BF4AD300",
    x"BF4AD6D5",
    x"BF4ADAAB",
    x"BF4ADE80",
    x"BF4AE255",
    x"BF4AE62A",
    x"BF4AE9FE",
    x"BF4AEDD3",
    x"BF4AF1A8",
    x"BF4AF57C",
    x"BF4AF950",
    x"BF4AFD24",
    x"BF4B00F8",
    x"BF4B04CC",
    x"BF4B08A0",
    x"BF4B0C74",
    x"BF4B1047",
    x"BF4B141B",
    x"BF4B17EE",
    x"BF4B1BC1",
    x"BF4B1F94",
    x"BF4B2367",
    x"BF4B273A",
    x"BF4B2B0D",
    x"BF4B2EDF",
    x"BF4B32B2",
    x"BF4B3684",
    x"BF4B3A56",
    x"BF4B3E28",
    x"BF4B41FA",
    x"BF4B45CC",
    x"BF4B499E",
    x"BF4B4D6F",
    x"BF4B5141",
    x"BF4B5512",
    x"BF4B58E3",
    x"BF4B5CB4",
    x"BF4B6085",
    x"BF4B6456",
    x"BF4B6827",
    x"BF4B6BF7",
    x"BF4B6FC8",
    x"BF4B7398",
    x"BF4B7768",
    x"BF4B7B39",
    x"BF4B7F09",
    x"BF4B82D8",
    x"BF4B86A8",
    x"BF4B8A78",
    x"BF4B8E47",
    x"BF4B9217",
    x"BF4B95E6",
    x"BF4B99B5",
    x"BF4B9D84",
    x"BF4BA153",
    x"BF4BA522",
    x"BF4BA8F0",
    x"BF4BACBF",
    x"BF4BB08D",
    x"BF4BB45B",
    x"BF4BB82A",
    x"BF4BBBF8",
    x"BF4BBFC6",
    x"BF4BC393",
    x"BF4BC761",
    x"BF4BCB2F",
    x"BF4BCEFC",
    x"BF4BD2C9",
    x"BF4BD696",
    x"BF4BDA63",
    x"BF4BDE30",
    x"BF4BE1FD",
    x"BF4BE5CA",
    x"BF4BE996",
    x"BF4BED63",
    x"BF4BF12F",
    x"BF4BF4FB",
    x"BF4BF8C7",
    x"BF4BFC93",
    x"BF4C005F",
    x"BF4C042B",
    x"BF4C07F6",
    x"BF4C0BC2",
    x"BF4C0F8D",
    x"BF4C1358",
    x"BF4C1723",
    x"BF4C1AEE",
    x"BF4C1EB9",
    x"BF4C2284",
    x"BF4C264E",
    x"BF4C2A19",
    x"BF4C2DE3",
    x"BF4C31AD",
    x"BF4C3578",
    x"BF4C3942",
    x"BF4C3D0B",
    x"BF4C40D5",
    x"BF4C449F",
    x"BF4C4868",
    x"BF4C4C32",
    x"BF4C4FFB",
    x"BF4C53C4",
    x"BF4C578D",
    x"BF4C5B56",
    x"BF4C5F1E",
    x"BF4C62E7",
    x"BF4C66B0",
    x"BF4C6A78",
    x"BF4C6E40",
    x"BF4C7208",
    x"BF4C75D0",
    x"BF4C7998",
    x"BF4C7D60",
    x"BF4C8128",
    x"BF4C84EF",
    x"BF4C88B6",
    x"BF4C8C7E",
    x"BF4C9045",
    x"BF4C940C",
    x"BF4C97D3",
    x"BF4C9B99",
    x"BF4C9F60",
    x"BF4CA327",
    x"BF4CA6ED",
    x"BF4CAAB3",
    x"BF4CAE79",
    x"BF4CB23F",
    x"BF4CB605",
    x"BF4CB9CB",
    x"BF4CBD91",
    x"BF4CC156",
    x"BF4CC51C",
    x"BF4CC8E1",
    x"BF4CCCA6",
    x"BF4CD06B",
    x"BF4CD430",
    x"BF4CD7F5",
    x"BF4CDBBA",
    x"BF4CDF7E",
    x"BF4CE343",
    x"BF4CE707",
    x"BF4CEACB",
    x"BF4CEE8F",
    x"BF4CF253",
    x"BF4CF617",
    x"BF4CF9DB",
    x"BF4CFD9E",
    x"BF4D0162",
    x"BF4D0525",
    x"BF4D08E8",
    x"BF4D0CAB",
    x"BF4D106E",
    x"BF4D1431",
    x"BF4D17F4",
    x"BF4D1BB6",
    x"BF4D1F79",
    x"BF4D233B",
    x"BF4D26FD",
    x"BF4D2ABF",
    x"BF4D2E81",
    x"BF4D3243",
    x"BF4D3605",
    x"BF4D39C6",
    x"BF4D3D88",
    x"BF4D4149",
    x"BF4D450A",
    x"BF4D48CB",
    x"BF4D4C8C",
    x"BF4D504D",
    x"BF4D540E",
    x"BF4D57CE",
    x"BF4D5B8F",
    x"BF4D5F4F",
    x"BF4D6310",
    x"BF4D66D0",
    x"BF4D6A90",
    x"BF4D6E4F",
    x"BF4D720F",
    x"BF4D75CF",
    x"BF4D798E",
    x"BF4D7D4E",
    x"BF4D810D",
    x"BF4D84CC",
    x"BF4D888B",
    x"BF4D8C4A",
    x"BF4D9009",
    x"BF4D93C7",
    x"BF4D9786",
    x"BF4D9B44",
    x"BF4D9F02",
    x"BF4DA2C0",
    x"BF4DA67E",
    x"BF4DAA3C",
    x"BF4DADFA",
    x"BF4DB1B8",
    x"BF4DB575",
    x"BF4DB932",
    x"BF4DBCF0",
    x"BF4DC0AD",
    x"BF4DC46A",
    x"BF4DC827",
    x"BF4DCBE3",
    x"BF4DCFA0",
    x"BF4DD35D",
    x"BF4DD719",
    x"BF4DDAD5",
    x"BF4DDE91",
    x"BF4DE24D",
    x"BF4DE609",
    x"BF4DE9C5",
    x"BF4DED81",
    x"BF4DF13C",
    x"BF4DF4F8",
    x"BF4DF8B3",
    x"BF4DFC6E",
    x"BF4E0029",
    x"BF4E03E4",
    x"BF4E079F",
    x"BF4E0B59",
    x"BF4E0F14",
    x"BF4E12CE",
    x"BF4E1689",
    x"BF4E1A43",
    x"BF4E1DFD",
    x"BF4E21B7",
    x"BF4E2570",
    x"BF4E292A",
    x"BF4E2CE4",
    x"BF4E309D",
    x"BF4E3456",
    x"BF4E380F",
    x"BF4E3BC8",
    x"BF4E3F81",
    x"BF4E433A",
    x"BF4E46F3",
    x"BF4E4AAB",
    x"BF4E4E64",
    x"BF4E521C",
    x"BF4E55D4",
    x"BF4E598C",
    x"BF4E5D44",
    x"BF4E60FC",
    x"BF4E64B4",
    x"BF4E686B",
    x"BF4E6C23",
    x"BF4E6FDA",
    x"BF4E7391",
    x"BF4E7748",
    x"BF4E7AFF",
    x"BF4E7EB6",
    x"BF4E826C",
    x"BF4E8623",
    x"BF4E89D9",
    x"BF4E8D90",
    x"BF4E9146",
    x"BF4E94FC",
    x"BF4E98B2",
    x"BF4E9C68",
    x"BF4EA01D",
    x"BF4EA3D3",
    x"BF4EA788",
    x"BF4EAB3E",
    x"BF4EAEF3",
    x"BF4EB2A8",
    x"BF4EB65D",
    x"BF4EBA12",
    x"BF4EBDC6",
    x"BF4EC17B",
    x"BF4EC52F",
    x"BF4EC8E4",
    x"BF4ECC98",
    x"BF4ED04C",
    x"BF4ED400",
    x"BF4ED7B3",
    x"BF4EDB67",
    x"BF4EDF1B",
    x"BF4EE2CE",
    x"BF4EE681",
    x"BF4EEA35",
    x"BF4EEDE8",
    x"BF4EF19B",
    x"BF4EF54D",
    x"BF4EF900",
    x"BF4EFCB3",
    x"BF4F0065",
    x"BF4F0417",
    x"BF4F07CA",
    x"BF4F0B7C",
    x"BF4F0F2E",
    x"BF4F12DF",
    x"BF4F1691",
    x"BF4F1A43",
    x"BF4F1DF4",
    x"BF4F21A5",
    x"BF4F2557",
    x"BF4F2908",
    x"BF4F2CB9",
    x"BF4F3069",
    x"BF4F341A",
    x"BF4F37CB",
    x"BF4F3B7B",
    x"BF4F3F2B",
    x"BF4F42DC",
    x"BF4F468C",
    x"BF4F4A3C",
    x"BF4F4DEB",
    x"BF4F519B",
    x"BF4F554B",
    x"BF4F58FA",
    x"BF4F5CA9",
    x"BF4F6059",
    x"BF4F6408",
    x"BF4F67B7",
    x"BF4F6B65",
    x"BF4F6F14",
    x"BF4F72C3",
    x"BF4F7671",
    x"BF4F7A1F",
    x"BF4F7DCE",
    x"BF4F817C",
    x"BF4F852A",
    x"BF4F88D7",
    x"BF4F8C85",
    x"BF4F9033",
    x"BF4F93E0",
    x"BF4F978D",
    x"BF4F9B3B",
    x"BF4F9EE8",
    x"BF4FA295",
    x"BF4FA642",
    x"BF4FA9EE",
    x"BF4FAD9B",
    x"BF4FB147",
    x"BF4FB4F4",
    x"BF4FB8A0",
    x"BF4FBC4C",
    x"BF4FBFF8",
    x"BF4FC3A4",
    x"BF4FC74F",
    x"BF4FCAFB",
    x"BF4FCEA6",
    x"BF4FD252",
    x"BF4FD5FD",
    x"BF4FD9A8",
    x"BF4FDD53",
    x"BF4FE0FE",
    x"BF4FE4A8",
    x"BF4FE853",
    x"BF4FEBFD",
    x"BF4FEFA8",
    x"BF4FF352",
    x"BF4FF6FC",
    x"BF4FFAA6",
    x"BF4FFE50",
    x"BF5001F9",
    x"BF5005A3",
    x"BF50094C",
    x"BF500CF6",
    x"BF50109F",
    x"BF501448",
    x"BF5017F1",
    x"BF501B9A",
    x"BF501F42",
    x"BF5022EB",
    x"BF502693",
    x"BF502A3B",
    x"BF502DE4",
    x"BF50318C",
    x"BF503534",
    x"BF5038DB",
    x"BF503C83",
    x"BF50402B",
    x"BF5043D2",
    x"BF504779",
    x"BF504B21",
    x"BF504EC8",
    x"BF50526F",
    x"BF505615",
    x"BF5059BC",
    x"BF505D63",
    x"BF506109",
    x"BF5064AF",
    x"BF506856",
    x"BF506BFC",
    x"BF506FA1",
    x"BF507347",
    x"BF5076ED",
    x"BF507A92",
    x"BF507E38",
    x"BF5081DD",
    x"BF508582",
    x"BF508927",
    x"BF508CCC",
    x"BF509071",
    x"BF509416",
    x"BF5097BA",
    x"BF509B5F",
    x"BF509F03",
    x"BF50A2A7",
    x"BF50A64B",
    x"BF50A9EF",
    x"BF50AD93",
    x"BF50B137",
    x"BF50B4DA",
    x"BF50B87E",
    x"BF50BC21",
    x"BF50BFC4",
    x"BF50C367",
    x"BF50C70A",
    x"BF50CAAD",
    x"BF50CE4F",
    x"BF50D1F2",
    x"BF50D594",
    x"BF50D937",
    x"BF50DCD9",
    x"BF50E07B",
    x"BF50E41D",
    x"BF50E7BE",
    x"BF50EB60",
    x"BF50EF02",
    x"BF50F2A3",
    x"BF50F644",
    x"BF50F9E5",
    x"BF50FD86",
    x"BF510127",
    x"BF5104C8",
    x"BF510869",
    x"BF510C09",
    x"BF510FAA",
    x"BF51134A",
    x"BF5116EA",
    x"BF511A8A",
    x"BF511E2A",
    x"BF5121CA",
    x"BF512569",
    x"BF512909",
    x"BF512CA8",
    x"BF513047",
    x"BF5133E7",
    x"BF513786",
    x"BF513B25",
    x"BF513EC3",
    x"BF514262",
    x"BF514600",
    x"BF51499F",
    x"BF514D3D",
    x"BF5150DB",
    x"BF515479",
    x"BF515817",
    x"BF515BB5",
    x"BF515F52",
    x"BF5162F0",
    x"BF51668D",
    x"BF516A2A",
    x"BF516DC8",
    x"BF517165",
    x"BF517501",
    x"BF51789E",
    x"BF517C3B",
    x"BF517FD7",
    x"BF518374",
    x"BF518710",
    x"BF518AAC",
    x"BF518E48",
    x"BF5191E4",
    x"BF51957F",
    x"BF51991B",
    x"BF519CB7",
    x"BF51A052",
    x"BF51A3ED",
    x"BF51A788",
    x"BF51AB23",
    x"BF51AEBE",
    x"BF51B259",
    x"BF51B5F3",
    x"BF51B98E",
    x"BF51BD28",
    x"BF51C0C2",
    x"BF51C45C",
    x"BF51C7F6",
    x"BF51CB90",
    x"BF51CF2A",
    x"BF51D2C3",
    x"BF51D65D",
    x"BF51D9F6",
    x"BF51DD8F",
    x"BF51E129",
    x"BF51E4C1",
    x"BF51E85A",
    x"BF51EBF3",
    x"BF51EF8C",
    x"BF51F324",
    x"BF51F6BC",
    x"BF51FA54",
    x"BF51FDED",
    x"BF520184",
    x"BF52051C",
    x"BF5208B4",
    x"BF520C4C",
    x"BF520FE3",
    x"BF52137A",
    x"BF521711",
    x"BF521AA8",
    x"BF521E3F",
    x"BF5221D6",
    x"BF52256D",
    x"BF522903",
    x"BF522C9A",
    x"BF523030",
    x"BF5233C6",
    x"BF52375C",
    x"BF523AF2",
    x"BF523E88",
    x"BF52421E",
    x"BF5245B3",
    x"BF524949",
    x"BF524CDE",
    x"BF525073",
    x"BF525408",
    x"BF52579D",
    x"BF525B32",
    x"BF525EC6",
    x"BF52625B",
    x"BF5265EF",
    x"BF526983",
    x"BF526D18",
    x"BF5270AC",
    x"BF52743F",
    x"BF5277D3",
    x"BF527B67",
    x"BF527EFA",
    x"BF52828E",
    x"BF528621",
    x"BF5289B4",
    x"BF528D47",
    x"BF5290DA",
    x"BF52946D",
    x"BF5297FF",
    x"BF529B92",
    x"BF529F24",
    x"BF52A2B6",
    x"BF52A649",
    x"BF52A9DA",
    x"BF52AD6C",
    x"BF52B0FE",
    x"BF52B490",
    x"BF52B821",
    x"BF52BBB2",
    x"BF52BF44",
    x"BF52C2D5",
    x"BF52C666",
    x"BF52C9F7",
    x"BF52CD87",
    x"BF52D118",
    x"BF52D4A8",
    x"BF52D839",
    x"BF52DBC9",
    x"BF52DF59",
    x"BF52E2E9",
    x"BF52E679",
    x"BF52EA08",
    x"BF52ED98",
    x"BF52F127",
    x"BF52F4B7",
    x"BF52F846",
    x"BF52FBD5",
    x"BF52FF64",
    x"BF5302F3",
    x"BF530681",
    x"BF530A10",
    x"BF530D9E",
    x"BF53112D",
    x"BF5314BB",
    x"BF531849",
    x"BF531BD7",
    x"BF531F65",
    x"BF5322F2",
    x"BF532680",
    x"BF532A0D",
    x"BF532D9A",
    x"BF533128",
    x"BF5334B5",
    x"BF533841",
    x"BF533BCE",
    x"BF533F5B",
    x"BF5342E7",
    x"BF534674",
    x"BF534A00",
    x"BF534D8C",
    x"BF535118",
    x"BF5354A4",
    x"BF535830",
    x"BF535BBB",
    x"BF535F47",
    x"BF5362D2",
    x"BF53665E",
    x"BF5369E9",
    x"BF536D74",
    x"BF5370FF",
    x"BF537489",
    x"BF537814",
    x"BF537B9E",
    x"BF537F29",
    x"BF5382B3",
    x"BF53863D",
    x"BF5389C7",
    x"BF538D51",
    x"BF5390DB",
    x"BF539464",
    x"BF5397EE",
    x"BF539B77",
    x"BF539F00",
    x"BF53A289",
    x"BF53A612",
    x"BF53A99B",
    x"BF53AD24",
    x"BF53B0AC",
    x"BF53B435",
    x"BF53B7BD",
    x"BF53BB45",
    x"BF53BECD",
    x"BF53C255",
    x"BF53C5DD",
    x"BF53C965",
    x"BF53CCEC",
    x"BF53D074",
    x"BF53D3FB",
    x"BF53D782",
    x"BF53DB09",
    x"BF53DE90",
    x"BF53E217",
    x"BF53E59D",
    x"BF53E924",
    x"BF53ECAA",
    x"BF53F031",
    x"BF53F3B7",
    x"BF53F73D",
    x"BF53FAC3",
    x"BF53FE48",
    x"BF5401CE",
    x"BF540553",
    x"BF5408D9",
    x"BF540C5E",
    x"BF540FE3",
    x"BF541368",
    x"BF5416ED",
    x"BF541A72",
    x"BF541DF6",
    x"BF54217B",
    x"BF5424FF",
    x"BF542883",
    x"BF542C08",
    x"BF542F8C",
    x"BF54330F",
    x"BF543693",
    x"BF543A17",
    x"BF543D9A",
    x"BF54411D",
    x"BF5444A1",
    x"BF544824",
    x"BF544BA7",
    x"BF544F2A",
    x"BF5452AC",
    x"BF54562F",
    x"BF5459B1",
    x"BF545D33",
    x"BF5460B6",
    x"BF546438",
    x"BF5467BA",
    x"BF546B3B",
    x"BF546EBD",
    x"BF54723F",
    x"BF5475C0",
    x"BF547941",
    x"BF547CC3",
    x"BF548044",
    x"BF5483C4",
    x"BF548745",
    x"BF548AC6",
    x"BF548E46",
    x"BF5491C7",
    x"BF549547",
    x"BF5498C7",
    x"BF549C47",
    x"BF549FC7",
    x"BF54A347",
    x"BF54A6C6",
    x"BF54AA46",
    x"BF54ADC5",
    x"BF54B144",
    x"BF54B4C4",
    x"BF54B843",
    x"BF54BBC1",
    x"BF54BF40",
    x"BF54C2BF",
    x"BF54C63D",
    x"BF54C9BC",
    x"BF54CD3A",
    x"BF54D0B8",
    x"BF54D436",
    x"BF54D7B4",
    x"BF54DB31",
    x"BF54DEAF",
    x"BF54E22C",
    x"BF54E5AA",
    x"BF54E927",
    x"BF54ECA4",
    x"BF54F021",
    x"BF54F39E",
    x"BF54F71A",
    x"BF54FA97",
    x"BF54FE13",
    x"BF55018F",
    x"BF55050C",
    x"BF550888",
    x"BF550C04",
    x"BF550F7F",
    x"BF5512FB",
    x"BF551676",
    x"BF5519F2",
    x"BF551D6D",
    x"BF5520E8",
    x"BF552463",
    x"BF5527DE",
    x"BF552B59",
    x"BF552ED4",
    x"BF55324E",
    x"BF5535C8",
    x"BF553943",
    x"BF553CBD",
    x"BF554037",
    x"BF5543B1",
    x"BF55472A",
    x"BF554AA4",
    x"BF554E1D",
    x"BF555197",
    x"BF555510",
    x"BF555889",
    x"BF555C02",
    x"BF555F7B",
    x"BF5562F3",
    x"BF55666C",
    x"BF5569E4",
    x"BF556D5D",
    x"BF5570D5",
    x"BF55744D",
    x"BF5577C5",
    x"BF557B3D",
    x"BF557EB4",
    x"BF55822C",
    x"BF5585A3",
    x"BF55891A",
    x"BF558C92",
    x"BF559009",
    x"BF55937F",
    x"BF5596F6",
    x"BF559A6D",
    x"BF559DE3",
    x"BF55A15A",
    x"BF55A4D0",
    x"BF55A846",
    x"BF55ABBC",
    x"BF55AF32",
    x"BF55B2A8",
    x"BF55B61D",
    x"BF55B993",
    x"BF55BD08",
    x"BF55C07D",
    x"BF55C3F2",
    x"BF55C767",
    x"BF55CADC",
    x"BF55CE51",
    x"BF55D1C5",
    x"BF55D53A",
    x"BF55D8AE",
    x"BF55DC22",
    x"BF55DF96",
    x"BF55E30A",
    x"BF55E67E",
    x"BF55E9F2",
    x"BF55ED65",
    x"BF55F0D9",
    x"BF55F44C",
    x"BF55F7BF",
    x"BF55FB32",
    x"BF55FEA5",
    x"BF560218",
    x"BF56058B",
    x"BF5608FD",
    x"BF560C70",
    x"BF560FE2",
    x"BF561354",
    x"BF5616C6",
    x"BF561A38",
    x"BF561DA9",
    x"BF56211B",
    x"BF56248D",
    x"BF5627FE",
    x"BF562B6F",
    x"BF562EE0",
    x"BF563251",
    x"BF5635C2",
    x"BF563933",
    x"BF563CA3",
    x"BF564014",
    x"BF564384",
    x"BF5646F4",
    x"BF564A64",
    x"BF564DD4",
    x"BF565144",
    x"BF5654B4",
    x"BF565823",
    x"BF565B93",
    x"BF565F02",
    x"BF566271",
    x"BF5665E0",
    x"BF56694F",
    x"BF566CBE",
    x"BF56702C",
    x"BF56739B",
    x"BF567709",
    x"BF567A78",
    x"BF567DE6",
    x"BF568154",
    x"BF5684C2",
    x"BF56882F",
    x"BF568B9D",
    x"BF568F0A",
    x"BF569278",
    x"BF5695E5",
    x"BF569952",
    x"BF569CBF",
    x"BF56A02C",
    x"BF56A399",
    x"BF56A705",
    x"BF56AA72",
    x"BF56ADDE",
    x"BF56B14A",
    x"BF56B4B6",
    x"BF56B822",
    x"BF56BB8E",
    x"BF56BEF9",
    x"BF56C265",
    x"BF56C5D0",
    x"BF56C93C",
    x"BF56CCA7",
    x"BF56D012",
    x"BF56D37D",
    x"BF56D6E8",
    x"BF56DA52",
    x"BF56DDBD",
    x"BF56E127",
    x"BF56E491",
    x"BF56E7FB",
    x"BF56EB65",
    x"BF56EECF",
    x"BF56F239",
    x"BF56F5A3",
    x"BF56F90C",
    x"BF56FC75",
    x"BF56FFDF",
    x"BF570348",
    x"BF5706B1",
    x"BF570A19",
    x"BF570D82",
    x"BF5710EB",
    x"BF571453",
    x"BF5717BB",
    x"BF571B24",
    x"BF571E8C",
    x"BF5721F3",
    x"BF57255B",
    x"BF5728C3",
    x"BF572C2A",
    x"BF572F92",
    x"BF5732F9",
    x"BF573660",
    x"BF5739C7",
    x"BF573D2E",
    x"BF574095",
    x"BF5743FB",
    x"BF574762",
    x"BF574AC8",
    x"BF574E2F",
    x"BF575195",
    x"BF5754FB",
    x"BF575860",
    x"BF575BC6",
    x"BF575F2C",
    x"BF576291",
    x"BF5765F6",
    x"BF57695C",
    x"BF576CC1",
    x"BF577026",
    x"BF57738A",
    x"BF5776EF",
    x"BF577A54",
    x"BF577DB8",
    x"BF57811C",
    x"BF578480",
    x"BF5787E4",
    x"BF578B48",
    x"BF578EAC",
    x"BF579210",
    x"BF579573",
    x"BF5798D7",
    x"BF579C3A",
    x"BF579F9D",
    x"BF57A300",
    x"BF57A663",
    x"BF57A9C6",
    x"BF57AD28",
    x"BF57B08B",
    x"BF57B3ED",
    x"BF57B74F",
    x"BF57BAB1",
    x"BF57BE13",
    x"BF57C175",
    x"BF57C4D7",
    x"BF57C838",
    x"BF57CB9A",
    x"BF57CEFB",
    x"BF57D25C",
    x"BF57D5BD",
    x"BF57D91E",
    x"BF57DC7F",
    x"BF57DFDF",
    x"BF57E340",
    x"BF57E6A0",
    x"BF57EA01",
    x"BF57ED61",
    x"BF57F0C1",
    x"BF57F421",
    x"BF57F780",
    x"BF57FAE0",
    x"BF57FE3F",
    x"BF58019F",
    x"BF5804FE",
    x"BF58085D",
    x"BF580BBC",
    x"BF580F1B",
    x"BF581279",
    x"BF5815D8",
    x"BF581936",
    x"BF581C95",
    x"BF581FF3",
    x"BF582351",
    x"BF5826AF",
    x"BF582A0D",
    x"BF582D6A",
    x"BF5830C8",
    x"BF583425",
    x"BF583782",
    x"BF583AE0",
    x"BF583E3D",
    x"BF584199",
    x"BF5844F6",
    x"BF584853",
    x"BF584BAF",
    x"BF584F0C",
    x"BF585268",
    x"BF5855C4",
    x"BF585920",
    x"BF585C7C",
    x"BF585FD7",
    x"BF586333",
    x"BF58668E",
    x"BF5869EA",
    x"BF586D45",
    x"BF5870A0",
    x"BF5873FB",
    x"BF587756",
    x"BF587AB0",
    x"BF587E0B",
    x"BF588165",
    x"BF5884BF",
    x"BF58881A",
    x"BF588B74",
    x"BF588ECD",
    x"BF589227",
    x"BF589581",
    x"BF5898DA",
    x"BF589C34",
    x"BF589F8D",
    x"BF58A2E6",
    x"BF58A63F",
    x"BF58A998",
    x"BF58ACF0",
    x"BF58B049",
    x"BF58B3A1",
    x"BF58B6FA",
    x"BF58BA52",
    x"BF58BDAA",
    x"BF58C102",
    x"BF58C45A",
    x"BF58C7B1",
    x"BF58CB09",
    x"BF58CE60",
    x"BF58D1B7",
    x"BF58D50E",
    x"BF58D865",
    x"BF58DBBC",
    x"BF58DF13",
    x"BF58E26A",
    x"BF58E5C0",
    x"BF58E916",
    x"BF58EC6D",
    x"BF58EFC3",
    x"BF58F319",
    x"BF58F66F",
    x"BF58F9C4",
    x"BF58FD1A",
    x"BF59006F",
    x"BF5903C5",
    x"BF59071A",
    x"BF590A6F",
    x"BF590DC4",
    x"BF591118",
    x"BF59146D",
    x"BF5917C2",
    x"BF591B16",
    x"BF591E6A",
    x"BF5921BE",
    x"BF592512",
    x"BF592866",
    x"BF592BBA",
    x"BF592F0E",
    x"BF593261",
    x"BF5935B4",
    x"BF593908",
    x"BF593C5B",
    x"BF593FAE",
    x"BF594300",
    x"BF594653",
    x"BF5949A6",
    x"BF594CF8",
    x"BF59504A",
    x"BF59539C",
    x"BF5956EE",
    x"BF595A40",
    x"BF595D92",
    x"BF5960E4",
    x"BF596435",
    x"BF596787",
    x"BF596AD8",
    x"BF596E29",
    x"BF59717A",
    x"BF5974CB",
    x"BF59781C",
    x"BF597B6C",
    x"BF597EBD",
    x"BF59820D",
    x"BF59855D",
    x"BF5988AD",
    x"BF598BFD",
    x"BF598F4D",
    x"BF59929D",
    x"BF5995EC",
    x"BF59993C",
    x"BF599C8B",
    x"BF599FDA",
    x"BF59A329",
    x"BF59A678",
    x"BF59A9C7",
    x"BF59AD15",
    x"BF59B064",
    x"BF59B3B2",
    x"BF59B700",
    x"BF59BA4E",
    x"BF59BD9C",
    x"BF59C0EA",
    x"BF59C438",
    x"BF59C785",
    x"BF59CAD3",
    x"BF59CE20",
    x"BF59D16D",
    x"BF59D4BA",
    x"BF59D807",
    x"BF59DB54",
    x"BF59DEA1",
    x"BF59E1ED",
    x"BF59E53A",
    x"BF59E886",
    x"BF59EBD2",
    x"BF59EF1E",
    x"BF59F26A",
    x"BF59F5B6",
    x"BF59F901",
    x"BF59FC4D",
    x"BF59FF98",
    x"BF5A02E3",
    x"BF5A062E",
    x"BF5A0979",
    x"BF5A0CC4",
    x"BF5A100F",
    x"BF5A1359",
    x"BF5A16A4",
    x"BF5A19EE",
    x"BF5A1D38",
    x"BF5A2082",
    x"BF5A23CC",
    x"BF5A2716",
    x"BF5A2A60",
    x"BF5A2DA9",
    x"BF5A30F2",
    x"BF5A343C",
    x"BF5A3785",
    x"BF5A3ACE",
    x"BF5A3E17",
    x"BF5A415F",
    x"BF5A44A8",
    x"BF5A47F0",
    x"BF5A4B39",
    x"BF5A4E81",
    x"BF5A51C9",
    x"BF5A5511",
    x"BF5A5859",
    x"BF5A5BA0",
    x"BF5A5EE8",
    x"BF5A622F",
    x"BF5A6577",
    x"BF5A68BE",
    x"BF5A6C05",
    x"BF5A6F4C",
    x"BF5A7292",
    x"BF5A75D9",
    x"BF5A791F",
    x"BF5A7C66",
    x"BF5A7FAC",
    x"BF5A82F2",
    x"BF5A8638",
    x"BF5A897E",
    x"BF5A8CC3",
    x"BF5A9009",
    x"BF5A934E",
    x"BF5A9694",
    x"BF5A99D9",
    x"BF5A9D1E",
    x"BF5AA063",
    x"BF5AA3A8",
    x"BF5AA6EC",
    x"BF5AAA31",
    x"BF5AAD75",
    x"BF5AB0B9",
    x"BF5AB3FD",
    x"BF5AB741",
    x"BF5ABA85",
    x"BF5ABDC9",
    x"BF5AC10D",
    x"BF5AC450",
    x"BF5AC793",
    x"BF5ACAD6",
    x"BF5ACE1A",
    x"BF5AD15C",
    x"BF5AD49F",
    x"BF5AD7E2",
    x"BF5ADB24",
    x"BF5ADE67",
    x"BF5AE1A9",
    x"BF5AE4EB",
    x"BF5AE82D",
    x"BF5AEB6F",
    x"BF5AEEB1",
    x"BF5AF1F2",
    x"BF5AF534",
    x"BF5AF875",
    x"BF5AFBB6",
    x"BF5AFEF7",
    x"BF5B0238",
    x"BF5B0579",
    x"BF5B08BA",
    x"BF5B0BFA",
    x"BF5B0F3B",
    x"BF5B127B",
    x"BF5B15BB",
    x"BF5B18FB",
    x"BF5B1C3B",
    x"BF5B1F7B",
    x"BF5B22BB",
    x"BF5B25FA",
    x"BF5B2939",
    x"BF5B2C79",
    x"BF5B2FB8",
    x"BF5B32F7",
    x"BF5B3636",
    x"BF5B3974",
    x"BF5B3CB3",
    x"BF5B3FF1",
    x"BF5B4330",
    x"BF5B466E",
    x"BF5B49AC",
    x"BF5B4CEA",
    x"BF5B5027",
    x"BF5B5365",
    x"BF5B56A3",
    x"BF5B59E0",
    x"BF5B5D1D",
    x"BF5B605A",
    x"BF5B6397",
    x"BF5B66D4",
    x"BF5B6A11",
    x"BF5B6D4D",
    x"BF5B708A",
    x"BF5B73C6",
    x"BF5B7702",
    x"BF5B7A3E",
    x"BF5B7D7A",
    x"BF5B80B6",
    x"BF5B83F2",
    x"BF5B872D",
    x"BF5B8A69",
    x"BF5B8DA4",
    x"BF5B90DF",
    x"BF5B941A",
    x"BF5B9755",
    x"BF5B9A90",
    x"BF5B9DCA",
    x"BF5BA105",
    x"BF5BA43F",
    x"BF5BA779",
    x"BF5BAAB3",
    x"BF5BADED",
    x"BF5BB127",
    x"BF5BB461",
    x"BF5BB79A",
    x"BF5BBAD4",
    x"BF5BBE0D",
    x"BF5BC146",
    x"BF5BC47F",
    x"BF5BC7B8",
    x"BF5BCAF1",
    x"BF5BCE29",
    x"BF5BD162",
    x"BF5BD49A",
    x"BF5BD7D3",
    x"BF5BDB0B",
    x"BF5BDE43",
    x"BF5BE17A",
    x"BF5BE4B2",
    x"BF5BE7EA",
    x"BF5BEB21",
    x"BF5BEE58",
    x"BF5BF190",
    x"BF5BF4C7",
    x"BF5BF7FD",
    x"BF5BFB34",
    x"BF5BFE6B",
    x"BF5C01A1",
    x"BF5C04D8",
    x"BF5C080E",
    x"BF5C0B44",
    x"BF5C0E7A",
    x"BF5C11B0",
    x"BF5C14E6",
    x"BF5C181B",
    x"BF5C1B51",
    x"BF5C1E86",
    x"BF5C21BB",
    x"BF5C24F0",
    x"BF5C2825",
    x"BF5C2B5A",
    x"BF5C2E8E",
    x"BF5C31C3",
    x"BF5C34F7",
    x"BF5C382B",
    x"BF5C3B60",
    x"BF5C3E94",
    x"BF5C41C7",
    x"BF5C44FB",
    x"BF5C482F",
    x"BF5C4B62",
    x"BF5C4E95",
    x"BF5C51C9",
    x"BF5C54FC",
    x"BF5C582F",
    x"BF5C5B61",
    x"BF5C5E94",
    x"BF5C61C7",
    x"BF5C64F9",
    x"BF5C682B",
    x"BF5C6B5D",
    x"BF5C6E8F",
    x"BF5C71C1",
    x"BF5C74F3",
    x"BF5C7824",
    x"BF5C7B56",
    x"BF5C7E87",
    x"BF5C81B8",
    x"BF5C84EA",
    x"BF5C881A",
    x"BF5C8B4B",
    x"BF5C8E7C",
    x"BF5C91AC",
    x"BF5C94DD",
    x"BF5C980D",
    x"BF5C9B3D",
    x"BF5C9E6D",
    x"BF5CA19D",
    x"BF5CA4CD",
    x"BF5CA7FC",
    x"BF5CAB2C",
    x"BF5CAE5B",
    x"BF5CB18A",
    x"BF5CB4B9",
    x"BF5CB7E8",
    x"BF5CBB17",
    x"BF5CBE46",
    x"BF5CC174",
    x"BF5CC4A3",
    x"BF5CC7D1",
    x"BF5CCAFF",
    x"BF5CCE2D",
    x"BF5CD15B",
    x"BF5CD489",
    x"BF5CD7B6",
    x"BF5CDAE4",
    x"BF5CDE11",
    x"BF5CE13E",
    x"BF5CE46B",
    x"BF5CE798",
    x"BF5CEAC5",
    x"BF5CEDF2",
    x"BF5CF11E",
    x"BF5CF44B",
    x"BF5CF777",
    x"BF5CFAA3",
    x"BF5CFDCF",
    x"BF5D00FB",
    x"BF5D0427",
    x"BF5D0752",
    x"BF5D0A7E",
    x"BF5D0DA9",
    x"BF5D10D4",
    x"BF5D13FF",
    x"BF5D172A",
    x"BF5D1A55",
    x"BF5D1D80",
    x"BF5D20AA",
    x"BF5D23D5",
    x"BF5D26FF",
    x"BF5D2A29",
    x"BF5D2D53",
    x"BF5D307D",
    x"BF5D33A7",
    x"BF5D36D0",
    x"BF5D39FA",
    x"BF5D3D23",
    x"BF5D404C",
    x"BF5D4376",
    x"BF5D469E",
    x"BF5D49C7",
    x"BF5D4CF0",
    x"BF5D5018",
    x"BF5D5341",
    x"BF5D5669",
    x"BF5D5991",
    x"BF5D5CB9",
    x"BF5D5FE1",
    x"BF5D6309",
    x"BF5D6631",
    x"BF5D6958",
    x"BF5D6C7F",
    x"BF5D6FA7",
    x"BF5D72CE",
    x"BF5D75F5",
    x"BF5D791B",
    x"BF5D7C42",
    x"BF5D7F69",
    x"BF5D828F",
    x"BF5D85B5",
    x"BF5D88DB",
    x"BF5D8C01",
    x"BF5D8F27",
    x"BF5D924D",
    x"BF5D9573",
    x"BF5D9898",
    x"BF5D9BBD",
    x"BF5D9EE3",
    x"BF5DA208",
    x"BF5DA52D",
    x"BF5DA851",
    x"BF5DAB76",
    x"BF5DAE9B",
    x"BF5DB1BF",
    x"BF5DB4E3",
    x"BF5DB807",
    x"BF5DBB2B",
    x"BF5DBE4F",
    x"BF5DC173",
    x"BF5DC497",
    x"BF5DC7BA",
    x"BF5DCADD",
    x"BF5DCE01",
    x"BF5DD124",
    x"BF5DD447",
    x"BF5DD769",
    x"BF5DDA8C",
    x"BF5DDDAF",
    x"BF5DE0D1",
    x"BF5DE3F3",
    x"BF5DE715",
    x"BF5DEA37",
    x"BF5DED59",
    x"BF5DF07B",
    x"BF5DF39D",
    x"BF5DF6BE",
    x"BF5DF9DF",
    x"BF5DFD01",
    x"BF5E0022",
    x"BF5E0343",
    x"BF5E0663",
    x"BF5E0984",
    x"BF5E0CA5",
    x"BF5E0FC5",
    x"BF5E12E5",
    x"BF5E1605",
    x"BF5E1925",
    x"BF5E1C45",
    x"BF5E1F65",
    x"BF5E2285",
    x"BF5E25A4",
    x"BF5E28C3",
    x"BF5E2BE3",
    x"BF5E2F02",
    x"BF5E3221",
    x"BF5E353F",
    x"BF5E385E",
    x"BF5E3B7D",
    x"BF5E3E9B",
    x"BF5E41B9",
    x"BF5E44D7",
    x"BF5E47F5",
    x"BF5E4B13",
    x"BF5E4E31",
    x"BF5E514E",
    x"BF5E546C",
    x"BF5E5789",
    x"BF5E5AA6",
    x"BF5E5DC3",
    x"BF5E60E0",
    x"BF5E63FD",
    x"BF5E671A",
    x"BF5E6A36",
    x"BF5E6D53",
    x"BF5E706F",
    x"BF5E738B",
    x"BF5E76A7",
    x"BF5E79C3",
    x"BF5E7CDE",
    x"BF5E7FFA",
    x"BF5E8316",
    x"BF5E8631",
    x"BF5E894C",
    x"BF5E8C67",
    x"BF5E8F82",
    x"BF5E929D",
    x"BF5E95B7",
    x"BF5E98D2",
    x"BF5E9BEC",
    x"BF5E9F06",
    x"BF5EA221",
    x"BF5EA53A",
    x"BF5EA854",
    x"BF5EAB6E",
    x"BF5EAE88",
    x"BF5EB1A1",
    x"BF5EB4BA",
    x"BF5EB7D3",
    x"BF5EBAEC",
    x"BF5EBE05",
    x"BF5EC11E",
    x"BF5EC437",
    x"BF5EC74F",
    x"BF5ECA68",
    x"BF5ECD80",
    x"BF5ED098",
    x"BF5ED3B0",
    x"BF5ED6C8",
    x"BF5ED9DF",
    x"BF5EDCF7",
    x"BF5EE00E",
    x"BF5EE326",
    x"BF5EE63D",
    x"BF5EE954",
    x"BF5EEC6B",
    x"BF5EEF81",
    x"BF5EF298",
    x"BF5EF5AE",
    x"BF5EF8C5",
    x"BF5EFBDB",
    x"BF5EFEF1",
    x"BF5F0207",
    x"BF5F051D",
    x"BF5F0833",
    x"BF5F0B48",
    x"BF5F0E5D",
    x"BF5F1173",
    x"BF5F1488",
    x"BF5F179D",
    x"BF5F1AB2",
    x"BF5F1DC6",
    x"BF5F20DB",
    x"BF5F23EF",
    x"BF5F2704",
    x"BF5F2A18",
    x"BF5F2D2C",
    x"BF5F3040",
    x"BF5F3354",
    x"BF5F3667",
    x"BF5F397B",
    x"BF5F3C8E",
    x"BF5F3FA2",
    x"BF5F42B5",
    x"BF5F45C8",
    x"BF5F48DB",
    x"BF5F4BED",
    x"BF5F4F00",
    x"BF5F5212",
    x"BF5F5525",
    x"BF5F5837",
    x"BF5F5B49",
    x"BF5F5E5B",
    x"BF5F616C",
    x"BF5F647E",
    x"BF5F6790",
    x"BF5F6AA1",
    x"BF5F6DB2",
    x"BF5F70C3",
    x"BF5F73D4",
    x"BF5F76E5",
    x"BF5F79F6",
    x"BF5F7D06",
    x"BF5F8017",
    x"BF5F8327",
    x"BF5F8637",
    x"BF5F8947",
    x"BF5F8C57",
    x"BF5F8F67",
    x"BF5F9276",
    x"BF5F9586",
    x"BF5F9895",
    x"BF5F9BA5",
    x"BF5F9EB4",
    x"BF5FA1C3",
    x"BF5FA4D1",
    x"BF5FA7E0",
    x"BF5FAAEF",
    x"BF5FADFD",
    x"BF5FB10B",
    x"BF5FB419",
    x"BF5FB727",
    x"BF5FBA35",
    x"BF5FBD43",
    x"BF5FC051",
    x"BF5FC35E",
    x"BF5FC66B",
    x"BF5FC979",
    x"BF5FCC86",
    x"BF5FCF93",
    x"BF5FD29F",
    x"BF5FD5AC",
    x"BF5FD8B8",
    x"BF5FDBC5",
    x"BF5FDED1",
    x"BF5FE1DD",
    x"BF5FE4E9",
    x"BF5FE7F5",
    x"BF5FEB01",
    x"BF5FEE0C",
    x"BF5FF118",
    x"BF5FF423",
    x"BF5FF72E",
    x"BF5FFA39",
    x"BF5FFD44",
    x"BF60004F",
    x"BF60035A",
    x"BF600664",
    x"BF60096E",
    x"BF600C79",
    x"BF600F83",
    x"BF60128D",
    x"BF601596",
    x"BF6018A0",
    x"BF601BAA",
    x"BF601EB3",
    x"BF6021BC",
    x"BF6024C6",
    x"BF6027CF",
    x"BF602AD7",
    x"BF602DE0",
    x"BF6030E9",
    x"BF6033F1",
    x"BF6036FA",
    x"BF603A02",
    x"BF603D0A",
    x"BF604012",
    x"BF60431A",
    x"BF604621",
    x"BF604929",
    x"BF604C30",
    x"BF604F37",
    x"BF60523E",
    x"BF605545",
    x"BF60584C",
    x"BF605B53",
    x"BF605E5A",
    x"BF606160",
    x"BF606466",
    x"BF60676D",
    x"BF606A73",
    x"BF606D78",
    x"BF60707E",
    x"BF607384",
    x"BF607689",
    x"BF60798F",
    x"BF607C94",
    x"BF607F99",
    x"BF60829E",
    x"BF6085A3",
    x"BF6088A7",
    x"BF608BAC",
    x"BF608EB0",
    x"BF6091B5",
    x"BF6094B9",
    x"BF6097BD",
    x"BF609AC1",
    x"BF609DC4",
    x"BF60A0C8",
    x"BF60A3CC",
    x"BF60A6CF",
    x"BF60A9D2",
    x"BF60ACD5",
    x"BF60AFD8",
    x"BF60B2DB",
    x"BF60B5DE",
    x"BF60B8E0",
    x"BF60BBE2",
    x"BF60BEE5",
    x"BF60C1E7",
    x"BF60C4E9",
    x"BF60C7EB",
    x"BF60CAEC",
    x"BF60CDEE",
    x"BF60D0EF",
    x"BF60D3F1",
    x"BF60D6F2",
    x"BF60D9F3",
    x"BF60DCF4",
    x"BF60DFF4",
    x"BF60E2F5",
    x"BF60E5F6",
    x"BF60E8F6",
    x"BF60EBF6",
    x"BF60EEF6",
    x"BF60F1F6",
    x"BF60F4F6",
    x"BF60F7F6",
    x"BF60FAF5",
    x"BF60FDF5",
    x"BF6100F4",
    x"BF6103F3",
    x"BF6106F2",
    x"BF6109F1",
    x"BF610CF0",
    x"BF610FEE",
    x"BF6112ED",
    x"BF6115EB",
    x"BF6118E9",
    x"BF611BE7",
    x"BF611EE5",
    x"BF6121E3",
    x"BF6124E1",
    x"BF6127DE",
    x"BF612ADB",
    x"BF612DD9",
    x"BF6130D6",
    x"BF6133D3",
    x"BF6136D0",
    x"BF6139CC",
    x"BF613CC9",
    x"BF613FC5",
    x"BF6142C1",
    x"BF6145BE",
    x"BF6148BA",
    x"BF614BB5",
    x"BF614EB1",
    x"BF6151AD",
    x"BF6154A8",
    x"BF6157A4",
    x"BF615A9F",
    x"BF615D9A",
    x"BF616095",
    x"BF616390",
    x"BF61668A",
    x"BF616985",
    x"BF616C7F",
    x"BF616F79",
    x"BF617274",
    x"BF61756E",
    x"BF617867",
    x"BF617B61",
    x"BF617E5B",
    x"BF618154",
    x"BF61844D",
    x"BF618747",
    x"BF618A40",
    x"BF618D38",
    x"BF619031",
    x"BF61932A",
    x"BF619622",
    x"BF61991B",
    x"BF619C13",
    x"BF619F0B",
    x"BF61A203",
    x"BF61A4FB",
    x"BF61A7F2",
    x"BF61AAEA",
    x"BF61ADE1",
    x"BF61B0D9",
    x"BF61B3D0",
    x"BF61B6C7",
    x"BF61B9BE",
    x"BF61BCB4",
    x"BF61BFAB",
    x"BF61C2A1",
    x"BF61C598",
    x"BF61C88E",
    x"BF61CB84",
    x"BF61CE7A",
    x"BF61D16F",
    x"BF61D465",
    x"BF61D75B",
    x"BF61DA50",
    x"BF61DD45",
    x"BF61E03A",
    x"BF61E32F",
    x"BF61E624",
    x"BF61E919",
    x"BF61EC0D",
    x"BF61EF02",
    x"BF61F1F6",
    x"BF61F4EA",
    x"BF61F7DE",
    x"BF61FAD2",
    x"BF61FDC6",
    x"BF6200B9",
    x"BF6203AD",
    x"BF6206A0",
    x"BF620993",
    x"BF620C86",
    x"BF620F79",
    x"BF62126C",
    x"BF62155E",
    x"BF621851",
    x"BF621B43",
    x"BF621E35",
    x"BF622128",
    x"BF62241A",
    x"BF62270B",
    x"BF6229FD",
    x"BF622CEF",
    x"BF622FE0",
    x"BF6232D1",
    x"BF6235C2",
    x"BF6238B3",
    x"BF623BA4",
    x"BF623E95",
    x"BF624186",
    x"BF624476",
    x"BF624766",
    x"BF624A57",
    x"BF624D47",
    x"BF625036",
    x"BF625326",
    x"BF625616",
    x"BF625905",
    x"BF625BF5",
    x"BF625EE4",
    x"BF6261D3",
    x"BF6264C2",
    x"BF6267B1",
    x"BF626AA0",
    x"BF626D8E",
    x"BF62707C",
    x"BF62736B",
    x"BF627659",
    x"BF627947",
    x"BF627C35",
    x"BF627F22",
    x"BF628210",
    x"BF6284FD",
    x"BF6287EB",
    x"BF628AD8",
    x"BF628DC5",
    x"BF6290B2",
    x"BF62939F",
    x"BF62968B",
    x"BF629978",
    x"BF629C64",
    x"BF629F50",
    x"BF62A23D",
    x"BF62A528",
    x"BF62A814",
    x"BF62AB00",
    x"BF62ADEB",
    x"BF62B0D7",
    x"BF62B3C2",
    x"BF62B6AD",
    x"BF62B998",
    x"BF62BC83",
    x"BF62BF6E",
    x"BF62C258",
    x"BF62C543",
    x"BF62C82D",
    x"BF62CB17",
    x"BF62CE01",
    x"BF62D0EB",
    x"BF62D3D5",
    x"BF62D6BF",
    x"BF62D9A8",
    x"BF62DC92",
    x"BF62DF7B",
    x"BF62E264",
    x"BF62E54D",
    x"BF62E836",
    x"BF62EB1E",
    x"BF62EE07",
    x"BF62F0EF",
    x"BF62F3D8",
    x"BF62F6C0",
    x"BF62F9A8",
    x"BF62FC8F",
    x"BF62FF77",
    x"BF63025F",
    x"BF630546",
    x"BF63082E",
    x"BF630B15",
    x"BF630DFC",
    x"BF6310E3",
    x"BF6313C9",
    x"BF6316B0",
    x"BF631996",
    x"BF631C7D",
    x"BF631F63",
    x"BF632249",
    x"BF63252F",
    x"BF632815",
    x"BF632AFB",
    x"BF632DE0",
    x"BF6330C5",
    x"BF6333AB",
    x"BF633690",
    x"BF633975",
    x"BF633C5A",
    x"BF633F3E",
    x"BF634223",
    x"BF634507",
    x"BF6347EC",
    x"BF634AD0",
    x"BF634DB4",
    x"BF635098",
    x"BF63537B",
    x"BF63565F",
    x"BF635943",
    x"BF635C26",
    x"BF635F09",
    x"BF6361EC",
    x"BF6364CF",
    x"BF6367B2",
    x"BF636A95",
    x"BF636D77",
    x"BF637059",
    x"BF63733C",
    x"BF63761E",
    x"BF637900",
    x"BF637BE2",
    x"BF637EC3",
    x"BF6381A5",
    x"BF638486",
    x"BF638767",
    x"BF638A49",
    x"BF638D2A",
    x"BF63900B",
    x"BF6392EB",
    x"BF6395CC",
    x"BF6398AC",
    x"BF639B8D",
    x"BF639E6D",
    x"BF63A14D",
    x"BF63A42D",
    x"BF63A70D",
    x"BF63A9EC",
    x"BF63ACCC",
    x"BF63AFAB",
    x"BF63B28A",
    x"BF63B569",
    x"BF63B848",
    x"BF63BB27",
    x"BF63BE06",
    x"BF63C0E4",
    x"BF63C3C3",
    x"BF63C6A1",
    x"BF63C97F",
    x"BF63CC5D",
    x"BF63CF3B",
    x"BF63D219",
    x"BF63D4F6",
    x"BF63D7D4",
    x"BF63DAB1",
    x"BF63DD8E",
    x"BF63E06B",
    x"BF63E348",
    x"BF63E625",
    x"BF63E901",
    x"BF63EBDE",
    x"BF63EEBA",
    x"BF63F196",
    x"BF63F473",
    x"BF63F74E",
    x"BF63FA2A",
    x"BF63FD06",
    x"BF63FFE1",
    x"BF6402BD",
    x"BF640598",
    x"BF640873",
    x"BF640B4E",
    x"BF640E29",
    x"BF641104",
    x"BF6413DE",
    x"BF6416B9",
    x"BF641993",
    x"BF641C6D",
    x"BF641F47",
    x"BF642221",
    x"BF6424FB",
    x"BF6427D4",
    x"BF642AAE",
    x"BF642D87",
    x"BF643060",
    x"BF643339",
    x"BF643612",
    x"BF6438EB",
    x"BF643BC4",
    x"BF643E9C",
    x"BF644174",
    x"BF64444D",
    x"BF644725",
    x"BF6449FD",
    x"BF644CD5",
    x"BF644FAC",
    x"BF645284",
    x"BF64555B",
    x"BF645832",
    x"BF645B0A",
    x"BF645DE1",
    x"BF6460B7",
    x"BF64638E",
    x"BF646665",
    x"BF64693B",
    x"BF646C11",
    x"BF646EE8",
    x"BF6471BE",
    x"BF647493",
    x"BF647769",
    x"BF647A3F",
    x"BF647D14",
    x"BF647FEA",
    x"BF6482BF",
    x"BF648594",
    x"BF648869",
    x"BF648B3E",
    x"BF648E12",
    x"BF6490E7",
    x"BF6493BB",
    x"BF64968F",
    x"BF649963",
    x"BF649C37",
    x"BF649F0B",
    x"BF64A1DF",
    x"BF64A4B2",
    x"BF64A786",
    x"BF64AA59",
    x"BF64AD2C",
    x"BF64AFFF",
    x"BF64B2D2",
    x"BF64B5A5",
    x"BF64B877",
    x"BF64BB4A",
    x"BF64BE1C",
    x"BF64C0EE",
    x"BF64C3C0",
    x"BF64C692",
    x"BF64C964",
    x"BF64CC35",
    x"BF64CF07",
    x"BF64D1D8",
    x"BF64D4AA",
    x"BF64D77B",
    x"BF64DA4B",
    x"BF64DD1C",
    x"BF64DFED",
    x"BF64E2BD",
    x"BF64E58E",
    x"BF64E85E",
    x"BF64EB2E",
    x"BF64EDFE",
    x"BF64F0CE",
    x"BF64F39E",
    x"BF64F66D",
    x"BF64F93D",
    x"BF64FC0C",
    x"BF64FEDB",
    x"BF6501AA",
    x"BF650479",
    x"BF650748",
    x"BF650A16",
    x"BF650CE5",
    x"BF650FB3",
    x"BF651281",
    x"BF65154F",
    x"BF65181D",
    x"BF651AEB",
    x"BF651DB8",
    x"BF652086",
    x"BF652353",
    x"BF652620",
    x"BF6528ED",
    x"BF652BBA",
    x"BF652E87",
    x"BF653154",
    x"BF653420",
    x"BF6536ED",
    x"BF6539B9",
    x"BF653C85",
    x"BF653F51",
    x"BF65421D",
    x"BF6544E8",
    x"BF6547B4",
    x"BF654A7F",
    x"BF654D4B",
    x"BF655016",
    x"BF6552E1",
    x"BF6555AC",
    x"BF655876",
    x"BF655B41",
    x"BF655E0B",
    x"BF6560D6",
    x"BF6563A0",
    x"BF65666A",
    x"BF656934",
    x"BF656BFD",
    x"BF656EC7",
    x"BF657190",
    x"BF65745A",
    x"BF657723",
    x"BF6579EC",
    x"BF657CB5",
    x"BF657F7E",
    x"BF658246",
    x"BF65850F",
    x"BF6587D7",
    x"BF658AA0",
    x"BF658D68",
    x"BF659030",
    x"BF6592F7",
    x"BF6595BF",
    x"BF659887",
    x"BF659B4E",
    x"BF659E15",
    x"BF65A0DC",
    x"BF65A3A3",
    x"BF65A66A",
    x"BF65A931",
    x"BF65ABF7",
    x"BF65AEBE",
    x"BF65B184",
    x"BF65B44A",
    x"BF65B710",
    x"BF65B9D6",
    x"BF65BC9C",
    x"BF65BF62",
    x"BF65C227",
    x"BF65C4EC",
    x"BF65C7B1",
    x"BF65CA77",
    x"BF65CD3B",
    x"BF65D000",
    x"BF65D2C5",
    x"BF65D589",
    x"BF65D84E",
    x"BF65DB12",
    x"BF65DDD6",
    x"BF65E09A",
    x"BF65E35E",
    x"BF65E621",
    x"BF65E8E5",
    x"BF65EBA8",
    x"BF65EE6C",
    x"BF65F12F",
    x"BF65F3F2",
    x"BF65F6B4",
    x"BF65F977",
    x"BF65FC3A",
    x"BF65FEFC",
    x"BF6601BE",
    x"BF660480",
    x"BF660742",
    x"BF660A04",
    x"BF660CC6",
    x"BF660F88",
    x"BF661249",
    x"BF66150A",
    x"BF6617CC",
    x"BF661A8D",
    x"BF661D4D",
    x"BF66200E",
    x"BF6622CF",
    x"BF66258F",
    x"BF662850",
    x"BF662B10",
    x"BF662DD0",
    x"BF663090",
    x"BF663350",
    x"BF66360F",
    x"BF6638CF",
    x"BF663B8E",
    x"BF663E4D",
    x"BF66410C",
    x"BF6643CB",
    x"BF66468A",
    x"BF664949",
    x"BF664C07",
    x"BF664EC6",
    x"BF665184",
    x"BF665442",
    x"BF665700",
    x"BF6659BE",
    x"BF665C7C",
    x"BF665F39",
    x"BF6661F7",
    x"BF6664B4",
    x"BF666771",
    x"BF666A2E",
    x"BF666CEB",
    x"BF666FA8",
    x"BF667264",
    x"BF667521",
    x"BF6677DD",
    x"BF667A99",
    x"BF667D55",
    x"BF668011",
    x"BF6682CD",
    x"BF668588",
    x"BF668844",
    x"BF668AFF",
    x"BF668DBA",
    x"BF669076",
    x"BF669330",
    x"BF6695EB",
    x"BF6698A6",
    x"BF669B60",
    x"BF669E1B",
    x"BF66A0D5",
    x"BF66A38F",
    x"BF66A649",
    x"BF66A903",
    x"BF66ABBC",
    x"BF66AE76",
    x"BF66B12F",
    x"BF66B3E9",
    x"BF66B6A2",
    x"BF66B95B",
    x"BF66BC14",
    x"BF66BECC",
    x"BF66C185",
    x"BF66C43D",
    x"BF66C6F6",
    x"BF66C9AE",
    x"BF66CC66",
    x"BF66CF1E",
    x"BF66D1D5",
    x"BF66D48D",
    x"BF66D744",
    x"BF66D9FC",
    x"BF66DCB3",
    x"BF66DF6A",
    x"BF66E221",
    x"BF66E4D7",
    x"BF66E78E",
    x"BF66EA45",
    x"BF66ECFB",
    x"BF66EFB1",
    x"BF66F267",
    x"BF66F51D",
    x"BF66F7D3",
    x"BF66FA88",
    x"BF66FD3E",
    x"BF66FFF3",
    x"BF6702A9",
    x"BF67055E",
    x"BF670813",
    x"BF670AC7",
    x"BF670D7C",
    x"BF671031",
    x"BF6712E5",
    x"BF671599",
    x"BF67184D",
    x"BF671B01",
    x"BF671DB5",
    x"BF672069",
    x"BF67231C",
    x"BF6725D0",
    x"BF672883",
    x"BF672B36",
    x"BF672DE9",
    x"BF67309C",
    x"BF67334F",
    x"BF673601",
    x"BF6738B4",
    x"BF673B66",
    x"BF673E18",
    x"BF6740CA",
    x"BF67437C",
    x"BF67462E",
    x"BF6748DF",
    x"BF674B91",
    x"BF674E42",
    x"BF6750F3",
    x"BF6753A5",
    x"BF675655",
    x"BF675906",
    x"BF675BB7",
    x"BF675E67",
    x"BF676118",
    x"BF6763C8",
    x"BF676678",
    x"BF676928",
    x"BF676BD8",
    x"BF676E87",
    x"BF677137",
    x"BF6773E6",
    x"BF677695",
    x"BF677944",
    x"BF677BF3",
    x"BF677EA2",
    x"BF678151",
    x"BF6783FF",
    x"BF6786AE",
    x"BF67895C",
    x"BF678C0A",
    x"BF678EB8",
    x"BF679166",
    x"BF679414",
    x"BF6796C1",
    x"BF67996F",
    x"BF679C1C",
    x"BF679EC9",
    x"BF67A176",
    x"BF67A423",
    x"BF67A6D0",
    x"BF67A97C",
    x"BF67AC29",
    x"BF67AED5",
    x"BF67B181",
    x"BF67B42D",
    x"BF67B6D9",
    x"BF67B985",
    x"BF67BC30",
    x"BF67BEDC",
    x"BF67C187",
    x"BF67C432",
    x"BF67C6DE",
    x"BF67C988",
    x"BF67CC33",
    x"BF67CEDE",
    x"BF67D188",
    x"BF67D433",
    x"BF67D6DD",
    x"BF67D987",
    x"BF67DC31",
    x"BF67DEDB",
    x"BF67E184",
    x"BF67E42E",
    x"BF67E6D7",
    x"BF67E980",
    x"BF67EC29",
    x"BF67EED2",
    x"BF67F17B",
    x"BF67F424",
    x"BF67F6CC",
    x"BF67F975",
    x"BF67FC1D",
    x"BF67FEC5",
    x"BF68016D",
    x"BF680415",
    x"BF6806BD",
    x"BF680964",
    x"BF680C0C",
    x"BF680EB3",
    x"BF68115A",
    x"BF681401",
    x"BF6816A8",
    x"BF68194F",
    x"BF681BF5",
    x"BF681E9C",
    x"BF682142",
    x"BF6823E8",
    x"BF68268E",
    x"BF682934",
    x"BF682BDA",
    x"BF682E7F",
    x"BF683125",
    x"BF6833CA",
    x"BF68366F",
    x"BF683914",
    x"BF683BB9",
    x"BF683E5E",
    x"BF684103",
    x"BF6843A7",
    x"BF68464B",
    x"BF6848F0",
    x"BF684B94",
    x"BF684E38",
    x"BF6850DB",
    x"BF68537F",
    x"BF685623",
    x"BF6858C6",
    x"BF685B69",
    x"BF685E0C",
    x"BF6860AF",
    x"BF686352",
    x"BF6865F5",
    x"BF686897",
    x"BF686B39",
    x"BF686DDC",
    x"BF68707E",
    x"BF687320",
    x"BF6875C2",
    x"BF687863",
    x"BF687B05",
    x"BF687DA6",
    x"BF688047",
    x"BF6882E9",
    x"BF68858A",
    x"BF68882A",
    x"BF688ACB",
    x"BF688D6C",
    x"BF68900C",
    x"BF6892AC",
    x"BF68954C",
    x"BF6897EC",
    x"BF689A8C",
    x"BF689D2C",
    x"BF689FCC",
    x"BF68A26B",
    x"BF68A50A",
    x"BF68A7AA",
    x"BF68AA49",
    x"BF68ACE7",
    x"BF68AF86",
    x"BF68B225",
    x"BF68B4C3",
    x"BF68B762",
    x"BF68BA00",
    x"BF68BC9E",
    x"BF68BF3C",
    x"BF68C1D9",
    x"BF68C477",
    x"BF68C714",
    x"BF68C9B2",
    x"BF68CC4F",
    x"BF68CEEC",
    x"BF68D189",
    x"BF68D426",
    x"BF68D6C2",
    x"BF68D95F",
    x"BF68DBFB",
    x"BF68DE97",
    x"BF68E134",
    x"BF68E3CF",
    x"BF68E66B",
    x"BF68E907",
    x"BF68EBA2",
    x"BF68EE3E",
    x"BF68F0D9",
    x"BF68F374",
    x"BF68F60F",
    x"BF68F8AA",
    x"BF68FB45",
    x"BF68FDDF",
    x"BF690079",
    x"BF690314",
    x"BF6905AE",
    x"BF690848",
    x"BF690AE2",
    x"BF690D7B",
    x"BF691015",
    x"BF6912AE",
    x"BF691547",
    x"BF6917E1",
    x"BF691A7A",
    x"BF691D12",
    x"BF691FAB",
    x"BF692244",
    x"BF6924DC",
    x"BF692774",
    x"BF692A0D",
    x"BF692CA5",
    x"BF692F3C",
    x"BF6931D4",
    x"BF69346C",
    x"BF693703",
    x"BF69399A",
    x"BF693C32",
    x"BF693EC9",
    x"BF694160",
    x"BF6943F6",
    x"BF69468D",
    x"BF694923",
    x"BF694BBA",
    x"BF694E50",
    x"BF6950E6",
    x"BF69537C",
    x"BF695611",
    x"BF6958A7",
    x"BF695B3D",
    x"BF695DD2",
    x"BF696067",
    x"BF6962FC",
    x"BF696591",
    x"BF696826",
    x"BF696ABA",
    x"BF696D4F",
    x"BF696FE3",
    x"BF697277",
    x"BF69750C",
    x"BF69779F",
    x"BF697A33",
    x"BF697CC7",
    x"BF697F5A",
    x"BF6981EE",
    x"BF698481",
    x"BF698714",
    x"BF6989A7",
    x"BF698C3A",
    x"BF698ECC",
    x"BF69915F",
    x"BF6993F1",
    x"BF699684",
    x"BF699916",
    x"BF699BA8",
    x"BF699E39",
    x"BF69A0CB",
    x"BF69A35D",
    x"BF69A5EE",
    x"BF69A87F",
    x"BF69AB10",
    x"BF69ADA1",
    x"BF69B032",
    x"BF69B2C3",
    x"BF69B553",
    x"BF69B7E4",
    x"BF69BA74",
    x"BF69BD04",
    x"BF69BF94",
    x"BF69C224",
    x"BF69C4B4",
    x"BF69C743",
    x"BF69C9D3",
    x"BF69CC62",
    x"BF69CEF1",
    x"BF69D180",
    x"BF69D40F",
    x"BF69D69E",
    x"BF69D92C",
    x"BF69DBBB",
    x"BF69DE49",
    x"BF69E0D7",
    x"BF69E365",
    x"BF69E5F3",
    x"BF69E881",
    x"BF69EB0E",
    x"BF69ED9C",
    x"BF69F029",
    x"BF69F2B6",
    x"BF69F543",
    x"BF69F7D0",
    x"BF69FA5D",
    x"BF69FCEA",
    x"BF69FF76",
    x"BF6A0202",
    x"BF6A048F",
    x"BF6A071B",
    x"BF6A09A7",
    x"BF6A0C32",
    x"BF6A0EBE",
    x"BF6A1149",
    x"BF6A13D5",
    x"BF6A1660",
    x"BF6A18EB",
    x"BF6A1B76",
    x"BF6A1E01",
    x"BF6A208B",
    x"BF6A2316",
    x"BF6A25A0",
    x"BF6A282A",
    x"BF6A2AB4",
    x"BF6A2D3E",
    x"BF6A2FC8",
    x"BF6A3252",
    x"BF6A34DB",
    x"BF6A3765",
    x"BF6A39EE",
    x"BF6A3C77",
    x"BF6A3F00",
    x"BF6A4189",
    x"BF6A4411",
    x"BF6A469A",
    x"BF6A4922",
    x"BF6A4BAA",
    x"BF6A4E33",
    x"BF6A50BA",
    x"BF6A5342",
    x"BF6A55CA",
    x"BF6A5851",
    x"BF6A5AD9",
    x"BF6A5D60",
    x"BF6A5FE7",
    x"BF6A626E",
    x"BF6A64F5",
    x"BF6A677C",
    x"BF6A6A02",
    x"BF6A6C89",
    x"BF6A6F0F",
    x"BF6A7195",
    x"BF6A741B",
    x"BF6A76A1",
    x"BF6A7926",
    x"BF6A7BAC",
    x"BF6A7E31",
    x"BF6A80B7",
    x"BF6A833C",
    x"BF6A85C1",
    x"BF6A8846",
    x"BF6A8ACA",
    x"BF6A8D4F",
    x"BF6A8FD3",
    x"BF6A9258",
    x"BF6A94DC",
    x"BF6A9760",
    x"BF6A99E4",
    x"BF6A9C67",
    x"BF6A9EEB",
    x"BF6AA16E",
    x"BF6AA3F2",
    x"BF6AA675",
    x"BF6AA8F8",
    x"BF6AAB7B",
    x"BF6AADFD",
    x"BF6AB080",
    x"BF6AB302",
    x"BF6AB585",
    x"BF6AB807",
    x"BF6ABA89",
    x"BF6ABD0B",
    x"BF6ABF8C",
    x"BF6AC20E",
    x"BF6AC48F",
    x"BF6AC711",
    x"BF6AC992",
    x"BF6ACC13",
    x"BF6ACE94",
    x"BF6AD115",
    x"BF6AD395",
    x"BF6AD616",
    x"BF6AD896",
    x"BF6ADB16",
    x"BF6ADD96",
    x"BF6AE016",
    x"BF6AE296",
    x"BF6AE515",
    x"BF6AE795",
    x"BF6AEA14",
    x"BF6AEC93",
    x"BF6AEF12",
    x"BF6AF191",
    x"BF6AF410",
    x"BF6AF68F",
    x"BF6AF90D",
    x"BF6AFB8C",
    x"BF6AFE0A",
    x"BF6B0088",
    x"BF6B0306",
    x"BF6B0584",
    x"BF6B0801",
    x"BF6B0A7F",
    x"BF6B0CFC",
    x"BF6B0F79",
    x"BF6B11F6",
    x"BF6B1473",
    x"BF6B16F0",
    x"BF6B196D",
    x"BF6B1BE9",
    x"BF6B1E65",
    x"BF6B20E2",
    x"BF6B235E",
    x"BF6B25DA",
    x"BF6B2855",
    x"BF6B2AD1",
    x"BF6B2D4D",
    x"BF6B2FC8",
    x"BF6B3243",
    x"BF6B34BE",
    x"BF6B3739",
    x"BF6B39B4",
    x"BF6B3C2F",
    x"BF6B3EA9",
    x"BF6B4124",
    x"BF6B439E",
    x"BF6B4618",
    x"BF6B4892",
    x"BF6B4B0C",
    x"BF6B4D85",
    x"BF6B4FFF",
    x"BF6B5278",
    x"BF6B54F1",
    x"BF6B576B",
    x"BF6B59E3",
    x"BF6B5C5C",
    x"BF6B5ED5",
    x"BF6B614D",
    x"BF6B63C6",
    x"BF6B663E",
    x"BF6B68B6",
    x"BF6B6B2E",
    x"BF6B6DA6",
    x"BF6B701E",
    x"BF6B7295",
    x"BF6B750D",
    x"BF6B7784",
    x"BF6B79FB",
    x"BF6B7C72",
    x"BF6B7EE9",
    x"BF6B815F",
    x"BF6B83D6",
    x"BF6B864C",
    x"BF6B88C3",
    x"BF6B8B39",
    x"BF6B8DAF",
    x"BF6B9025",
    x"BF6B929A",
    x"BF6B9510",
    x"BF6B9785",
    x"BF6B99FB",
    x"BF6B9C70",
    x"BF6B9EE5",
    x"BF6BA159",
    x"BF6BA3CE",
    x"BF6BA643",
    x"BF6BA8B7",
    x"BF6BAB2B",
    x"BF6BADA0",
    x"BF6BB014",
    x"BF6BB287",
    x"BF6BB4FB",
    x"BF6BB76F",
    x"BF6BB9E2",
    x"BF6BBC55",
    x"BF6BBEC8",
    x"BF6BC13B",
    x"BF6BC3AE",
    x"BF6BC621",
    x"BF6BC894",
    x"BF6BCB06",
    x"BF6BCD78",
    x"BF6BCFEA",
    x"BF6BD25C",
    x"BF6BD4CE",
    x"BF6BD740",
    x"BF6BD9B2",
    x"BF6BDC23",
    x"BF6BDE94",
    x"BF6BE105",
    x"BF6BE376",
    x"BF6BE5E7",
    x"BF6BE858",
    x"BF6BEAC9",
    x"BF6BED39",
    x"BF6BEFA9",
    x"BF6BF21A",
    x"BF6BF48A",
    x"BF6BF6F9",
    x"BF6BF969",
    x"BF6BFBD9",
    x"BF6BFE48",
    x"BF6C00B7",
    x"BF6C0327",
    x"BF6C0596",
    x"BF6C0805",
    x"BF6C0A73",
    x"BF6C0CE2",
    x"BF6C0F50",
    x"BF6C11BF",
    x"BF6C142D",
    x"BF6C169B",
    x"BF6C1909",
    x"BF6C1B76",
    x"BF6C1DE4",
    x"BF6C2051",
    x"BF6C22BF",
    x"BF6C252C",
    x"BF6C2799",
    x"BF6C2A06",
    x"BF6C2C73",
    x"BF6C2EDF",
    x"BF6C314C",
    x"BF6C33B8",
    x"BF6C3624",
    x"BF6C3890",
    x"BF6C3AFC",
    x"BF6C3D68",
    x"BF6C3FD3",
    x"BF6C423F",
    x"BF6C44AA",
    x"BF6C4715",
    x"BF6C4980",
    x"BF6C4BEB",
    x"BF6C4E56",
    x"BF6C50C1",
    x"BF6C532B",
    x"BF6C5595",
    x"BF6C5800",
    x"BF6C5A6A",
    x"BF6C5CD4",
    x"BF6C5F3D",
    x"BF6C61A7",
    x"BF6C6410",
    x"BF6C667A",
    x"BF6C68E3",
    x"BF6C6B4C",
    x"BF6C6DB5",
    x"BF6C701E",
    x"BF6C7286",
    x"BF6C74EF",
    x"BF6C7757",
    x"BF6C79BF",
    x"BF6C7C27",
    x"BF6C7E8F",
    x"BF6C80F7",
    x"BF6C835E",
    x"BF6C85C6",
    x"BF6C882D",
    x"BF6C8A94",
    x"BF6C8CFC",
    x"BF6C8F62",
    x"BF6C91C9",
    x"BF6C9430",
    x"BF6C9696",
    x"BF6C98FD",
    x"BF6C9B63",
    x"BF6C9DC9",
    x"BF6CA02F",
    x"BF6CA295",
    x"BF6CA4FA",
    x"BF6CA760",
    x"BF6CA9C5",
    x"BF6CAC2A",
    x"BF6CAE8F",
    x"BF6CB0F4",
    x"BF6CB359",
    x"BF6CB5BD",
    x"BF6CB822",
    x"BF6CBA86",
    x"BF6CBCEA",
    x"BF6CBF4F",
    x"BF6CC1B2",
    x"BF6CC416",
    x"BF6CC67A",
    x"BF6CC8DD",
    x"BF6CCB41",
    x"BF6CCDA4",
    x"BF6CD007",
    x"BF6CD26A",
    x"BF6CD4CD",
    x"BF6CD72F",
    x"BF6CD992",
    x"BF6CDBF4",
    x"BF6CDE56",
    x"BF6CE0B8",
    x"BF6CE31A",
    x"BF6CE57C",
    x"BF6CE7DE",
    x"BF6CEA3F",
    x"BF6CECA0",
    x"BF6CEF02",
    x"BF6CF163",
    x"BF6CF3C4",
    x"BF6CF624",
    x"BF6CF885",
    x"BF6CFAE5",
    x"BF6CFD46",
    x"BF6CFFA6",
    x"BF6D0206",
    x"BF6D0466",
    x"BF6D06C6",
    x"BF6D0925",
    x"BF6D0B85",
    x"BF6D0DE4",
    x"BF6D1043",
    x"BF6D12A2",
    x"BF6D1501",
    x"BF6D1760",
    x"BF6D19BF",
    x"BF6D1C1D",
    x"BF6D1E7C",
    x"BF6D20DA",
    x"BF6D2338",
    x"BF6D2596",
    x"BF6D27F4",
    x"BF6D2A51",
    x"BF6D2CAF",
    x"BF6D2F0C",
    x"BF6D3169",
    x"BF6D33C6",
    x"BF6D3623",
    x"BF6D3880",
    x"BF6D3ADD",
    x"BF6D3D39",
    x"BF6D3F95",
    x"BF6D41F2",
    x"BF6D444E",
    x"BF6D46AA",
    x"BF6D4905",
    x"BF6D4B61",
    x"BF6D4DBC",
    x"BF6D5018",
    x"BF6D5273",
    x"BF6D54CE",
    x"BF6D5729",
    x"BF6D5984",
    x"BF6D5BDE",
    x"BF6D5E39",
    x"BF6D6093",
    x"BF6D62ED",
    x"BF6D6547",
    x"BF6D67A1",
    x"BF6D69FB",
    x"BF6D6C55",
    x"BF6D6EAE",
    x"BF6D7108",
    x"BF6D7361",
    x"BF6D75BA",
    x"BF6D7813",
    x"BF6D7A6C",
    x"BF6D7CC4",
    x"BF6D7F1D",
    x"BF6D8175",
    x"BF6D83CD",
    x"BF6D8625",
    x"BF6D887D",
    x"BF6D8AD5",
    x"BF6D8D2D",
    x"BF6D8F84",
    x"BF6D91DB",
    x"BF6D9433",
    x"BF6D968A",
    x"BF6D98E1",
    x"BF6D9B37",
    x"BF6D9D8E",
    x"BF6D9FE4",
    x"BF6DA23B",
    x"BF6DA491",
    x"BF6DA6E7",
    x"BF6DA93D",
    x"BF6DAB93",
    x"BF6DADE8",
    x"BF6DB03E",
    x"BF6DB293",
    x"BF6DB4E8",
    x"BF6DB73D",
    x"BF6DB992",
    x"BF6DBBE7",
    x"BF6DBE3C",
    x"BF6DC090",
    x"BF6DC2E4",
    x"BF6DC539",
    x"BF6DC78D",
    x"BF6DC9E1",
    x"BF6DCC34",
    x"BF6DCE88",
    x"BF6DD0DB",
    x"BF6DD32F",
    x"BF6DD582",
    x"BF6DD7D5",
    x"BF6DDA28",
    x"BF6DDC7B",
    x"BF6DDECD",
    x"BF6DE120",
    x"BF6DE372",
    x"BF6DE5C4",
    x"BF6DE816",
    x"BF6DEA68",
    x"BF6DECBA",
    x"BF6DEF0B",
    x"BF6DF15D",
    x"BF6DF3AE",
    x"BF6DF5FF",
    x"BF6DF850",
    x"BF6DFAA1",
    x"BF6DFCF2",
    x"BF6DFF43",
    x"BF6E0193",
    x"BF6E03E3",
    x"BF6E0634",
    x"BF6E0884",
    x"BF6E0AD4",
    x"BF6E0D23",
    x"BF6E0F73",
    x"BF6E11C2",
    x"BF6E1412",
    x"BF6E1661",
    x"BF6E18B0",
    x"BF6E1AFF",
    x"BF6E1D4E",
    x"BF6E1F9C",
    x"BF6E21EB",
    x"BF6E2439",
    x"BF6E2687",
    x"BF6E28D5",
    x"BF6E2B23",
    x"BF6E2D71",
    x"BF6E2FBE",
    x"BF6E320C",
    x"BF6E3459",
    x"BF6E36A6",
    x"BF6E38F3",
    x"BF6E3B40",
    x"BF6E3D8D",
    x"BF6E3FD9",
    x"BF6E4226",
    x"BF6E4472",
    x"BF6E46BE",
    x"BF6E490A",
    x"BF6E4B56",
    x"BF6E4DA2",
    x"BF6E4FEE",
    x"BF6E5239",
    x"BF6E5484",
    x"BF6E56CF",
    x"BF6E591A",
    x"BF6E5B65",
    x"BF6E5DB0",
    x"BF6E5FFB",
    x"BF6E6245",
    x"BF6E648F",
    x"BF6E66D9",
    x"BF6E6924",
    x"BF6E6B6D",
    x"BF6E6DB7",
    x"BF6E7001",
    x"BF6E724A",
    x"BF6E7493",
    x"BF6E76DD",
    x"BF6E7926",
    x"BF6E7B6E",
    x"BF6E7DB7",
    x"BF6E8000",
    x"BF6E8248",
    x"BF6E8490",
    x"BF6E86D8",
    x"BF6E8920",
    x"BF6E8B68",
    x"BF6E8DB0",
    x"BF6E8FF8",
    x"BF6E923F",
    x"BF6E9486",
    x"BF6E96CD",
    x"BF6E9914",
    x"BF6E9B5B",
    x"BF6E9DA2",
    x"BF6E9FE9",
    x"BF6EA22F",
    x"BF6EA475",
    x"BF6EA6BB",
    x"BF6EA901",
    x"BF6EAB47",
    x"BF6EAD8D",
    x"BF6EAFD2",
    x"BF6EB218",
    x"BF6EB45D",
    x"BF6EB6A2",
    x"BF6EB8E7",
    x"BF6EBB2C",
    x"BF6EBD71",
    x"BF6EBFB5",
    x"BF6EC1FA",
    x"BF6EC43E",
    x"BF6EC682",
    x"BF6EC8C6",
    x"BF6ECB0A",
    x"BF6ECD4D",
    x"BF6ECF91",
    x"BF6ED1D4",
    x"BF6ED418",
    x"BF6ED65B",
    x"BF6ED89E",
    x"BF6EDAE1",
    x"BF6EDD23",
    x"BF6EDF66",
    x"BF6EE1A8",
    x"BF6EE3EA",
    x"BF6EE62C",
    x"BF6EE86E",
    x"BF6EEAB0",
    x"BF6EECF2",
    x"BF6EEF33",
    x"BF6EF175",
    x"BF6EF3B6",
    x"BF6EF5F7",
    x"BF6EF838",
    x"BF6EFA79",
    x"BF6EFCBA",
    x"BF6EFEFA",
    x"BF6F013A",
    x"BF6F037B",
    x"BF6F05BB",
    x"BF6F07FB",
    x"BF6F0A3A",
    x"BF6F0C7A",
    x"BF6F0EBA",
    x"BF6F10F9",
    x"BF6F1338",
    x"BF6F1577",
    x"BF6F17B6",
    x"BF6F19F5",
    x"BF6F1C34",
    x"BF6F1E72",
    x"BF6F20B0",
    x"BF6F22EF",
    x"BF6F252D",
    x"BF6F276B",
    x"BF6F29A8",
    x"BF6F2BE6",
    x"BF6F2E24",
    x"BF6F3061",
    x"BF6F329E",
    x"BF6F34DB",
    x"BF6F3718",
    x"BF6F3955",
    x"BF6F3B92",
    x"BF6F3DCE",
    x"BF6F400A",
    x"BF6F4247",
    x"BF6F4483",
    x"BF6F46BE",
    x"BF6F48FA",
    x"BF6F4B36",
    x"BF6F4D71",
    x"BF6F4FAD",
    x"BF6F51E8",
    x"BF6F5423",
    x"BF6F565E",
    x"BF6F5899",
    x"BF6F5AD3",
    x"BF6F5D0E",
    x"BF6F5F48",
    x"BF6F6182",
    x"BF6F63BC",
    x"BF6F65F6",
    x"BF6F6830",
    x"BF6F6A69",
    x"BF6F6CA3",
    x"BF6F6EDC",
    x"BF6F7115",
    x"BF6F734E",
    x"BF6F7587",
    x"BF6F77C0",
    x"BF6F79F8",
    x"BF6F7C31",
    x"BF6F7E69",
    x"BF6F80A1",
    x"BF6F82D9",
    x"BF6F8511",
    x"BF6F8749",
    x"BF6F8981",
    x"BF6F8BB8",
    x"BF6F8DEF",
    x"BF6F9026",
    x"BF6F925D",
    x"BF6F9494",
    x"BF6F96CB",
    x"BF6F9902",
    x"BF6F9B38",
    x"BF6F9D6E",
    x"BF6F9FA4",
    x"BF6FA1DA",
    x"BF6FA410",
    x"BF6FA646",
    x"BF6FA87C",
    x"BF6FAAB1",
    x"BF6FACE6",
    x"BF6FAF1B",
    x"BF6FB150",
    x"BF6FB385",
    x"BF6FB5BA",
    x"BF6FB7EE",
    x"BF6FBA23",
    x"BF6FBC57",
    x"BF6FBE8B",
    x"BF6FC0BF",
    x"BF6FC2F3",
    x"BF6FC527",
    x"BF6FC75A",
    x"BF6FC98E",
    x"BF6FCBC1",
    x"BF6FCDF4",
    x"BF6FD027",
    x"BF6FD25A",
    x"BF6FD48C",
    x"BF6FD6BF",
    x"BF6FD8F1",
    x"BF6FDB24",
    x"BF6FDD56",
    x"BF6FDF88",
    x"BF6FE1B9",
    x"BF6FE3EB",
    x"BF6FE61D",
    x"BF6FE84E",
    x"BF6FEA7F",
    x"BF6FECB0",
    x"BF6FEEE1",
    x"BF6FF112",
    x"BF6FF343",
    x"BF6FF573",
    x"BF6FF7A3",
    x"BF6FF9D4",
    x"BF6FFC04",
    x"BF6FFE34",
    x"BF700063",
    x"BF700293",
    x"BF7004C3",
    x"BF7006F2",
    x"BF700921",
    x"BF700B50",
    x"BF700D7F",
    x"BF700FAE",
    x"BF7011DC",
    x"BF70140B",
    x"BF701639",
    x"BF701867",
    x"BF701A95",
    x"BF701CC3",
    x"BF701EF1",
    x"BF70211F",
    x"BF70234C",
    x"BF70257A",
    x"BF7027A7",
    x"BF7029D4",
    x"BF702C01",
    x"BF702E2D",
    x"BF70305A",
    x"BF703286",
    x"BF7034B3",
    x"BF7036DF",
    x"BF70390B",
    x"BF703B37",
    x"BF703D63",
    x"BF703F8E",
    x"BF7041BA",
    x"BF7043E5",
    x"BF704610",
    x"BF70483B",
    x"BF704A66",
    x"BF704C91",
    x"BF704EBB",
    x"BF7050E6",
    x"BF705310",
    x"BF70553A",
    x"BF705764",
    x"BF70598E",
    x"BF705BB8",
    x"BF705DE1",
    x"BF70600A",
    x"BF706234",
    x"BF70645D",
    x"BF706686",
    x"BF7068AF",
    x"BF706AD7",
    x"BF706D00",
    x"BF706F28",
    x"BF707151",
    x"BF707379",
    x"BF7075A1",
    x"BF7077C8",
    x"BF7079F0",
    x"BF707C18",
    x"BF707E3F",
    x"BF708066",
    x"BF70828D",
    x"BF7084B4",
    x"BF7086DB",
    x"BF708902",
    x"BF708B28",
    x"BF708D4F",
    x"BF708F75",
    x"BF70919B",
    x"BF7093C1",
    x"BF7095E7",
    x"BF70980C",
    x"BF709A32",
    x"BF709C57",
    x"BF709E7C",
    x"BF70A0A2",
    x"BF70A2C6",
    x"BF70A4EB",
    x"BF70A710",
    x"BF70A934",
    x"BF70AB59",
    x"BF70AD7D",
    x"BF70AFA1",
    x"BF70B1C5",
    x"BF70B3E9",
    x"BF70B60C",
    x"BF70B830",
    x"BF70BA53",
    x"BF70BC76",
    x"BF70BE99",
    x"BF70C0BC",
    x"BF70C2DF",
    x"BF70C501",
    x"BF70C724",
    x"BF70C946",
    x"BF70CB68",
    x"BF70CD8A",
    x"BF70CFAC",
    x"BF70D1CE",
    x"BF70D3F0",
    x"BF70D611",
    x"BF70D832",
    x"BF70DA54",
    x"BF70DC75",
    x"BF70DE95",
    x"BF70E0B6",
    x"BF70E2D7",
    x"BF70E4F7",
    x"BF70E717",
    x"BF70E938",
    x"BF70EB58",
    x"BF70ED77",
    x"BF70EF97",
    x"BF70F1B7",
    x"BF70F3D6",
    x"BF70F5F5",
    x"BF70F814",
    x"BF70FA33",
    x"BF70FC52",
    x"BF70FE71",
    x"BF71008F",
    x"BF7102AE",
    x"BF7104CC",
    x"BF7106EA",
    x"BF710908",
    x"BF710B26",
    x"BF710D44",
    x"BF710F61",
    x"BF71117F",
    x"BF71139C",
    x"BF7115B9",
    x"BF7117D6",
    x"BF7119F3",
    x"BF711C0F",
    x"BF711E2C",
    x"BF712048",
    x"BF712264",
    x"BF712480",
    x"BF71269C",
    x"BF7128B8",
    x"BF712AD4",
    x"BF712CEF",
    x"BF712F0B",
    x"BF713126",
    x"BF713341",
    x"BF71355C",
    x"BF713776",
    x"BF713991",
    x"BF713BAC",
    x"BF713DC6",
    x"BF713FE0",
    x"BF7141FA",
    x"BF714414",
    x"BF71462E",
    x"BF714847",
    x"BF714A61",
    x"BF714C7A",
    x"BF714E93",
    x"BF7150AC",
    x"BF7152C5",
    x"BF7154DE",
    x"BF7156F6",
    x"BF71590F",
    x"BF715B27",
    x"BF715D3F",
    x"BF715F57",
    x"BF71616F",
    x"BF716387",
    x"BF71659F",
    x"BF7167B6",
    x"BF7169CD",
    x"BF716BE4",
    x"BF716DFB",
    x"BF717012",
    x"BF717229",
    x"BF71743F",
    x"BF717656",
    x"BF71786C",
    x"BF717A82",
    x"BF717C98",
    x"BF717EAE",
    x"BF7180C4",
    x"BF7182D9",
    x"BF7184EF",
    x"BF718704",
    x"BF718919",
    x"BF718B2E",
    x"BF718D43",
    x"BF718F57",
    x"BF71916C",
    x"BF719380",
    x"BF719594",
    x"BF7197A8",
    x"BF7199BC",
    x"BF719BD0",
    x"BF719DE4",
    x"BF719FF7",
    x"BF71A20B",
    x"BF71A41E",
    x"BF71A631",
    x"BF71A844",
    x"BF71AA57",
    x"BF71AC69",
    x"BF71AE7C",
    x"BF71B08E",
    x"BF71B2A0",
    x"BF71B4B2",
    x"BF71B6C4",
    x"BF71B8D6",
    x"BF71BAE7",
    x"BF71BCF9",
    x"BF71BF0A",
    x"BF71C11B",
    x"BF71C32C",
    x"BF71C53D",
    x"BF71C74E",
    x"BF71C95F",
    x"BF71CB6F",
    x"BF71CD7F",
    x"BF71CF8F",
    x"BF71D19F",
    x"BF71D3AF",
    x"BF71D5BF",
    x"BF71D7CF",
    x"BF71D9DE",
    x"BF71DBED",
    x"BF71DDFC",
    x"BF71E00B",
    x"BF71E21A",
    x"BF71E429",
    x"BF71E637",
    x"BF71E846",
    x"BF71EA54",
    x"BF71EC62",
    x"BF71EE70",
    x"BF71F07E",
    x"BF71F28C",
    x"BF71F499",
    x"BF71F6A6",
    x"BF71F8B4",
    x"BF71FAC1",
    x"BF71FCCE",
    x"BF71FEDA",
    x"BF7200E7",
    x"BF7202F4",
    x"BF720500",
    x"BF72070C",
    x"BF720918",
    x"BF720B24",
    x"BF720D30",
    x"BF720F3C",
    x"BF721147",
    x"BF721352",
    x"BF72155E",
    x"BF721769",
    x"BF721973",
    x"BF721B7E",
    x"BF721D89",
    x"BF721F93",
    x"BF72219E",
    x"BF7223A8",
    x"BF7225B2",
    x"BF7227BC",
    x"BF7229C5",
    x"BF722BCF",
    x"BF722DD8",
    x"BF722FE2",
    x"BF7231EB",
    x"BF7233F4",
    x"BF7235FD",
    x"BF723805",
    x"BF723A0E",
    x"BF723C16",
    x"BF723E1F",
    x"BF724027",
    x"BF72422F",
    x"BF724437",
    x"BF72463E",
    x"BF724846",
    x"BF724A4D",
    x"BF724C54",
    x"BF724E5C",
    x"BF725063",
    x"BF725269",
    x"BF725470",
    x"BF725677",
    x"BF72587D",
    x"BF725A83",
    x"BF725C89",
    x"BF725E8F",
    x"BF726095",
    x"BF72629B",
    x"BF7264A0",
    x"BF7266A5",
    x"BF7268AB",
    x"BF726AB0",
    x"BF726CB5",
    x"BF726EB9",
    x"BF7270BE",
    x"BF7272C2",
    x"BF7274C7",
    x"BF7276CB",
    x"BF7278CF",
    x"BF727AD3",
    x"BF727CD7",
    x"BF727EDA",
    x"BF7280DE",
    x"BF7282E1",
    x"BF7284E4",
    x"BF7286E7",
    x"BF7288EA",
    x"BF728AED",
    x"BF728CEF",
    x"BF728EF2",
    x"BF7290F4",
    x"BF7292F6",
    x"BF7294F8",
    x"BF7296FA",
    x"BF7298FC",
    x"BF729AFD",
    x"BF729CFF",
    x"BF729F00",
    x"BF72A101",
    x"BF72A302",
    x"BF72A503",
    x"BF72A703",
    x"BF72A904",
    x"BF72AB04",
    x"BF72AD05",
    x"BF72AF05",
    x"BF72B105",
    x"BF72B304",
    x"BF72B504",
    x"BF72B704",
    x"BF72B903",
    x"BF72BB02",
    x"BF72BD01",
    x"BF72BF00",
    x"BF72C0FF",
    x"BF72C2FE",
    x"BF72C4FC",
    x"BF72C6FA",
    x"BF72C8F9",
    x"BF72CAF7",
    x"BF72CCF5",
    x"BF72CEF2",
    x"BF72D0F0",
    x"BF72D2ED",
    x"BF72D4EB",
    x"BF72D6E8",
    x"BF72D8E5",
    x"BF72DAE2",
    x"BF72DCDE",
    x"BF72DEDB",
    x"BF72E0D7",
    x"BF72E2D4",
    x"BF72E4D0",
    x"BF72E6CC",
    x"BF72E8C8",
    x"BF72EAC3",
    x"BF72ECBF",
    x"BF72EEBA",
    x"BF72F0B6",
    x"BF72F2B1",
    x"BF72F4AC",
    x"BF72F6A7",
    x"BF72F8A1",
    x"BF72FA9C",
    x"BF72FC96",
    x"BF72FE90",
    x"BF73008B",
    x"BF730284",
    x"BF73047E",
    x"BF730678",
    x"BF730871",
    x"BF730A6B",
    x"BF730C64",
    x"BF730E5D",
    x"BF731056",
    x"BF73124F",
    x"BF731447",
    x"BF731640",
    x"BF731838",
    x"BF731A30",
    x"BF731C28",
    x"BF731E20",
    x"BF732018",
    x"BF732210",
    x"BF732407",
    x"BF7325FE",
    x"BF7327F6",
    x"BF7329ED",
    x"BF732BE4",
    x"BF732DDA",
    x"BF732FD1",
    x"BF7331C7",
    x"BF7333BE",
    x"BF7335B4",
    x"BF7337AA",
    x"BF7339A0",
    x"BF733B95",
    x"BF733D8B",
    x"BF733F80",
    x"BF734175",
    x"BF73436B",
    x"BF734560",
    x"BF734754",
    x"BF734949",
    x"BF734B3E",
    x"BF734D32",
    x"BF734F26",
    x"BF73511A",
    x"BF73530E",
    x"BF735502",
    x"BF7356F6",
    x"BF7358E9",
    x"BF735ADC",
    x"BF735CD0",
    x"BF735EC3",
    x"BF7360B6",
    x"BF7362A8",
    x"BF73649B",
    x"BF73668E",
    x"BF736880",
    x"BF736A72",
    x"BF736C64",
    x"BF736E56",
    x"BF737048",
    x"BF737239",
    x"BF73742B",
    x"BF73761C",
    x"BF73780D",
    x"BF7379FE",
    x"BF737BEF",
    x"BF737DE0",
    x"BF737FD0",
    x"BF7381C1",
    x"BF7383B1",
    x"BF7385A1",
    x"BF738791",
    x"BF738981",
    x"BF738B71",
    x"BF738D60",
    x"BF738F50",
    x"BF73913F",
    x"BF73932E",
    x"BF73951D",
    x"BF73970C",
    x"BF7398FA",
    x"BF739AE9",
    x"BF739CD7",
    x"BF739EC5",
    x"BF73A0B4",
    x"BF73A2A1",
    x"BF73A48F",
    x"BF73A67D",
    x"BF73A86A",
    x"BF73AA58",
    x"BF73AC45",
    x"BF73AE32",
    x"BF73B01F",
    x"BF73B20C",
    x"BF73B3F8",
    x"BF73B5E5",
    x"BF73B7D1",
    x"BF73B9BD",
    x"BF73BBA9",
    x"BF73BD95",
    x"BF73BF81",
    x"BF73C16C",
    x"BF73C358",
    x"BF73C543",
    x"BF73C72E",
    x"BF73C919",
    x"BF73CB04",
    x"BF73CCEF",
    x"BF73CED9",
    x"BF73D0C4",
    x"BF73D2AE",
    x"BF73D498",
    x"BF73D682",
    x"BF73D86C",
    x"BF73DA56",
    x"BF73DC3F",
    x"BF73DE28",
    x"BF73E012",
    x"BF73E1FB",
    x"BF73E3E4",
    x"BF73E5CC",
    x"BF73E7B5",
    x"BF73E99E",
    x"BF73EB86",
    x"BF73ED6E",
    x"BF73EF56",
    x"BF73F13E",
    x"BF73F326",
    x"BF73F50D",
    x"BF73F6F5",
    x"BF73F8DC",
    x"BF73FAC3",
    x"BF73FCAA",
    x"BF73FE91",
    x"BF740078",
    x"BF74025F",
    x"BF740445",
    x"BF74062B",
    x"BF740812",
    x"BF7409F8",
    x"BF740BDD",
    x"BF740DC3",
    x"BF740FA9",
    x"BF74118E",
    x"BF741373",
    x"BF741558",
    x"BF74173D",
    x"BF741922",
    x"BF741B07",
    x"BF741CEB",
    x"BF741ED0",
    x"BF7420B4",
    x"BF742298",
    x"BF74247C",
    x"BF742660",
    x"BF742843",
    x"BF742A27",
    x"BF742C0A",
    x"BF742DED",
    x"BF742FD1",
    x"BF7431B3",
    x"BF743396",
    x"BF743579",
    x"BF74375B",
    x"BF74393E",
    x"BF743B20",
    x"BF743D02",
    x"BF743EE4",
    x"BF7440C5",
    x"BF7442A7",
    x"BF744488",
    x"BF74466A",
    x"BF74484B",
    x"BF744A2C",
    x"BF744C0D",
    x"BF744DED",
    x"BF744FCE",
    x"BF7451AE",
    x"BF74538F",
    x"BF74556F",
    x"BF74574F",
    x"BF74592F",
    x"BF745B0E",
    x"BF745CEE",
    x"BF745ECD",
    x"BF7460AC",
    x"BF74628B",
    x"BF74646A",
    x"BF746649",
    x"BF746828",
    x"BF746A06",
    x"BF746BE5",
    x"BF746DC3",
    x"BF746FA1",
    x"BF74717F",
    x"BF74735D",
    x"BF74753A",
    x"BF747718",
    x"BF7478F5",
    x"BF747AD2",
    x"BF747CAF",
    x"BF747E8C",
    x"BF748069",
    x"BF748245",
    x"BF748422",
    x"BF7485FE",
    x"BF7487DA",
    x"BF7489B6",
    x"BF748B92",
    x"BF748D6E",
    x"BF748F49",
    x"BF749125",
    x"BF749300",
    x"BF7494DB",
    x"BF7496B6",
    x"BF749891",
    x"BF749A6B",
    x"BF749C46",
    x"BF749E20",
    x"BF749FFA",
    x"BF74A1D5",
    x"BF74A3AE",
    x"BF74A588",
    x"BF74A762",
    x"BF74A93B",
    x"BF74AB15",
    x"BF74ACEE",
    x"BF74AEC7",
    x"BF74B0A0",
    x"BF74B279",
    x"BF74B451",
    x"BF74B62A",
    x"BF74B802",
    x"BF74B9DA",
    x"BF74BBB2",
    x"BF74BD8A",
    x"BF74BF62",
    x"BF74C139",
    x"BF74C311",
    x"BF74C4E8",
    x"BF74C6BF",
    x"BF74C896",
    x"BF74CA6D",
    x"BF74CC44",
    x"BF74CE1A",
    x"BF74CFF0",
    x"BF74D1C7",
    x"BF74D39D",
    x"BF74D573",
    x"BF74D749",
    x"BF74D91E",
    x"BF74DAF4",
    x"BF74DCC9",
    x"BF74DE9E",
    x"BF74E073",
    x"BF74E248",
    x"BF74E41D",
    x"BF74E5F2",
    x"BF74E7C6",
    x"BF74E99A",
    x"BF74EB6F",
    x"BF74ED43",
    x"BF74EF17",
    x"BF74F0EA",
    x"BF74F2BE",
    x"BF74F491",
    x"BF74F665",
    x"BF74F838",
    x"BF74FA0B",
    x"BF74FBDE",
    x"BF74FDB0",
    x"BF74FF83",
    x"BF750155",
    x"BF750327",
    x"BF7504FA",
    x"BF7506CC",
    x"BF75089D",
    x"BF750A6F",
    x"BF750C41",
    x"BF750E12",
    x"BF750FE3",
    x"BF7511B4",
    x"BF751385",
    x"BF751556",
    x"BF751727",
    x"BF7518F7",
    x"BF751AC7",
    x"BF751C98",
    x"BF751E68",
    x"BF752038",
    x"BF752207",
    x"BF7523D7",
    x"BF7525A6",
    x"BF752776",
    x"BF752945",
    x"BF752B14",
    x"BF752CE3",
    x"BF752EB1",
    x"BF753080",
    x"BF75324E",
    x"BF75341D",
    x"BF7535EB",
    x"BF7537B9",
    x"BF753987",
    x"BF753B54",
    x"BF753D22",
    x"BF753EEF",
    x"BF7540BC",
    x"BF754289",
    x"BF754456",
    x"BF754623",
    x"BF7547F0",
    x"BF7549BC",
    x"BF754B89",
    x"BF754D55",
    x"BF754F21",
    x"BF7550ED",
    x"BF7552B9",
    x"BF755484",
    x"BF755650",
    x"BF75581B",
    x"BF7559E6",
    x"BF755BB1",
    x"BF755D7C",
    x"BF755F47",
    x"BF756111",
    x"BF7562DC",
    x"BF7564A6",
    x"BF756670",
    x"BF75683A",
    x"BF756A04",
    x"BF756BCE",
    x"BF756D97",
    x"BF756F61",
    x"BF75712A",
    x"BF7572F3",
    x"BF7574BC",
    x"BF757685",
    x"BF75784D",
    x"BF757A16",
    x"BF757BDE",
    x"BF757DA7",
    x"BF757F6F",
    x"BF758136",
    x"BF7582FE",
    x"BF7584C6",
    x"BF75868D",
    x"BF758855",
    x"BF758A1C",
    x"BF758BE3",
    x"BF758DAA",
    x"BF758F70",
    x"BF759137",
    x"BF7592FE",
    x"BF7594C4",
    x"BF75968A",
    x"BF759850",
    x"BF759A16",
    x"BF759BDB",
    x"BF759DA1",
    x"BF759F66",
    x"BF75A12C",
    x"BF75A2F1",
    x"BF75A4B6",
    x"BF75A67B",
    x"BF75A83F",
    x"BF75AA04",
    x"BF75ABC8",
    x"BF75AD8C",
    x"BF75AF50",
    x"BF75B114",
    x"BF75B2D8",
    x"BF75B49C",
    x"BF75B65F",
    x"BF75B822",
    x"BF75B9E6",
    x"BF75BBA9",
    x"BF75BD6C",
    x"BF75BF2E",
    x"BF75C0F1",
    x"BF75C2B3",
    x"BF75C476",
    x"BF75C638",
    x"BF75C7FA",
    x"BF75C9BC",
    x"BF75CB7D",
    x"BF75CD3F",
    x"BF75CF00",
    x"BF75D0C2",
    x"BF75D283",
    x"BF75D444",
    x"BF75D604",
    x"BF75D7C5",
    x"BF75D986",
    x"BF75DB46",
    x"BF75DD06",
    x"BF75DEC6",
    x"BF75E086",
    x"BF75E246",
    x"BF75E406",
    x"BF75E5C5",
    x"BF75E784",
    x"BF75E944",
    x"BF75EB03",
    x"BF75ECC2",
    x"BF75EE80",
    x"BF75F03F",
    x"BF75F1FD",
    x"BF75F3BC",
    x"BF75F57A",
    x"BF75F738",
    x"BF75F8F6",
    x"BF75FAB3",
    x"BF75FC71",
    x"BF75FE2E",
    x"BF75FFEB",
    x"BF7601A9",
    x"BF760366",
    x"BF760522",
    x"BF7606DF",
    x"BF76089C",
    x"BF760A58",
    x"BF760C14",
    x"BF760DD0",
    x"BF760F8C",
    x"BF761148",
    x"BF761304",
    x"BF7614BF",
    x"BF76167A",
    x"BF761836",
    x"BF7619F1",
    x"BF761BAB",
    x"BF761D66",
    x"BF761F21",
    x"BF7620DB",
    x"BF762296",
    x"BF762450",
    x"BF76260A",
    x"BF7627C3",
    x"BF76297D",
    x"BF762B37",
    x"BF762CF0",
    x"BF762EA9",
    x"BF763063",
    x"BF76321B",
    x"BF7633D4",
    x"BF76358D",
    x"BF763745",
    x"BF7638FE",
    x"BF763AB6",
    x"BF763C6E",
    x"BF763E26",
    x"BF763FDE",
    x"BF764195",
    x"BF76434D",
    x"BF764504",
    x"BF7646BB",
    x"BF764872",
    x"BF764A29",
    x"BF764BE0",
    x"BF764D97",
    x"BF764F4D",
    x"BF765103",
    x"BF7652B9",
    x"BF76546F",
    x"BF765625",
    x"BF7657DB",
    x"BF765991",
    x"BF765B46",
    x"BF765CFB",
    x"BF765EB0",
    x"BF766065",
    x"BF76621A",
    x"BF7663CF",
    x"BF766583",
    x"BF766738",
    x"BF7668EC",
    x"BF766AA0",
    x"BF766C54",
    x"BF766E08",
    x"BF766FBB",
    x"BF76716F",
    x"BF767322",
    x"BF7674D5",
    x"BF767688",
    x"BF76783B",
    x"BF7679EE",
    x"BF767BA0",
    x"BF767D53",
    x"BF767F05",
    x"BF7680B7",
    x"BF768269",
    x"BF76841B",
    x"BF7685CD",
    x"BF76877E",
    x"BF768930",
    x"BF768AE1",
    x"BF768C92",
    x"BF768E43",
    x"BF768FF4",
    x"BF7691A4",
    x"BF769355",
    x"BF769505",
    x"BF7696B5",
    x"BF769865",
    x"BF769A15",
    x"BF769BC5",
    x"BF769D75",
    x"BF769F24",
    x"BF76A0D3",
    x"BF76A283",
    x"BF76A432",
    x"BF76A5E0",
    x"BF76A78F",
    x"BF76A93E",
    x"BF76AAEC",
    x"BF76AC9A",
    x"BF76AE49",
    x"BF76AFF7",
    x"BF76B1A4",
    x"BF76B352",
    x"BF76B500",
    x"BF76B6AD",
    x"BF76B85A",
    x"BF76BA07",
    x"BF76BBB4",
    x"BF76BD61",
    x"BF76BF0E",
    x"BF76C0BA",
    x"BF76C266",
    x"BF76C413",
    x"BF76C5BF",
    x"BF76C76B",
    x"BF76C916",
    x"BF76CAC2",
    x"BF76CC6D",
    x"BF76CE19",
    x"BF76CFC4",
    x"BF76D16F",
    x"BF76D31A",
    x"BF76D4C4",
    x"BF76D66F",
    x"BF76D819",
    x"BF76D9C4",
    x"BF76DB6E",
    x"BF76DD18",
    x"BF76DEC1",
    x"BF76E06B",
    x"BF76E215",
    x"BF76E3BE",
    x"BF76E567",
    x"BF76E710",
    x"BF76E8B9",
    x"BF76EA62",
    x"BF76EC0B",
    x"BF76EDB3",
    x"BF76EF5B",
    x"BF76F103",
    x"BF76F2AC",
    x"BF76F453",
    x"BF76F5FB",
    x"BF76F7A3",
    x"BF76F94A",
    x"BF76FAF1",
    x"BF76FC99",
    x"BF76FE40",
    x"BF76FFE6",
    x"BF77018D",
    x"BF770334",
    x"BF7704DA",
    x"BF770680",
    x"BF770826",
    x"BF7709CC",
    x"BF770B72",
    x"BF770D18",
    x"BF770EBD",
    x"BF771063",
    x"BF771208",
    x"BF7713AD",
    x"BF771552",
    x"BF7716F6",
    x"BF77189B",
    x"BF771A3F",
    x"BF771BE4",
    x"BF771D88",
    x"BF771F2C",
    x"BF7720D0",
    x"BF772274",
    x"BF772417",
    x"BF7725BA",
    x"BF77275E",
    x"BF772901",
    x"BF772AA4",
    x"BF772C47",
    x"BF772DE9",
    x"BF772F8C",
    x"BF77312E",
    x"BF7732D0",
    x"BF773472",
    x"BF773614",
    x"BF7737B6",
    x"BF773958",
    x"BF773AF9",
    x"BF773C9B",
    x"BF773E3C",
    x"BF773FDD",
    x"BF77417E",
    x"BF77431E",
    x"BF7744BF",
    x"BF77465F",
    x"BF774800",
    x"BF7749A0",
    x"BF774B40",
    x"BF774CE0",
    x"BF774E7F",
    x"BF77501F",
    x"BF7751BE",
    x"BF77535E",
    x"BF7754FD",
    x"BF77569C",
    x"BF77583A",
    x"BF7759D9",
    x"BF775B78",
    x"BF775D16",
    x"BF775EB4",
    x"BF776052",
    x"BF7761F0",
    x"BF77638E",
    x"BF77652B",
    x"BF7766C9",
    x"BF776866",
    x"BF776A03",
    x"BF776BA0",
    x"BF776D3D",
    x"BF776EDA",
    x"BF777076",
    x"BF777213",
    x"BF7773AF",
    x"BF77754B",
    x"BF7776E7",
    x"BF777883",
    x"BF777A1F",
    x"BF777BBA",
    x"BF777D56",
    x"BF777EF1",
    x"BF77808C",
    x"BF778227",
    x"BF7783C2",
    x"BF77855C",
    x"BF7786F7",
    x"BF778891",
    x"BF778A2B",
    x"BF778BC5",
    x"BF778D5F",
    x"BF778EF9",
    x"BF779092",
    x"BF77922C",
    x"BF7793C5",
    x"BF77955E",
    x"BF7796F7",
    x"BF779890",
    x"BF779A29",
    x"BF779BC1",
    x"BF779D5A",
    x"BF779EF2",
    x"BF77A08A",
    x"BF77A222",
    x"BF77A3BA",
    x"BF77A551",
    x"BF77A6E9",
    x"BF77A880",
    x"BF77AA17",
    x"BF77ABAE",
    x"BF77AD45",
    x"BF77AEDC",
    x"BF77B073",
    x"BF77B209",
    x"BF77B39F",
    x"BF77B535",
    x"BF77B6CB",
    x"BF77B861",
    x"BF77B9F7",
    x"BF77BB8D",
    x"BF77BD22",
    x"BF77BEB7",
    x"BF77C04C",
    x"BF77C1E1",
    x"BF77C376",
    x"BF77C50B",
    x"BF77C69F",
    x"BF77C834",
    x"BF77C9C8",
    x"BF77CB5C",
    x"BF77CCF0",
    x"BF77CE83",
    x"BF77D017",
    x"BF77D1AB",
    x"BF77D33E",
    x"BF77D4D1",
    x"BF77D664",
    x"BF77D7F7",
    x"BF77D98A",
    x"BF77DB1C",
    x"BF77DCAF",
    x"BF77DE41",
    x"BF77DFD3",
    x"BF77E165",
    x"BF77E2F7",
    x"BF77E488",
    x"BF77E61A",
    x"BF77E7AB",
    x"BF77E93D",
    x"BF77EACE",
    x"BF77EC5F",
    x"BF77EDEF",
    x"BF77EF80",
    x"BF77F110",
    x"BF77F2A1",
    x"BF77F431",
    x"BF77F5C1",
    x"BF77F751",
    x"BF77F8E1",
    x"BF77FA70",
    x"BF77FC00",
    x"BF77FD8F",
    x"BF77FF1E",
    x"BF7800AD",
    x"BF78023C",
    x"BF7803CA",
    x"BF780559",
    x"BF7806E7",
    x"BF780876",
    x"BF780A04",
    x"BF780B92",
    x"BF780D1F",
    x"BF780EAD",
    x"BF78103A",
    x"BF7811C8",
    x"BF781355",
    x"BF7814E2",
    x"BF78166F",
    x"BF7817FC",
    x"BF781988",
    x"BF781B15",
    x"BF781CA1",
    x"BF781E2D",
    x"BF781FB9",
    x"BF782145",
    x"BF7822D1",
    x"BF78245C",
    x"BF7825E8",
    x"BF782773",
    x"BF7828FE",
    x"BF782A89",
    x"BF782C14",
    x"BF782D9E",
    x"BF782F29",
    x"BF7830B3",
    x"BF78323D",
    x"BF7833C7",
    x"BF783551",
    x"BF7836DB",
    x"BF783865",
    x"BF7839EE",
    x"BF783B77",
    x"BF783D01",
    x"BF783E8A",
    x"BF784012",
    x"BF78419B",
    x"BF784324",
    x"BF7844AC",
    x"BF784634",
    x"BF7847BC",
    x"BF784944",
    x"BF784ACC",
    x"BF784C54",
    x"BF784DDB",
    x"BF784F63",
    x"BF7850EA",
    x"BF785271",
    x"BF7853F8",
    x"BF78557F",
    x"BF785705",
    x"BF78588C",
    x"BF785A12",
    x"BF785B98",
    x"BF785D1E",
    x"BF785EA4",
    x"BF78602A",
    x"BF7861AF",
    x"BF786335",
    x"BF7864BA",
    x"BF78663F",
    x"BF7867C4",
    x"BF786949",
    x"BF786ACE",
    x"BF786C52",
    x"BF786DD6",
    x"BF786F5B",
    x"BF7870DF",
    x"BF787263",
    x"BF7873E6",
    x"BF78756A",
    x"BF7876ED",
    x"BF787871",
    x"BF7879F4",
    x"BF787B77",
    x"BF787CFA",
    x"BF787E7D",
    x"BF787FFF",
    x"BF788182",
    x"BF788304",
    x"BF788486",
    x"BF788608",
    x"BF78878A",
    x"BF78890B",
    x"BF788A8D",
    x"BF788C0E",
    x"BF788D8F",
    x"BF788F11",
    x"BF789091",
    x"BF789212",
    x"BF789393",
    x"BF789513",
    x"BF789694",
    x"BF789814",
    x"BF789994",
    x"BF789B14",
    x"BF789C93",
    x"BF789E13",
    x"BF789F92",
    x"BF78A112",
    x"BF78A291",
    x"BF78A410",
    x"BF78A58F",
    x"BF78A70D",
    x"BF78A88C",
    x"BF78AA0A",
    x"BF78AB88",
    x"BF78AD06",
    x"BF78AE84",
    x"BF78B002",
    x"BF78B180",
    x"BF78B2FD",
    x"BF78B47B",
    x"BF78B5F8",
    x"BF78B775",
    x"BF78B8F2",
    x"BF78BA6E",
    x"BF78BBEB",
    x"BF78BD67",
    x"BF78BEE4",
    x"BF78C060",
    x"BF78C1DC",
    x"BF78C358",
    x"BF78C4D3",
    x"BF78C64F",
    x"BF78C7CA",
    x"BF78C945",
    x"BF78CAC1",
    x"BF78CC3B",
    x"BF78CDB6",
    x"BF78CF31",
    x"BF78D0AB",
    x"BF78D226",
    x"BF78D3A0",
    x"BF78D51A",
    x"BF78D694",
    x"BF78D80E",
    x"BF78D987",
    x"BF78DB01",
    x"BF78DC7A",
    x"BF78DDF3",
    x"BF78DF6C",
    x"BF78E0E5",
    x"BF78E25D",
    x"BF78E3D6",
    x"BF78E54E",
    x"BF78E6C7",
    x"BF78E83F",
    x"BF78E9B7",
    x"BF78EB2E",
    x"BF78ECA6",
    x"BF78EE1D",
    x"BF78EF95",
    x"BF78F10C",
    x"BF78F283",
    x"BF78F3FA",
    x"BF78F571",
    x"BF78F6E7",
    x"BF78F85E",
    x"BF78F9D4",
    x"BF78FB4A",
    x"BF78FCC0",
    x"BF78FE36",
    x"BF78FFAC",
    x"BF790121",
    x"BF790296",
    x"BF79040C",
    x"BF790581",
    x"BF7906F6",
    x"BF79086A",
    x"BF7909DF",
    x"BF790B54",
    x"BF790CC8",
    x"BF790E3C",
    x"BF790FB0",
    x"BF791124",
    x"BF791298",
    x"BF79140B",
    x"BF79157F",
    x"BF7916F2",
    x"BF791865",
    x"BF7919D8",
    x"BF791B4B",
    x"BF791CBE",
    x"BF791E30",
    x"BF791FA3",
    x"BF792115",
    x"BF792287",
    x"BF7923F9",
    x"BF79256B",
    x"BF7926DC",
    x"BF79284E",
    x"BF7929BF",
    x"BF792B30",
    x"BF792CA1",
    x"BF792E12",
    x"BF792F83",
    x"BF7930F3",
    x"BF793264",
    x"BF7933D4",
    x"BF793544",
    x"BF7936B4",
    x"BF793824",
    x"BF793994",
    x"BF793B03",
    x"BF793C73",
    x"BF793DE2",
    x"BF793F51",
    x"BF7940C0",
    x"BF79422F",
    x"BF79439D",
    x"BF79450C",
    x"BF79467A",
    x"BF7947E8",
    x"BF794956",
    x"BF794AC4",
    x"BF794C32",
    x"BF794D9F",
    x"BF794F0D",
    x"BF79507A",
    x"BF7951E7",
    x"BF795354",
    x"BF7954C1",
    x"BF79562E",
    x"BF79579A",
    x"BF795907",
    x"BF795A73",
    x"BF795BDF",
    x"BF795D4B",
    x"BF795EB7",
    x"BF796022",
    x"BF79618E",
    x"BF7962F9",
    x"BF796464",
    x"BF7965CF",
    x"BF79673A",
    x"BF7968A5",
    x"BF796A0F",
    x"BF796B7A",
    x"BF796CE4",
    x"BF796E4E",
    x"BF796FB8",
    x"BF797122",
    x"BF79728C",
    x"BF7973F5",
    x"BF79755F",
    x"BF7976C8",
    x"BF797831",
    x"BF79799A",
    x"BF797B03",
    x"BF797C6B",
    x"BF797DD4",
    x"BF797F3C",
    x"BF7980A4",
    x"BF79820C",
    x"BF798374",
    x"BF7984DC",
    x"BF798643",
    x"BF7987AB",
    x"BF798912",
    x"BF798A79",
    x"BF798BE0",
    x"BF798D47",
    x"BF798EAE",
    x"BF799014",
    x"BF79917A",
    x"BF7992E1",
    x"BF799447",
    x"BF7995AD",
    x"BF799712",
    x"BF799878",
    x"BF7999DE",
    x"BF799B43",
    x"BF799CA8",
    x"BF799E0D",
    x"BF799F72",
    x"BF79A0D7",
    x"BF79A23B",
    x"BF79A3A0",
    x"BF79A504",
    x"BF79A668",
    x"BF79A7CC",
    x"BF79A930",
    x"BF79AA93",
    x"BF79ABF7",
    x"BF79AD5A",
    x"BF79AEBD",
    x"BF79B020",
    x"BF79B183",
    x"BF79B2E6",
    x"BF79B449",
    x"BF79B5AB",
    x"BF79B70D",
    x"BF79B870",
    x"BF79B9D2",
    x"BF79BB33",
    x"BF79BC95",
    x"BF79BDF7",
    x"BF79BF58",
    x"BF79C0B9",
    x"BF79C21A",
    x"BF79C37B",
    x"BF79C4DC",
    x"BF79C63D",
    x"BF79C79D",
    x"BF79C8FE",
    x"BF79CA5E",
    x"BF79CBBE",
    x"BF79CD1E",
    x"BF79CE7E",
    x"BF79CFDD",
    x"BF79D13D",
    x"BF79D29C",
    x"BF79D3FB",
    x"BF79D55A",
    x"BF79D6B9",
    x"BF79D818",
    x"BF79D976",
    x"BF79DAD5",
    x"BF79DC33",
    x"BF79DD91",
    x"BF79DEEF",
    x"BF79E04D",
    x"BF79E1AA",
    x"BF79E308",
    x"BF79E465",
    x"BF79E5C2",
    x"BF79E71F",
    x"BF79E87C",
    x"BF79E9D9",
    x"BF79EB36",
    x"BF79EC92",
    x"BF79EDEE",
    x"BF79EF4A",
    x"BF79F0A6",
    x"BF79F202",
    x"BF79F35E",
    x"BF79F4B9",
    x"BF79F615",
    x"BF79F770",
    x"BF79F8CB",
    x"BF79FA26",
    x"BF79FB81",
    x"BF79FCDB",
    x"BF79FE36",
    x"BF79FF90",
    x"BF7A00EA",
    x"BF7A0244",
    x"BF7A039E",
    x"BF7A04F8",
    x"BF7A0652",
    x"BF7A07AB",
    x"BF7A0904",
    x"BF7A0A5D",
    x"BF7A0BB6",
    x"BF7A0D0F",
    x"BF7A0E68",
    x"BF7A0FC0",
    x"BF7A1119",
    x"BF7A1271",
    x"BF7A13C9",
    x"BF7A1521",
    x"BF7A1679",
    x"BF7A17D0",
    x"BF7A1928",
    x"BF7A1A7F",
    x"BF7A1BD6",
    x"BF7A1D2D",
    x"BF7A1E84",
    x"BF7A1FDB",
    x"BF7A2131",
    x"BF7A2288",
    x"BF7A23DE",
    x"BF7A2534",
    x"BF7A268A",
    x"BF7A27E0",
    x"BF7A2936",
    x"BF7A2A8B",
    x"BF7A2BE1",
    x"BF7A2D36",
    x"BF7A2E8B",
    x"BF7A2FE0",
    x"BF7A3134",
    x"BF7A3289",
    x"BF7A33DD",
    x"BF7A3532",
    x"BF7A3686",
    x"BF7A37DA",
    x"BF7A392E",
    x"BF7A3A81",
    x"BF7A3BD5",
    x"BF7A3D28",
    x"BF7A3E7C",
    x"BF7A3FCF",
    x"BF7A4122",
    x"BF7A4275",
    x"BF7A43C7",
    x"BF7A451A",
    x"BF7A466C",
    x"BF7A47BE",
    x"BF7A4910",
    x"BF7A4A62",
    x"BF7A4BB4",
    x"BF7A4D05",
    x"BF7A4E57",
    x"BF7A4FA8",
    x"BF7A50F9",
    x"BF7A524A",
    x"BF7A539B",
    x"BF7A54EC",
    x"BF7A563C",
    x"BF7A578D",
    x"BF7A58DD",
    x"BF7A5A2D",
    x"BF7A5B7D",
    x"BF7A5CCD",
    x"BF7A5E1C",
    x"BF7A5F6C",
    x"BF7A60BB",
    x"BF7A620A",
    x"BF7A6359",
    x"BF7A64A8",
    x"BF7A65F7",
    x"BF7A6745",
    x"BF7A6894",
    x"BF7A69E2",
    x"BF7A6B30",
    x"BF7A6C7E",
    x"BF7A6DCC",
    x"BF7A6F1A",
    x"BF7A7067",
    x"BF7A71B5",
    x"BF7A7302",
    x"BF7A744F",
    x"BF7A759C",
    x"BF7A76E9",
    x"BF7A7835",
    x"BF7A7982",
    x"BF7A7ACE",
    x"BF7A7C1A",
    x"BF7A7D66",
    x"BF7A7EB2",
    x"BF7A7FFE",
    x"BF7A8149",
    x"BF7A8295",
    x"BF7A83E0",
    x"BF7A852B",
    x"BF7A8676",
    x"BF7A87C1",
    x"BF7A890B",
    x"BF7A8A56",
    x"BF7A8BA0",
    x"BF7A8CEA",
    x"BF7A8E34",
    x"BF7A8F7E",
    x"BF7A90C8",
    x"BF7A9212",
    x"BF7A935B",
    x"BF7A94A4",
    x"BF7A95EE",
    x"BF7A9737",
    x"BF7A987F",
    x"BF7A99C8",
    x"BF7A9B11",
    x"BF7A9C59",
    x"BF7A9DA1",
    x"BF7A9EE9",
    x"BF7AA031",
    x"BF7AA179",
    x"BF7AA2C1",
    x"BF7AA408",
    x"BF7AA54F",
    x"BF7AA697",
    x"BF7AA7DE",
    x"BF7AA925",
    x"BF7AAA6B",
    x"BF7AABB2",
    x"BF7AACF8",
    x"BF7AAE3F",
    x"BF7AAF85",
    x"BF7AB0CB",
    x"BF7AB210",
    x"BF7AB356",
    x"BF7AB49C",
    x"BF7AB5E1",
    x"BF7AB726",
    x"BF7AB86B",
    x"BF7AB9B0",
    x"BF7ABAF5",
    x"BF7ABC3A",
    x"BF7ABD7E",
    x"BF7ABEC2",
    x"BF7AC006",
    x"BF7AC14A",
    x"BF7AC28E",
    x"BF7AC3D2",
    x"BF7AC516",
    x"BF7AC659",
    x"BF7AC79C",
    x"BF7AC8DF",
    x"BF7ACA22",
    x"BF7ACB65",
    x"BF7ACCA8",
    x"BF7ACDEA",
    x"BF7ACF2D",
    x"BF7AD06F",
    x"BF7AD1B1",
    x"BF7AD2F3",
    x"BF7AD434",
    x"BF7AD576",
    x"BF7AD6B7",
    x"BF7AD7F9",
    x"BF7AD93A",
    x"BF7ADA7B",
    x"BF7ADBBC",
    x"BF7ADCFC",
    x"BF7ADE3D",
    x"BF7ADF7D",
    x"BF7AE0BD",
    x"BF7AE1FE",
    x"BF7AE33D",
    x"BF7AE47D",
    x"BF7AE5BD",
    x"BF7AE6FC",
    x"BF7AE83C",
    x"BF7AE97B",
    x"BF7AEABA",
    x"BF7AEBF9",
    x"BF7AED37",
    x"BF7AEE76",
    x"BF7AEFB4",
    x"BF7AF0F3",
    x"BF7AF231",
    x"BF7AF36F",
    x"BF7AF4AD",
    x"BF7AF5EA",
    x"BF7AF728",
    x"BF7AF865",
    x"BF7AF9A2",
    x"BF7AFADF",
    x"BF7AFC1C",
    x"BF7AFD59",
    x"BF7AFE96",
    x"BF7AFFD2",
    x"BF7B010E",
    x"BF7B024A",
    x"BF7B0386",
    x"BF7B04C2",
    x"BF7B05FE",
    x"BF7B073A",
    x"BF7B0875",
    x"BF7B09B0",
    x"BF7B0AEB",
    x"BF7B0C26",
    x"BF7B0D61",
    x"BF7B0E9C",
    x"BF7B0FD6",
    x"BF7B1110",
    x"BF7B124B",
    x"BF7B1385",
    x"BF7B14BE",
    x"BF7B15F8",
    x"BF7B1732",
    x"BF7B186B",
    x"BF7B19A4",
    x"BF7B1ADE",
    x"BF7B1C17",
    x"BF7B1D4F",
    x"BF7B1E88",
    x"BF7B1FC1",
    x"BF7B20F9",
    x"BF7B2231",
    x"BF7B2369",
    x"BF7B24A1",
    x"BF7B25D9",
    x"BF7B2711",
    x"BF7B2848",
    x"BF7B297F",
    x"BF7B2AB6",
    x"BF7B2BED",
    x"BF7B2D24",
    x"BF7B2E5B",
    x"BF7B2F92",
    x"BF7B30C8",
    x"BF7B31FE",
    x"BF7B3334",
    x"BF7B346A",
    x"BF7B35A0",
    x"BF7B36D6",
    x"BF7B380B",
    x"BF7B3940",
    x"BF7B3A76",
    x"BF7B3BAB",
    x"BF7B3CE0",
    x"BF7B3E14",
    x"BF7B3F49",
    x"BF7B407D",
    x"BF7B41B2",
    x"BF7B42E6",
    x"BF7B441A",
    x"BF7B454E",
    x"BF7B4681",
    x"BF7B47B5",
    x"BF7B48E8",
    x"BF7B4A1B",
    x"BF7B4B4E",
    x"BF7B4C81",
    x"BF7B4DB4",
    x"BF7B4EE7",
    x"BF7B5019",
    x"BF7B514B",
    x"BF7B527E",
    x"BF7B53B0",
    x"BF7B54E1",
    x"BF7B5613",
    x"BF7B5745",
    x"BF7B5876",
    x"BF7B59A7",
    x"BF7B5AD9",
    x"BF7B5C09",
    x"BF7B5D3A",
    x"BF7B5E6B",
    x"BF7B5F9B",
    x"BF7B60CC",
    x"BF7B61FC",
    x"BF7B632C",
    x"BF7B645C",
    x"BF7B658C",
    x"BF7B66BB",
    x"BF7B67EB",
    x"BF7B691A",
    x"BF7B6A49",
    x"BF7B6B78",
    x"BF7B6CA7",
    x"BF7B6DD6",
    x"BF7B6F04",
    x"BF7B7032",
    x"BF7B7161",
    x"BF7B728F",
    x"BF7B73BD",
    x"BF7B74EA",
    x"BF7B7618",
    x"BF7B7745",
    x"BF7B7873",
    x"BF7B79A0",
    x"BF7B7ACD",
    x"BF7B7BFA",
    x"BF7B7D27",
    x"BF7B7E53",
    x"BF7B7F80",
    x"BF7B80AC",
    x"BF7B81D8",
    x"BF7B8304",
    x"BF7B8430",
    x"BF7B855B",
    x"BF7B8687",
    x"BF7B87B2",
    x"BF7B88DD",
    x"BF7B8A08",
    x"BF7B8B33",
    x"BF7B8C5E",
    x"BF7B8D89",
    x"BF7B8EB3",
    x"BF7B8FDD",
    x"BF7B9107",
    x"BF7B9231",
    x"BF7B935B",
    x"BF7B9485",
    x"BF7B95AE",
    x"BF7B96D8",
    x"BF7B9801",
    x"BF7B992A",
    x"BF7B9A53",
    x"BF7B9B7C",
    x"BF7B9CA4",
    x"BF7B9DCD",
    x"BF7B9EF5",
    x"BF7BA01D",
    x"BF7BA145",
    x"BF7BA26D",
    x"BF7BA395",
    x"BF7BA4BC",
    x"BF7BA5E4",
    x"BF7BA70B",
    x"BF7BA832",
    x"BF7BA959",
    x"BF7BAA80",
    x"BF7BABA7",
    x"BF7BACCD",
    x"BF7BADF3",
    x"BF7BAF1A",
    x"BF7BB040",
    x"BF7BB166",
    x"BF7BB28B",
    x"BF7BB3B1",
    x"BF7BB4D6",
    x"BF7BB5FC",
    x"BF7BB721",
    x"BF7BB846",
    x"BF7BB96B",
    x"BF7BBA8F",
    x"BF7BBBB4",
    x"BF7BBCD8",
    x"BF7BBDFC",
    x"BF7BBF20",
    x"BF7BC044",
    x"BF7BC168",
    x"BF7BC28C",
    x"BF7BC3AF",
    x"BF7BC4D2",
    x"BF7BC5F6",
    x"BF7BC719",
    x"BF7BC83B",
    x"BF7BC95E",
    x"BF7BCA81",
    x"BF7BCBA3",
    x"BF7BCCC5",
    x"BF7BCDE7",
    x"BF7BCF09",
    x"BF7BD02B",
    x"BF7BD14D",
    x"BF7BD26E",
    x"BF7BD390",
    x"BF7BD4B1",
    x"BF7BD5D2",
    x"BF7BD6F3",
    x"BF7BD814",
    x"BF7BD934",
    x"BF7BDA55",
    x"BF7BDB75",
    x"BF7BDC95",
    x"BF7BDDB5",
    x"BF7BDED5",
    x"BF7BDFF4",
    x"BF7BE114",
    x"BF7BE233",
    x"BF7BE353",
    x"BF7BE472",
    x"BF7BE590",
    x"BF7BE6AF",
    x"BF7BE7CE",
    x"BF7BE8EC",
    x"BF7BEA0B",
    x"BF7BEB29",
    x"BF7BEC47",
    x"BF7BED65",
    x"BF7BEE82",
    x"BF7BEFA0",
    x"BF7BF0BD",
    x"BF7BF1DA",
    x"BF7BF2F8",
    x"BF7BF415",
    x"BF7BF531",
    x"BF7BF64E",
    x"BF7BF76A",
    x"BF7BF887",
    x"BF7BF9A3",
    x"BF7BFABF",
    x"BF7BFBDB",
    x"BF7BFCF7",
    x"BF7BFE12",
    x"BF7BFF2E",
    x"BF7C0049",
    x"BF7C0164",
    x"BF7C027F",
    x"BF7C039A",
    x"BF7C04B4",
    x"BF7C05CF",
    x"BF7C06E9",
    x"BF7C0803",
    x"BF7C091E",
    x"BF7C0A37",
    x"BF7C0B51",
    x"BF7C0C6B",
    x"BF7C0D84",
    x"BF7C0E9D",
    x"BF7C0FB7",
    x"BF7C10D0",
    x"BF7C11E8",
    x"BF7C1301",
    x"BF7C141A",
    x"BF7C1532",
    x"BF7C164A",
    x"BF7C1762",
    x"BF7C187A",
    x"BF7C1992",
    x"BF7C1AAA",
    x"BF7C1BC1",
    x"BF7C1CD9",
    x"BF7C1DF0",
    x"BF7C1F07",
    x"BF7C201E",
    x"BF7C2134",
    x"BF7C224B",
    x"BF7C2361",
    x"BF7C2478",
    x"BF7C258E",
    x"BF7C26A4",
    x"BF7C27B9",
    x"BF7C28CF",
    x"BF7C29E5",
    x"BF7C2AFA",
    x"BF7C2C0F",
    x"BF7C2D24",
    x"BF7C2E39",
    x"BF7C2F4E",
    x"BF7C3062",
    x"BF7C3177",
    x"BF7C328B",
    x"BF7C339F",
    x"BF7C34B3",
    x"BF7C35C7",
    x"BF7C36DB",
    x"BF7C37EE",
    x"BF7C3902",
    x"BF7C3A15",
    x"BF7C3B28",
    x"BF7C3C3B",
    x"BF7C3D4E",
    x"BF7C3E60",
    x"BF7C3F73",
    x"BF7C4085",
    x"BF7C4197",
    x"BF7C42A9",
    x"BF7C43BB",
    x"BF7C44CD",
    x"BF7C45DE",
    x"BF7C46F0",
    x"BF7C4801",
    x"BF7C4912",
    x"BF7C4A23",
    x"BF7C4B34",
    x"BF7C4C44",
    x"BF7C4D55",
    x"BF7C4E65",
    x"BF7C4F75",
    x"BF7C5085",
    x"BF7C5195",
    x"BF7C52A5",
    x"BF7C53B4",
    x"BF7C54C4",
    x"BF7C55D3",
    x"BF7C56E2",
    x"BF7C57F1",
    x"BF7C5900",
    x"BF7C5A0F",
    x"BF7C5B1D",
    x"BF7C5C2C",
    x"BF7C5D3A",
    x"BF7C5E48",
    x"BF7C5F56",
    x"BF7C6063",
    x"BF7C6171",
    x"BF7C627E",
    x"BF7C638C",
    x"BF7C6499",
    x"BF7C65A6",
    x"BF7C66B3",
    x"BF7C67BF",
    x"BF7C68CC",
    x"BF7C69D8",
    x"BF7C6AE5",
    x"BF7C6BF1",
    x"BF7C6CFD",
    x"BF7C6E08",
    x"BF7C6F14",
    x"BF7C701F",
    x"BF7C712B",
    x"BF7C7236",
    x"BF7C7341",
    x"BF7C744C",
    x"BF7C7556",
    x"BF7C7661",
    x"BF7C776B",
    x"BF7C7876",
    x"BF7C7980",
    x"BF7C7A8A",
    x"BF7C7B94",
    x"BF7C7C9D",
    x"BF7C7DA7",
    x"BF7C7EB0",
    x"BF7C7FB9",
    x"BF7C80C2",
    x"BF7C81CB",
    x"BF7C82D4",
    x"BF7C83DC",
    x"BF7C84E5",
    x"BF7C85ED",
    x"BF7C86F5",
    x"BF7C87FD",
    x"BF7C8905",
    x"BF7C8A0D",
    x"BF7C8B14",
    x"BF7C8C1C",
    x"BF7C8D23",
    x"BF7C8E2A",
    x"BF7C8F31",
    x"BF7C9037",
    x"BF7C913E",
    x"BF7C9245",
    x"BF7C934B",
    x"BF7C9451",
    x"BF7C9557",
    x"BF7C965D",
    x"BF7C9762",
    x"BF7C9868",
    x"BF7C996D",
    x"BF7C9A73",
    x"BF7C9B78",
    x"BF7C9C7D",
    x"BF7C9D81",
    x"BF7C9E86",
    x"BF7C9F8A",
    x"BF7CA08F",
    x"BF7CA193",
    x"BF7CA297",
    x"BF7CA39B",
    x"BF7CA49F",
    x"BF7CA5A2",
    x"BF7CA6A6",
    x"BF7CA7A9",
    x"BF7CA8AC",
    x"BF7CA9AF",
    x"BF7CAAB2",
    x"BF7CABB4",
    x"BF7CACB7",
    x"BF7CADB9",
    x"BF7CAEBB",
    x"BF7CAFBD",
    x"BF7CB0BF",
    x"BF7CB1C1",
    x"BF7CB2C2",
    x"BF7CB3C4",
    x"BF7CB4C5",
    x"BF7CB5C6",
    x"BF7CB6C7",
    x"BF7CB7C8",
    x"BF7CB8C9",
    x"BF7CB9C9",
    x"BF7CBACA",
    x"BF7CBBCA",
    x"BF7CBCCA",
    x"BF7CBDCA",
    x"BF7CBECA",
    x"BF7CBFC9",
    x"BF7CC0C9",
    x"BF7CC1C8",
    x"BF7CC2C7",
    x"BF7CC3C6",
    x"BF7CC4C5",
    x"BF7CC5C4",
    x"BF7CC6C2",
    x"BF7CC7C0",
    x"BF7CC8BF",
    x"BF7CC9BD",
    x"BF7CCABB",
    x"BF7CCBB8",
    x"BF7CCCB6",
    x"BF7CCDB4",
    x"BF7CCEB1",
    x"BF7CCFAE",
    x"BF7CD0AB",
    x"BF7CD1A8",
    x"BF7CD2A5",
    x"BF7CD3A1",
    x"BF7CD49E",
    x"BF7CD59A",
    x"BF7CD696",
    x"BF7CD792",
    x"BF7CD88E",
    x"BF7CD989",
    x"BF7CDA85",
    x"BF7CDB80",
    x"BF7CDC7B",
    x"BF7CDD76",
    x"BF7CDE71",
    x"BF7CDF6C",
    x"BF7CE066",
    x"BF7CE161",
    x"BF7CE25B",
    x"BF7CE355",
    x"BF7CE44F",
    x"BF7CE549",
    x"BF7CE643",
    x"BF7CE73C",
    x"BF7CE836",
    x"BF7CE92F",
    x"BF7CEA28",
    x"BF7CEB21",
    x"BF7CEC19",
    x"BF7CED12",
    x"BF7CEE0B",
    x"BF7CEF03",
    x"BF7CEFFB",
    x"BF7CF0F3",
    x"BF7CF1EB",
    x"BF7CF2E2",
    x"BF7CF3DA",
    x"BF7CF4D1",
    x"BF7CF5C9",
    x"BF7CF6C0",
    x"BF7CF7B7",
    x"BF7CF8AD",
    x"BF7CF9A4",
    x"BF7CFA9A",
    x"BF7CFB91",
    x"BF7CFC87",
    x"BF7CFD7D",
    x"BF7CFE73",
    x"BF7CFF68",
    x"BF7D005E",
    x"BF7D0153",
    x"BF7D0249",
    x"BF7D033E",
    x"BF7D0433",
    x"BF7D0527",
    x"BF7D061C",
    x"BF7D0710",
    x"BF7D0805",
    x"BF7D08F9",
    x"BF7D09ED",
    x"BF7D0AE1",
    x"BF7D0BD5",
    x"BF7D0CC8",
    x"BF7D0DBC",
    x"BF7D0EAF",
    x"BF7D0FA2",
    x"BF7D1095",
    x"BF7D1188",
    x"BF7D127A",
    x"BF7D136D",
    x"BF7D145F",
    x"BF7D1551",
    x"BF7D1643",
    x"BF7D1735",
    x"BF7D1827",
    x"BF7D1919",
    x"BF7D1A0A",
    x"BF7D1AFB",
    x"BF7D1BEC",
    x"BF7D1CDD",
    x"BF7D1DCE",
    x"BF7D1EBF",
    x"BF7D1FAF",
    x"BF7D20A0",
    x"BF7D2190",
    x"BF7D2280",
    x"BF7D2370",
    x"BF7D2460",
    x"BF7D254F",
    x"BF7D263F",
    x"BF7D272E",
    x"BF7D281D",
    x"BF7D290C",
    x"BF7D29FB",
    x"BF7D2AEA",
    x"BF7D2BD8",
    x"BF7D2CC7",
    x"BF7D2DB5",
    x"BF7D2EA3",
    x"BF7D2F91",
    x"BF7D307F",
    x"BF7D316C",
    x"BF7D325A",
    x"BF7D3347",
    x"BF7D3434",
    x"BF7D3521",
    x"BF7D360E",
    x"BF7D36FB",
    x"BF7D37E7",
    x"BF7D38D4",
    x"BF7D39C0",
    x"BF7D3AAC",
    x"BF7D3B98",
    x"BF7D3C84",
    x"BF7D3D6F",
    x"BF7D3E5B",
    x"BF7D3F46",
    x"BF7D4031",
    x"BF7D411C",
    x"BF7D4207",
    x"BF7D42F2",
    x"BF7D43DC",
    x"BF7D44C7",
    x"BF7D45B1",
    x"BF7D469B",
    x"BF7D4785",
    x"BF7D486F",
    x"BF7D4959",
    x"BF7D4A42",
    x"BF7D4B2C",
    x"BF7D4C15",
    x"BF7D4CFE",
    x"BF7D4DE7",
    x"BF7D4ECF",
    x"BF7D4FB8",
    x"BF7D50A0",
    x"BF7D5189",
    x"BF7D5271",
    x"BF7D5359",
    x"BF7D5441",
    x"BF7D5528",
    x"BF7D5610",
    x"BF7D56F7",
    x"BF7D57DE",
    x"BF7D58C5",
    x"BF7D59AC",
    x"BF7D5A93",
    x"BF7D5B7A",
    x"BF7D5C60",
    x"BF7D5D46",
    x"BF7D5E2D",
    x"BF7D5F13",
    x"BF7D5FF8",
    x"BF7D60DE",
    x"BF7D61C4",
    x"BF7D62A9",
    x"BF7D638E",
    x"BF7D6473",
    x"BF7D6558",
    x"BF7D663D",
    x"BF7D6722",
    x"BF7D6806",
    x"BF7D68EA",
    x"BF7D69CE",
    x"BF7D6AB2",
    x"BF7D6B96",
    x"BF7D6C7A",
    x"BF7D6D5E",
    x"BF7D6E41",
    x"BF7D6F24",
    x"BF7D7007",
    x"BF7D70EA",
    x"BF7D71CD",
    x"BF7D72B0",
    x"BF7D7392",
    x"BF7D7474",
    x"BF7D7557",
    x"BF7D7639",
    x"BF7D771B",
    x"BF7D77FC",
    x"BF7D78DE",
    x"BF7D79BF",
    x"BF7D7AA0",
    x"BF7D7B82",
    x"BF7D7C62",
    x"BF7D7D43",
    x"BF7D7E24",
    x"BF7D7F04",
    x"BF7D7FE5",
    x"BF7D80C5",
    x"BF7D81A5",
    x"BF7D8285",
    x"BF7D8365",
    x"BF7D8444",
    x"BF7D8524",
    x"BF7D8603",
    x"BF7D86E2",
    x"BF7D87C1",
    x"BF7D88A0",
    x"BF7D897E",
    x"BF7D8A5D",
    x"BF7D8B3B",
    x"BF7D8C19",
    x"BF7D8CF8",
    x"BF7D8DD5",
    x"BF7D8EB3",
    x"BF7D8F91",
    x"BF7D906E",
    x"BF7D914B",
    x"BF7D9229",
    x"BF7D9306",
    x"BF7D93E2",
    x"BF7D94BF",
    x"BF7D959C",
    x"BF7D9678",
    x"BF7D9754",
    x"BF7D9830",
    x"BF7D990C",
    x"BF7D99E8",
    x"BF7D9AC4",
    x"BF7D9B9F",
    x"BF7D9C7A",
    x"BF7D9D55",
    x"BF7D9E30",
    x"BF7D9F0B",
    x"BF7D9FE6",
    x"BF7DA0C0",
    x"BF7DA19B",
    x"BF7DA275",
    x"BF7DA34F",
    x"BF7DA429",
    x"BF7DA503",
    x"BF7DA5DC",
    x"BF7DA6B6",
    x"BF7DA78F",
    x"BF7DA868",
    x"BF7DA941",
    x"BF7DAA1A",
    x"BF7DAAF3",
    x"BF7DABCC",
    x"BF7DACA4",
    x"BF7DAD7C",
    x"BF7DAE54",
    x"BF7DAF2C",
    x"BF7DB004",
    x"BF7DB0DC",
    x"BF7DB1B3",
    x"BF7DB28A",
    x"BF7DB362",
    x"BF7DB439",
    x"BF7DB510",
    x"BF7DB5E6",
    x"BF7DB6BD",
    x"BF7DB793",
    x"BF7DB869",
    x"BF7DB940",
    x"BF7DBA15",
    x"BF7DBAEB",
    x"BF7DBBC1",
    x"BF7DBC96",
    x"BF7DBD6C",
    x"BF7DBE41",
    x"BF7DBF16",
    x"BF7DBFEB",
    x"BF7DC0C0",
    x"BF7DC194",
    x"BF7DC269",
    x"BF7DC33D",
    x"BF7DC411",
    x"BF7DC4E5",
    x"BF7DC5B9",
    x"BF7DC68C",
    x"BF7DC760",
    x"BF7DC833",
    x"BF7DC906",
    x"BF7DC9DA",
    x"BF7DCAAC",
    x"BF7DCB7F",
    x"BF7DCC52",
    x"BF7DCD24",
    x"BF7DCDF6",
    x"BF7DCEC9",
    x"BF7DCF9B",
    x"BF7DD06C",
    x"BF7DD13E",
    x"BF7DD210",
    x"BF7DD2E1",
    x"BF7DD3B2",
    x"BF7DD483",
    x"BF7DD554",
    x"BF7DD625",
    x"BF7DD6F5",
    x"BF7DD7C6",
    x"BF7DD896",
    x"BF7DD966",
    x"BF7DDA36",
    x"BF7DDB06",
    x"BF7DDBD6",
    x"BF7DDCA5",
    x"BF7DDD75",
    x"BF7DDE44",
    x"BF7DDF13",
    x"BF7DDFE2",
    x"BF7DE0B1",
    x"BF7DE17F",
    x"BF7DE24E",
    x"BF7DE31C",
    x"BF7DE3EA",
    x"BF7DE4B8",
    x"BF7DE586",
    x"BF7DE654",
    x"BF7DE721",
    x"BF7DE7EF",
    x"BF7DE8BC",
    x"BF7DE989",
    x"BF7DEA56",
    x"BF7DEB23",
    x"BF7DEBEF",
    x"BF7DECBC",
    x"BF7DED88",
    x"BF7DEE54",
    x"BF7DEF20",
    x"BF7DEFEC",
    x"BF7DF0B8",
    x"BF7DF183",
    x"BF7DF24F",
    x"BF7DF31A",
    x"BF7DF3E5",
    x"BF7DF4B0",
    x"BF7DF57B",
    x"BF7DF646",
    x"BF7DF710",
    x"BF7DF7DA",
    x"BF7DF8A5",
    x"BF7DF96F",
    x"BF7DFA38",
    x"BF7DFB02",
    x"BF7DFBCC",
    x"BF7DFC95",
    x"BF7DFD5E",
    x"BF7DFE28",
    x"BF7DFEF0",
    x"BF7DFFB9",
    x"BF7E0082",
    x"BF7E014A",
    x"BF7E0213",
    x"BF7E02DB",
    x"BF7E03A3",
    x"BF7E046B",
    x"BF7E0533",
    x"BF7E05FA",
    x"BF7E06C2",
    x"BF7E0789",
    x"BF7E0850",
    x"BF7E0917",
    x"BF7E09DE",
    x"BF7E0AA4",
    x"BF7E0B6B",
    x"BF7E0C31",
    x"BF7E0CF7",
    x"BF7E0DBD",
    x"BF7E0E83",
    x"BF7E0F49",
    x"BF7E100F",
    x"BF7E10D4",
    x"BF7E1199",
    x"BF7E125F",
    x"BF7E1324",
    x"BF7E13E8",
    x"BF7E14AD",
    x"BF7E1572",
    x"BF7E1636",
    x"BF7E16FA",
    x"BF7E17BE",
    x"BF7E1882",
    x"BF7E1946",
    x"BF7E1A09",
    x"BF7E1ACD",
    x"BF7E1B90",
    x"BF7E1C53",
    x"BF7E1D16",
    x"BF7E1DD9",
    x"BF7E1E9C",
    x"BF7E1F5E",
    x"BF7E2021",
    x"BF7E20E3",
    x"BF7E21A5",
    x"BF7E2267",
    x"BF7E2329",
    x"BF7E23EA",
    x"BF7E24AC",
    x"BF7E256D",
    x"BF7E262E",
    x"BF7E26EF",
    x"BF7E27B0",
    x"BF7E2871",
    x"BF7E2931",
    x"BF7E29F2",
    x"BF7E2AB2",
    x"BF7E2B72",
    x"BF7E2C32",
    x"BF7E2CF2",
    x"BF7E2DB1",
    x"BF7E2E71",
    x"BF7E2F30",
    x"BF7E2FEF",
    x"BF7E30AE",
    x"BF7E316D",
    x"BF7E322C",
    x"BF7E32EA",
    x"BF7E33A9",
    x"BF7E3467",
    x"BF7E3525",
    x"BF7E35E3",
    x"BF7E36A1",
    x"BF7E375E",
    x"BF7E381C",
    x"BF7E38D9",
    x"BF7E3996",
    x"BF7E3A53",
    x"BF7E3B10",
    x"BF7E3BCD",
    x"BF7E3C89",
    x"BF7E3D46",
    x"BF7E3E02",
    x"BF7E3EBE",
    x"BF7E3F7A",
    x"BF7E4036",
    x"BF7E40F1",
    x"BF7E41AD",
    x"BF7E4268",
    x"BF7E4323",
    x"BF7E43DE",
    x"BF7E4499",
    x"BF7E4554",
    x"BF7E460F",
    x"BF7E46C9",
    x"BF7E4783",
    x"BF7E483D",
    x"BF7E48F7",
    x"BF7E49B1",
    x"BF7E4A6B",
    x"BF7E4B24",
    x"BF7E4BDE",
    x"BF7E4C97",
    x"BF7E4D50",
    x"BF7E4E09",
    x"BF7E4EC1",
    x"BF7E4F7A",
    x"BF7E5032",
    x"BF7E50EB",
    x"BF7E51A3",
    x"BF7E525B",
    x"BF7E5312",
    x"BF7E53CA",
    x"BF7E5482",
    x"BF7E5539",
    x"BF7E55F0",
    x"BF7E56A7",
    x"BF7E575E",
    x"BF7E5815",
    x"BF7E58CB",
    x"BF7E5982",
    x"BF7E5A38",
    x"BF7E5AEE",
    x"BF7E5BA4",
    x"BF7E5C5A",
    x"BF7E5D10",
    x"BF7E5DC5",
    x"BF7E5E7B",
    x"BF7E5F30",
    x"BF7E5FE5",
    x"BF7E609A",
    x"BF7E614E",
    x"BF7E6203",
    x"BF7E62B7",
    x"BF7E636C",
    x"BF7E6420",
    x"BF7E64D4",
    x"BF7E6588",
    x"BF7E663B",
    x"BF7E66EF",
    x"BF7E67A2",
    x"BF7E6855",
    x"BF7E6908",
    x"BF7E69BB",
    x"BF7E6A6E",
    x"BF7E6B21",
    x"BF7E6BD3",
    x"BF7E6C85",
    x"BF7E6D38",
    x"BF7E6DEA",
    x"BF7E6E9B",
    x"BF7E6F4D",
    x"BF7E6FFF",
    x"BF7E70B0",
    x"BF7E7161",
    x"BF7E7212",
    x"BF7E72C3",
    x"BF7E7374",
    x"BF7E7424",
    x"BF7E74D5",
    x"BF7E7585",
    x"BF7E7635",
    x"BF7E76E5",
    x"BF7E7795",
    x"BF7E7845",
    x"BF7E78F4",
    x"BF7E79A4",
    x"BF7E7A53",
    x"BF7E7B02",
    x"BF7E7BB1",
    x"BF7E7C60",
    x"BF7E7D0E",
    x"BF7E7DBD",
    x"BF7E7E6B",
    x"BF7E7F19",
    x"BF7E7FC7",
    x"BF7E8075",
    x"BF7E8123",
    x"BF7E81D0",
    x"BF7E827E",
    x"BF7E832B",
    x"BF7E83D8",
    x"BF7E8485",
    x"BF7E8532",
    x"BF7E85DE",
    x"BF7E868B",
    x"BF7E8737",
    x"BF7E87E3",
    x"BF7E888F",
    x"BF7E893B",
    x"BF7E89E7",
    x"BF7E8A92",
    x"BF7E8B3E",
    x"BF7E8BE9",
    x"BF7E8C94",
    x"BF7E8D3F",
    x"BF7E8DEA",
    x"BF7E8E94",
    x"BF7E8F3F",
    x"BF7E8FE9",
    x"BF7E9093",
    x"BF7E913D",
    x"BF7E91E7",
    x"BF7E9291",
    x"BF7E933A",
    x"BF7E93E4",
    x"BF7E948D",
    x"BF7E9536",
    x"BF7E95DF",
    x"BF7E9688",
    x"BF7E9731",
    x"BF7E97D9",
    x"BF7E9881",
    x"BF7E9929",
    x"BF7E99D2",
    x"BF7E9A79",
    x"BF7E9B21",
    x"BF7E9BC9",
    x"BF7E9C70",
    x"BF7E9D17",
    x"BF7E9DBE",
    x"BF7E9E65",
    x"BF7E9F0C",
    x"BF7E9FB3",
    x"BF7EA059",
    x"BF7EA100",
    x"BF7EA1A6",
    x"BF7EA24C",
    x"BF7EA2F2",
    x"BF7EA397",
    x"BF7EA43D",
    x"BF7EA4E2",
    x"BF7EA588",
    x"BF7EA62D",
    x"BF7EA6D2",
    x"BF7EA776",
    x"BF7EA81B",
    x"BF7EA8C0",
    x"BF7EA964",
    x"BF7EAA08",
    x"BF7EAAAC",
    x"BF7EAB50",
    x"BF7EABF4",
    x"BF7EAC97",
    x"BF7EAD3B",
    x"BF7EADDE",
    x"BF7EAE81",
    x"BF7EAF24",
    x"BF7EAFC7",
    x"BF7EB069",
    x"BF7EB10C",
    x"BF7EB1AE",
    x"BF7EB250",
    x"BF7EB2F2",
    x"BF7EB394",
    x"BF7EB436",
    x"BF7EB4D8",
    x"BF7EB579",
    x"BF7EB61A",
    x"BF7EB6BB",
    x"BF7EB75C",
    x"BF7EB7FD",
    x"BF7EB89E",
    x"BF7EB93E",
    x"BF7EB9DF",
    x"BF7EBA7F",
    x"BF7EBB1F",
    x"BF7EBBBF",
    x"BF7EBC5F",
    x"BF7EBCFE",
    x"BF7EBD9E",
    x"BF7EBE3D",
    x"BF7EBEDC",
    x"BF7EBF7B",
    x"BF7EC01A",
    x"BF7EC0B8",
    x"BF7EC157",
    x"BF7EC1F5",
    x"BF7EC293",
    x"BF7EC331",
    x"BF7EC3CF",
    x"BF7EC46D",
    x"BF7EC50B",
    x"BF7EC5A8",
    x"BF7EC645",
    x"BF7EC6E3",
    x"BF7EC780",
    x"BF7EC81C",
    x"BF7EC8B9",
    x"BF7EC955",
    x"BF7EC9F2",
    x"BF7ECA8E",
    x"BF7ECB2A",
    x"BF7ECBC6",
    x"BF7ECC62",
    x"BF7ECCFD",
    x"BF7ECD99",
    x"BF7ECE34",
    x"BF7ECECF",
    x"BF7ECF6A",
    x"BF7ED005",
    x"BF7ED0A0",
    x"BF7ED13A",
    x"BF7ED1D4",
    x"BF7ED26F",
    x"BF7ED309",
    x"BF7ED3A3",
    x"BF7ED43C",
    x"BF7ED4D6",
    x"BF7ED56F",
    x"BF7ED609",
    x"BF7ED6A2",
    x"BF7ED73B",
    x"BF7ED7D4",
    x"BF7ED86C",
    x"BF7ED905",
    x"BF7ED99D",
    x"BF7EDA35",
    x"BF7EDACD",
    x"BF7EDB65",
    x"BF7EDBFD",
    x"BF7EDC95",
    x"BF7EDD2C",
    x"BF7EDDC3",
    x"BF7EDE5B",
    x"BF7EDEF2",
    x"BF7EDF88",
    x"BF7EE01F",
    x"BF7EE0B6",
    x"BF7EE14C",
    x"BF7EE1E2",
    x"BF7EE278",
    x"BF7EE30E",
    x"BF7EE3A4",
    x"BF7EE43A",
    x"BF7EE4CF",
    x"BF7EE564",
    x"BF7EE5F9",
    x"BF7EE68E",
    x"BF7EE723",
    x"BF7EE7B8",
    x"BF7EE84C",
    x"BF7EE8E1",
    x"BF7EE975",
    x"BF7EEA09",
    x"BF7EEA9D",
    x"BF7EEB31",
    x"BF7EEBC4",
    x"BF7EEC58",
    x"BF7EECEB",
    x"BF7EED7E",
    x"BF7EEE11",
    x"BF7EEEA4",
    x"BF7EEF37",
    x"BF7EEFC9",
    x"BF7EF05C",
    x"BF7EF0EE",
    x"BF7EF180",
    x"BF7EF212",
    x"BF7EF2A4",
    x"BF7EF335",
    x"BF7EF3C7",
    x"BF7EF458",
    x"BF7EF4E9",
    x"BF7EF57A",
    x"BF7EF60B",
    x"BF7EF69C",
    x"BF7EF72C",
    x"BF7EF7BD",
    x"BF7EF84D",
    x"BF7EF8DD",
    x"BF7EF96D",
    x"BF7EF9FD",
    x"BF7EFA8C",
    x"BF7EFB1C",
    x"BF7EFBAB",
    x"BF7EFC3A",
    x"BF7EFCC9",
    x"BF7EFD58",
    x"BF7EFDE7",
    x"BF7EFE75",
    x"BF7EFF04",
    x"BF7EFF92",
    x"BF7F0020",
    x"BF7F00AE",
    x"BF7F013C",
    x"BF7F01C9",
    x"BF7F0257",
    x"BF7F02E4",
    x"BF7F0371",
    x"BF7F03FE",
    x"BF7F048B",
    x"BF7F0518",
    x"BF7F05A4",
    x"BF7F0631",
    x"BF7F06BD",
    x"BF7F0749",
    x"BF7F07D5",
    x"BF7F0861",
    x"BF7F08EC",
    x"BF7F0978",
    x"BF7F0A03",
    x"BF7F0A8E",
    x"BF7F0B19",
    x"BF7F0BA4",
    x"BF7F0C2F",
    x"BF7F0CB9",
    x"BF7F0D44",
    x"BF7F0DCE",
    x"BF7F0E58",
    x"BF7F0EE2",
    x"BF7F0F6C",
    x"BF7F0FF5",
    x"BF7F107F",
    x"BF7F1108",
    x"BF7F1191",
    x"BF7F121A",
    x"BF7F12A3",
    x"BF7F132C",
    x"BF7F13B4",
    x"BF7F143D",
    x"BF7F14C5",
    x"BF7F154D",
    x"BF7F15D5",
    x"BF7F165D",
    x"BF7F16E4",
    x"BF7F176C",
    x"BF7F17F3",
    x"BF7F187A",
    x"BF7F1901",
    x"BF7F1988",
    x"BF7F1A0F",
    x"BF7F1A95",
    x"BF7F1B1C",
    x"BF7F1BA2",
    x"BF7F1C28",
    x"BF7F1CAE",
    x"BF7F1D34",
    x"BF7F1DB9",
    x"BF7F1E3F",
    x"BF7F1EC4",
    x"BF7F1F49",
    x"BF7F1FCE",
    x"BF7F2053",
    x"BF7F20D8",
    x"BF7F215C",
    x"BF7F21E1",
    x"BF7F2265",
    x"BF7F22E9",
    x"BF7F236D",
    x"BF7F23F1",
    x"BF7F2475",
    x"BF7F24F8",
    x"BF7F257B",
    x"BF7F25FF",
    x"BF7F2682",
    x"BF7F2704",
    x"BF7F2787",
    x"BF7F280A",
    x"BF7F288C",
    x"BF7F290E",
    x"BF7F2990",
    x"BF7F2A12",
    x"BF7F2A94",
    x"BF7F2B16",
    x"BF7F2B97",
    x"BF7F2C19",
    x"BF7F2C9A",
    x"BF7F2D1B",
    x"BF7F2D9C",
    x"BF7F2E1C",
    x"BF7F2E9D",
    x"BF7F2F1D",
    x"BF7F2F9D",
    x"BF7F301E",
    x"BF7F309E",
    x"BF7F311D",
    x"BF7F319D",
    x"BF7F321C",
    x"BF7F329C",
    x"BF7F331B",
    x"BF7F339A",
    x"BF7F3419",
    x"BF7F3497",
    x"BF7F3516",
    x"BF7F3594",
    x"BF7F3613",
    x"BF7F3691",
    x"BF7F370F",
    x"BF7F378C",
    x"BF7F380A",
    x"BF7F3888",
    x"BF7F3905",
    x"BF7F3982",
    x"BF7F39FF",
    x"BF7F3A7C",
    x"BF7F3AF9",
    x"BF7F3B75",
    x"BF7F3BF2",
    x"BF7F3C6E",
    x"BF7F3CEA",
    x"BF7F3D66",
    x"BF7F3DE2",
    x"BF7F3E5D",
    x"BF7F3ED9",
    x"BF7F3F54",
    x"BF7F3FCF",
    x"BF7F404A",
    x"BF7F40C5",
    x"BF7F4140",
    x"BF7F41BA",
    x"BF7F4235",
    x"BF7F42AF",
    x"BF7F4329",
    x"BF7F43A3",
    x"BF7F441D",
    x"BF7F4497",
    x"BF7F4510",
    x"BF7F4589",
    x"BF7F4603",
    x"BF7F467C",
    x"BF7F46F4",
    x"BF7F476D",
    x"BF7F47E6",
    x"BF7F485E",
    x"BF7F48D6",
    x"BF7F494E",
    x"BF7F49C6",
    x"BF7F4A3E",
    x"BF7F4AB6",
    x"BF7F4B2D",
    x"BF7F4BA5",
    x"BF7F4C1C",
    x"BF7F4C93",
    x"BF7F4D0A",
    x"BF7F4D80",
    x"BF7F4DF7",
    x"BF7F4E6D",
    x"BF7F4EE4",
    x"BF7F4F5A",
    x"BF7F4FD0",
    x"BF7F5045",
    x"BF7F50BB",
    x"BF7F5131",
    x"BF7F51A6",
    x"BF7F521B",
    x"BF7F5290",
    x"BF7F5305",
    x"BF7F537A",
    x"BF7F53EE",
    x"BF7F5463",
    x"BF7F54D7",
    x"BF7F554B",
    x"BF7F55BF",
    x"BF7F5633",
    x"BF7F56A6",
    x"BF7F571A",
    x"BF7F578D",
    x"BF7F5800",
    x"BF7F5873",
    x"BF7F58E6",
    x"BF7F5959",
    x"BF7F59CC",
    x"BF7F5A3E",
    x"BF7F5AB0",
    x"BF7F5B22",
    x"BF7F5B94",
    x"BF7F5C06",
    x"BF7F5C78",
    x"BF7F5CE9",
    x"BF7F5D5A",
    x"BF7F5DCC",
    x"BF7F5E3D",
    x"BF7F5EAE",
    x"BF7F5F1E",
    x"BF7F5F8F",
    x"BF7F5FFF",
    x"BF7F606F",
    x"BF7F60E0",
    x"BF7F6150",
    x"BF7F61BF",
    x"BF7F622F",
    x"BF7F629E",
    x"BF7F630E",
    x"BF7F637D",
    x"BF7F63EC",
    x"BF7F645B",
    x"BF7F64CA",
    x"BF7F6538",
    x"BF7F65A7",
    x"BF7F6615",
    x"BF7F6683",
    x"BF7F66F1",
    x"BF7F675F",
    x"BF7F67CC",
    x"BF7F683A",
    x"BF7F68A7",
    x"BF7F6914",
    x"BF7F6981",
    x"BF7F69EE",
    x"BF7F6A5B",
    x"BF7F6AC7",
    x"BF7F6B34",
    x"BF7F6BA0",
    x"BF7F6C0C",
    x"BF7F6C78",
    x"BF7F6CE4",
    x"BF7F6D50",
    x"BF7F6DBB",
    x"BF7F6E26",
    x"BF7F6E92",
    x"BF7F6EFD",
    x"BF7F6F67",
    x"BF7F6FD2",
    x"BF7F703D",
    x"BF7F70A7",
    x"BF7F7111",
    x"BF7F717B",
    x"BF7F71E5",
    x"BF7F724F",
    x"BF7F72B9",
    x"BF7F7322",
    x"BF7F738C",
    x"BF7F73F5",
    x"BF7F745E",
    x"BF7F74C7",
    x"BF7F752F",
    x"BF7F7598",
    x"BF7F7600",
    x"BF7F7669",
    x"BF7F76D1",
    x"BF7F7739",
    x"BF7F77A0",
    x"BF7F7808",
    x"BF7F7870",
    x"BF7F78D7",
    x"BF7F793E",
    x"BF7F79A5",
    x"BF7F7A0C",
    x"BF7F7A73",
    x"BF7F7AD9",
    x"BF7F7B40",
    x"BF7F7BA6",
    x"BF7F7C0C",
    x"BF7F7C72",
    x"BF7F7CD8",
    x"BF7F7D3D",
    x"BF7F7DA3",
    x"BF7F7E08",
    x"BF7F7E6D",
    x"BF7F7ED2",
    x"BF7F7F37",
    x"BF7F7F9C",
    x"BF7F8000",
    x"BF7F8065",
    x"BF7F80C9",
    x"BF7F812D",
    x"BF7F8191",
    x"BF7F81F5",
    x"BF7F8259",
    x"BF7F82BC",
    x"BF7F831F",
    x"BF7F8383",
    x"BF7F83E6",
    x"BF7F8448",
    x"BF7F84AB",
    x"BF7F850E",
    x"BF7F8570",
    x"BF7F85D2",
    x"BF7F8634",
    x"BF7F8696",
    x"BF7F86F8",
    x"BF7F875A",
    x"BF7F87BB",
    x"BF7F881D",
    x"BF7F887E",
    x"BF7F88DF",
    x"BF7F8940",
    x"BF7F89A0",
    x"BF7F8A01",
    x"BF7F8A61",
    x"BF7F8AC2",
    x"BF7F8B22",
    x"BF7F8B82",
    x"BF7F8BE1",
    x"BF7F8C41",
    x"BF7F8CA1",
    x"BF7F8D00",
    x"BF7F8D5F",
    x"BF7F8DBE",
    x"BF7F8E1D",
    x"BF7F8E7C",
    x"BF7F8EDA",
    x"BF7F8F39",
    x"BF7F8F97",
    x"BF7F8FF5",
    x"BF7F9053",
    x"BF7F90B1",
    x"BF7F910E",
    x"BF7F916C",
    x"BF7F91C9",
    x"BF7F9226",
    x"BF7F9283",
    x"BF7F92E0",
    x"BF7F933D",
    x"BF7F9399",
    x"BF7F93F6",
    x"BF7F9452",
    x"BF7F94AE",
    x"BF7F950A",
    x"BF7F9566",
    x"BF7F95C1",
    x"BF7F961D",
    x"BF7F9678",
    x"BF7F96D3",
    x"BF7F972E",
    x"BF7F9789",
    x"BF7F97E4",
    x"BF7F983F",
    x"BF7F9899",
    x"BF7F98F3",
    x"BF7F994D",
    x"BF7F99A7",
    x"BF7F9A01",
    x"BF7F9A5B",
    x"BF7F9AB4",
    x"BF7F9B0D",
    x"BF7F9B67",
    x"BF7F9BC0",
    x"BF7F9C18",
    x"BF7F9C71",
    x"BF7F9CCA",
    x"BF7F9D22",
    x"BF7F9D7A",
    x"BF7F9DD2",
    x"BF7F9E2A",
    x"BF7F9E82",
    x"BF7F9EDA",
    x"BF7F9F31",
    x"BF7F9F89",
    x"BF7F9FE0",
    x"BF7FA037",
    x"BF7FA08E",
    x"BF7FA0E4",
    x"BF7FA13B",
    x"BF7FA191",
    x"BF7FA1E8",
    x"BF7FA23E",
    x"BF7FA294",
    x"BF7FA2E9",
    x"BF7FA33F",
    x"BF7FA394",
    x"BF7FA3EA",
    x"BF7FA43F",
    x"BF7FA494",
    x"BF7FA4E9",
    x"BF7FA53D",
    x"BF7FA592",
    x"BF7FA5E6",
    x"BF7FA63B",
    x"BF7FA68F",
    x"BF7FA6E3",
    x"BF7FA736",
    x"BF7FA78A",
    x"BF7FA7DE",
    x"BF7FA831",
    x"BF7FA884",
    x"BF7FA8D7",
    x"BF7FA92A",
    x"BF7FA97D",
    x"BF7FA9CF",
    x"BF7FAA21",
    x"BF7FAA74",
    x"BF7FAAC6",
    x"BF7FAB18",
    x"BF7FAB6A",
    x"BF7FABBB",
    x"BF7FAC0D",
    x"BF7FAC5E",
    x"BF7FACAF",
    x"BF7FAD00",
    x"BF7FAD51",
    x"BF7FADA2",
    x"BF7FADF2",
    x"BF7FAE43",
    x"BF7FAE93",
    x"BF7FAEE3",
    x"BF7FAF33",
    x"BF7FAF83",
    x"BF7FAFD2",
    x"BF7FB022",
    x"BF7FB071",
    x"BF7FB0C0",
    x"BF7FB10F",
    x"BF7FB15E",
    x"BF7FB1AD",
    x"BF7FB1FB",
    x"BF7FB24A",
    x"BF7FB298",
    x"BF7FB2E6",
    x"BF7FB334",
    x"BF7FB382",
    x"BF7FB3CF",
    x"BF7FB41D",
    x"BF7FB46A",
    x"BF7FB4B7",
    x"BF7FB504",
    x"BF7FB551",
    x"BF7FB59E",
    x"BF7FB5EA",
    x"BF7FB637",
    x"BF7FB683",
    x"BF7FB6CF",
    x"BF7FB71B",
    x"BF7FB767",
    x"BF7FB7B2",
    x"BF7FB7FE",
    x"BF7FB849",
    x"BF7FB894",
    x"BF7FB8DF",
    x"BF7FB92A",
    x"BF7FB975",
    x"BF7FB9BF",
    x"BF7FBA0A",
    x"BF7FBA54",
    x"BF7FBA9E",
    x"BF7FBAE8",
    x"BF7FBB32",
    x"BF7FBB7B",
    x"BF7FBBC5",
    x"BF7FBC0E",
    x"BF7FBC57",
    x"BF7FBCA0",
    x"BF7FBCE9",
    x"BF7FBD32",
    x"BF7FBD7A",
    x"BF7FBDC2",
    x"BF7FBE0B",
    x"BF7FBE53",
    x"BF7FBE9B",
    x"BF7FBEE2",
    x"BF7FBF2A",
    x"BF7FBF72",
    x"BF7FBFB9",
    x"BF7FC000",
    x"BF7FC047",
    x"BF7FC08E",
    x"BF7FC0D4",
    x"BF7FC11B",
    x"BF7FC161",
    x"BF7FC1A8",
    x"BF7FC1EE",
    x"BF7FC234",
    x"BF7FC279",
    x"BF7FC2BF",
    x"BF7FC304",
    x"BF7FC34A",
    x"BF7FC38F",
    x"BF7FC3D4",
    x"BF7FC419",
    x"BF7FC45D",
    x"BF7FC4A2",
    x"BF7FC4E6",
    x"BF7FC52A",
    x"BF7FC56F",
    x"BF7FC5B2",
    x"BF7FC5F6",
    x"BF7FC63A",
    x"BF7FC67D",
    x"BF7FC6C1",
    x"BF7FC704",
    x"BF7FC747",
    x"BF7FC789",
    x"BF7FC7CC",
    x"BF7FC80F",
    x"BF7FC851",
    x"BF7FC893",
    x"BF7FC8D5",
    x"BF7FC917",
    x"BF7FC959",
    x"BF7FC99B",
    x"BF7FC9DC",
    x"BF7FCA1D",
    x"BF7FCA5E",
    x"BF7FCA9F",
    x"BF7FCAE0",
    x"BF7FCB21",
    x"BF7FCB61",
    x"BF7FCBA2",
    x"BF7FCBE2",
    x"BF7FCC22",
    x"BF7FCC62",
    x"BF7FCCA2",
    x"BF7FCCE1",
    x"BF7FCD21",
    x"BF7FCD60",
    x"BF7FCD9F",
    x"BF7FCDDE",
    x"BF7FCE1D",
    x"BF7FCE5C",
    x"BF7FCE9A",
    x"BF7FCED9",
    x"BF7FCF17",
    x"BF7FCF55",
    x"BF7FCF93",
    x"BF7FCFD1",
    x"BF7FD00E",
    x"BF7FD04C",
    x"BF7FD089",
    x"BF7FD0C6",
    x"BF7FD103",
    x"BF7FD140",
    x"BF7FD17C",
    x"BF7FD1B9",
    x"BF7FD1F5",
    x"BF7FD232",
    x"BF7FD26E",
    x"BF7FD2A9",
    x"BF7FD2E5",
    x"BF7FD321",
    x"BF7FD35C",
    x"BF7FD397",
    x"BF7FD3D3",
    x"BF7FD40E",
    x"BF7FD448",
    x"BF7FD483",
    x"BF7FD4BE",
    x"BF7FD4F8",
    x"BF7FD532",
    x"BF7FD56C",
    x"BF7FD5A6",
    x"BF7FD5E0",
    x"BF7FD619",
    x"BF7FD653",
    x"BF7FD68C",
    x"BF7FD6C5",
    x"BF7FD6FE",
    x"BF7FD737",
    x"BF7FD770",
    x"BF7FD7A8",
    x"BF7FD7E1",
    x"BF7FD819",
    x"BF7FD851",
    x"BF7FD889",
    x"BF7FD8C0",
    x"BF7FD8F8",
    x"BF7FD92F",
    x"BF7FD967",
    x"BF7FD99E",
    x"BF7FD9D5",
    x"BF7FDA0C",
    x"BF7FDA42",
    x"BF7FDA79",
    x"BF7FDAAF",
    x"BF7FDAE5",
    x"BF7FDB1B",
    x"BF7FDB51",
    x"BF7FDB87",
    x"BF7FDBBD",
    x"BF7FDBF2",
    x"BF7FDC27",
    x"BF7FDC5C",
    x"BF7FDC91",
    x"BF7FDCC6",
    x"BF7FDCFB",
    x"BF7FDD2F",
    x"BF7FDD64",
    x"BF7FDD98",
    x"BF7FDDCC",
    x"BF7FDE00",
    x"BF7FDE33",
    x"BF7FDE67",
    x"BF7FDE9A",
    x"BF7FDECE",
    x"BF7FDF01",
    x"BF7FDF34",
    x"BF7FDF67",
    x"BF7FDF99",
    x"BF7FDFCC",
    x"BF7FDFFE",
    x"BF7FE030",
    x"BF7FE062",
    x"BF7FE094",
    x"BF7FE0C6",
    x"BF7FE0F8",
    x"BF7FE129",
    x"BF7FE15A",
    x"BF7FE18B",
    x"BF7FE1BC",
    x"BF7FE1ED",
    x"BF7FE21E",
    x"BF7FE24E",
    x"BF7FE27F",
    x"BF7FE2AF",
    x"BF7FE2DF",
    x"BF7FE30F",
    x"BF7FE33E",
    x"BF7FE36E",
    x"BF7FE39D",
    x"BF7FE3CD",
    x"BF7FE3FC",
    x"BF7FE42B",
    x"BF7FE459",
    x"BF7FE488",
    x"BF7FE4B7",
    x"BF7FE4E5",
    x"BF7FE513",
    x"BF7FE541",
    x"BF7FE56F",
    x"BF7FE59D",
    x"BF7FE5CA",
    x"BF7FE5F8",
    x"BF7FE625",
    x"BF7FE652",
    x"BF7FE67F",
    x"BF7FE6AC",
    x"BF7FE6D8",
    x"BF7FE705",
    x"BF7FE731",
    x"BF7FE75D",
    x"BF7FE789",
    x"BF7FE7B5",
    x"BF7FE7E1",
    x"BF7FE80D",
    x"BF7FE838",
    x"BF7FE863",
    x"BF7FE88E",
    x"BF7FE8B9",
    x"BF7FE8E4",
    x"BF7FE90F",
    x"BF7FE939",
    x"BF7FE964",
    x"BF7FE98E",
    x"BF7FE9B8",
    x"BF7FE9E2",
    x"BF7FEA0B",
    x"BF7FEA35",
    x"BF7FEA5E",
    x"BF7FEA87",
    x"BF7FEAB1",
    x"BF7FEADA",
    x"BF7FEB02",
    x"BF7FEB2B",
    x"BF7FEB53",
    x"BF7FEB7C",
    x"BF7FEBA4",
    x"BF7FEBCC",
    x"BF7FEBF4",
    x"BF7FEC1B",
    x"BF7FEC43",
    x"BF7FEC6A",
    x"BF7FEC92",
    x"BF7FECB9",
    x"BF7FECE0",
    x"BF7FED06",
    x"BF7FED2D",
    x"BF7FED54",
    x"BF7FED7A",
    x"BF7FEDA0",
    x"BF7FEDC6",
    x"BF7FEDEC",
    x"BF7FEE12",
    x"BF7FEE37",
    x"BF7FEE5D",
    x"BF7FEE82",
    x"BF7FEEA7",
    x"BF7FEECC",
    x"BF7FEEF1",
    x"BF7FEF15",
    x"BF7FEF3A",
    x"BF7FEF5E",
    x"BF7FEF82",
    x"BF7FEFA6",
    x"BF7FEFCA",
    x"BF7FEFEE",
    x"BF7FF011",
    x"BF7FF035",
    x"BF7FF058",
    x"BF7FF07B",
    x"BF7FF09E",
    x"BF7FF0C1",
    x"BF7FF0E3",
    x"BF7FF106",
    x"BF7FF128",
    x"BF7FF14A",
    x"BF7FF16C",
    x"BF7FF18E",
    x"BF7FF1B0",
    x"BF7FF1D1",
    x"BF7FF1F3",
    x"BF7FF214",
    x"BF7FF235",
    x"BF7FF256",
    x"BF7FF277",
    x"BF7FF297",
    x"BF7FF2B8",
    x"BF7FF2D8",
    x"BF7FF2F8",
    x"BF7FF318",
    x"BF7FF338",
    x"BF7FF358",
    x"BF7FF377",
    x"BF7FF397",
    x"BF7FF3B6",
    x"BF7FF3D5",
    x"BF7FF3F4",
    x"BF7FF413",
    x"BF7FF431",
    x"BF7FF450",
    x"BF7FF46E",
    x"BF7FF48C",
    x"BF7FF4AA",
    x"BF7FF4C8",
    x"BF7FF4E6",
    x"BF7FF503",
    x"BF7FF521",
    x"BF7FF53E",
    x"BF7FF55B",
    x"BF7FF578",
    x"BF7FF595",
    x"BF7FF5B1",
    x"BF7FF5CE",
    x"BF7FF5EA",
    x"BF7FF606",
    x"BF7FF622",
    x"BF7FF63E",
    x"BF7FF659",
    x"BF7FF675",
    x"BF7FF690",
    x"BF7FF6AC",
    x"BF7FF6C7",
    x"BF7FF6E2",
    x"BF7FF6FC",
    x"BF7FF717",
    x"BF7FF731",
    x"BF7FF74C",
    x"BF7FF766",
    x"BF7FF780",
    x"BF7FF79A",
    x"BF7FF7B3",
    x"BF7FF7CD",
    x"BF7FF7E6",
    x"BF7FF7FF",
    x"BF7FF818",
    x"BF7FF831",
    x"BF7FF84A",
    x"BF7FF863",
    x"BF7FF87B",
    x"BF7FF893",
    x"BF7FF8AC",
    x"BF7FF8C4",
    x"BF7FF8DB",
    x"BF7FF8F3",
    x"BF7FF90B",
    x"BF7FF922",
    x"BF7FF939",
    x"BF7FF950",
    x"BF7FF967",
    x"BF7FF97E",
    x"BF7FF994",
    x"BF7FF9AB",
    x"BF7FF9C1",
    x"BF7FF9D7",
    x"BF7FF9ED",
    x"BF7FFA03",
    x"BF7FFA19",
    x"BF7FFA2E",
    x"BF7FFA44",
    x"BF7FFA59",
    x"BF7FFA6E",
    x"BF7FFA83",
    x"BF7FFA97",
    x"BF7FFAAC",
    x"BF7FFAC1",
    x"BF7FFAD5",
    x"BF7FFAE9",
    x"BF7FFAFD",
    x"BF7FFB11",
    x"BF7FFB24",
    x"BF7FFB38",
    x"BF7FFB4B",
    x"BF7FFB5E",
    x"BF7FFB71",
    x"BF7FFB84",
    x"BF7FFB97",
    x"BF7FFBAA",
    x"BF7FFBBC",
    x"BF7FFBCE",
    x"BF7FFBE1",
    x"BF7FFBF2",
    x"BF7FFC04",
    x"BF7FFC16",
    x"BF7FFC27",
    x"BF7FFC39",
    x"BF7FFC4A",
    x"BF7FFC5B",
    x"BF7FFC6C",
    x"BF7FFC7D",
    x"BF7FFC8D",
    x"BF7FFC9E",
    x"BF7FFCAE",
    x"BF7FFCBE",
    x"BF7FFCCE",
    x"BF7FFCDE",
    x"BF7FFCED",
    x"BF7FFCFD",
    x"BF7FFD0C",
    x"BF7FFD1B",
    x"BF7FFD2B",
    x"BF7FFD39",
    x"BF7FFD48",
    x"BF7FFD57",
    x"BF7FFD65",
    x"BF7FFD73",
    x"BF7FFD81",
    x"BF7FFD8F",
    x"BF7FFD9D",
    x"BF7FFDAB",
    x"BF7FFDB8",
    x"BF7FFDC6",
    x"BF7FFDD3",
    x"BF7FFDE0",
    x"BF7FFDED",
    x"BF7FFDFA",
    x"BF7FFE06",
    x"BF7FFE13",
    x"BF7FFE1F",
    x"BF7FFE2B",
    x"BF7FFE37",
    x"BF7FFE43",
    x"BF7FFE4E",
    x"BF7FFE5A",
    x"BF7FFE65",
    x"BF7FFE70",
    x"BF7FFE7B",
    x"BF7FFE86",
    x"BF7FFE91",
    x"BF7FFE9B",
    x"BF7FFEA6",
    x"BF7FFEB0",
    x"BF7FFEBA",
    x"BF7FFEC4",
    x"BF7FFECE",
    x"BF7FFED8",
    x"BF7FFEE1",
    x"BF7FFEEA",
    x"BF7FFEF4",
    x"BF7FFEFD",
    x"BF7FFF05",
    x"BF7FFF0E",
    x"BF7FFF17",
    x"BF7FFF1F",
    x"BF7FFF27",
    x"BF7FFF30",
    x"BF7FFF37",
    x"BF7FFF3F",
    x"BF7FFF47",
    x"BF7FFF4E",
    x"BF7FFF56",
    x"BF7FFF5D",
    x"BF7FFF64",
    x"BF7FFF6B",
    x"BF7FFF71",
    x"BF7FFF78",
    x"BF7FFF7E",
    x"BF7FFF85",
    x"BF7FFF8B",
    x"BF7FFF91",
    x"BF7FFF96",
    x"BF7FFF9C",
    x"BF7FFFA2",
    x"BF7FFFA7",
    x"BF7FFFAC",
    x"BF7FFFB1",
    x"BF7FFFB6",
    x"BF7FFFBB",
    x"BF7FFFBF",
    x"BF7FFFC4",
    x"BF7FFFC8",
    x"BF7FFFCC",
    x"BF7FFFD0",
    x"BF7FFFD4",
    x"BF7FFFD7",
    x"BF7FFFDB",
    x"BF7FFFDE",
    x"BF7FFFE1",
    x"BF7FFFE4",
    x"BF7FFFE7",
    x"BF7FFFEA",
    x"BF7FFFEC",
    x"BF7FFFEF",
    x"BF7FFFF1",
    x"BF7FFFF3",
    x"BF7FFFF5",
    x"BF7FFFF7",
    x"BF7FFFF8",
    x"BF7FFFFA",
    x"BF7FFFFB",
    x"BF7FFFFC",
    x"BF7FFFFD",
    x"BF7FFFFE",
    x"BF7FFFFF",
    x"BF7FFFFF",
    x"BF800000",
    x"BF800000",
    x"BF800000",
    x"BF800000",
    x"BF800000",
    x"BF7FFFFF",
    x"BF7FFFFF",
    x"BF7FFFFE",
    x"BF7FFFFD",
    x"BF7FFFFC",
    x"BF7FFFFB",
    x"BF7FFFFA",
    x"BF7FFFF8",
    x"BF7FFFF7",
    x"BF7FFFF5",
    x"BF7FFFF3",
    x"BF7FFFF1",
    x"BF7FFFEF",
    x"BF7FFFEC",
    x"BF7FFFEA",
    x"BF7FFFE7",
    x"BF7FFFE4",
    x"BF7FFFE1",
    x"BF7FFFDE",
    x"BF7FFFDB",
    x"BF7FFFD7",
    x"BF7FFFD4",
    x"BF7FFFD0",
    x"BF7FFFCC",
    x"BF7FFFC8",
    x"BF7FFFC4",
    x"BF7FFFBF",
    x"BF7FFFBB",
    x"BF7FFFB6",
    x"BF7FFFB1",
    x"BF7FFFAC",
    x"BF7FFFA7",
    x"BF7FFFA2",
    x"BF7FFF9C",
    x"BF7FFF96",
    x"BF7FFF91",
    x"BF7FFF8B",
    x"BF7FFF85",
    x"BF7FFF7E",
    x"BF7FFF78",
    x"BF7FFF71",
    x"BF7FFF6B",
    x"BF7FFF64",
    x"BF7FFF5D",
    x"BF7FFF56",
    x"BF7FFF4E",
    x"BF7FFF47",
    x"BF7FFF3F",
    x"BF7FFF37",
    x"BF7FFF30",
    x"BF7FFF27",
    x"BF7FFF1F",
    x"BF7FFF17",
    x"BF7FFF0E",
    x"BF7FFF05",
    x"BF7FFEFD",
    x"BF7FFEF4",
    x"BF7FFEEA",
    x"BF7FFEE1",
    x"BF7FFED8",
    x"BF7FFECE",
    x"BF7FFEC4",
    x"BF7FFEBA",
    x"BF7FFEB0",
    x"BF7FFEA6",
    x"BF7FFE9B",
    x"BF7FFE91",
    x"BF7FFE86",
    x"BF7FFE7B",
    x"BF7FFE70",
    x"BF7FFE65",
    x"BF7FFE5A",
    x"BF7FFE4E",
    x"BF7FFE43",
    x"BF7FFE37",
    x"BF7FFE2B",
    x"BF7FFE1F",
    x"BF7FFE13",
    x"BF7FFE06",
    x"BF7FFDFA",
    x"BF7FFDED",
    x"BF7FFDE0",
    x"BF7FFDD3",
    x"BF7FFDC6",
    x"BF7FFDB8",
    x"BF7FFDAB",
    x"BF7FFD9D",
    x"BF7FFD8F",
    x"BF7FFD81",
    x"BF7FFD73",
    x"BF7FFD65",
    x"BF7FFD57",
    x"BF7FFD48",
    x"BF7FFD39",
    x"BF7FFD2B",
    x"BF7FFD1B",
    x"BF7FFD0C",
    x"BF7FFCFD",
    x"BF7FFCED",
    x"BF7FFCDE",
    x"BF7FFCCE",
    x"BF7FFCBE",
    x"BF7FFCAE",
    x"BF7FFC9E",
    x"BF7FFC8D",
    x"BF7FFC7D",
    x"BF7FFC6C",
    x"BF7FFC5B",
    x"BF7FFC4A",
    x"BF7FFC39",
    x"BF7FFC27",
    x"BF7FFC16",
    x"BF7FFC04",
    x"BF7FFBF2",
    x"BF7FFBE1",
    x"BF7FFBCE",
    x"BF7FFBBC",
    x"BF7FFBAA",
    x"BF7FFB97",
    x"BF7FFB84",
    x"BF7FFB71",
    x"BF7FFB5E",
    x"BF7FFB4B",
    x"BF7FFB38",
    x"BF7FFB24",
    x"BF7FFB11",
    x"BF7FFAFD",
    x"BF7FFAE9",
    x"BF7FFAD5",
    x"BF7FFAC1",
    x"BF7FFAAC",
    x"BF7FFA97",
    x"BF7FFA83",
    x"BF7FFA6E",
    x"BF7FFA59",
    x"BF7FFA44",
    x"BF7FFA2E",
    x"BF7FFA19",
    x"BF7FFA03",
    x"BF7FF9ED",
    x"BF7FF9D7",
    x"BF7FF9C1",
    x"BF7FF9AB",
    x"BF7FF994",
    x"BF7FF97E",
    x"BF7FF967",
    x"BF7FF950",
    x"BF7FF939",
    x"BF7FF922",
    x"BF7FF90B",
    x"BF7FF8F3",
    x"BF7FF8DB",
    x"BF7FF8C4",
    x"BF7FF8AC",
    x"BF7FF893",
    x"BF7FF87B",
    x"BF7FF863",
    x"BF7FF84A",
    x"BF7FF831",
    x"BF7FF818",
    x"BF7FF7FF",
    x"BF7FF7E6",
    x"BF7FF7CD",
    x"BF7FF7B3",
    x"BF7FF79A",
    x"BF7FF780",
    x"BF7FF766",
    x"BF7FF74C",
    x"BF7FF731",
    x"BF7FF717",
    x"BF7FF6FC",
    x"BF7FF6E2",
    x"BF7FF6C7",
    x"BF7FF6AC",
    x"BF7FF690",
    x"BF7FF675",
    x"BF7FF659",
    x"BF7FF63E",
    x"BF7FF622",
    x"BF7FF606",
    x"BF7FF5EA",
    x"BF7FF5CE",
    x"BF7FF5B1",
    x"BF7FF595",
    x"BF7FF578",
    x"BF7FF55B",
    x"BF7FF53E",
    x"BF7FF521",
    x"BF7FF503",
    x"BF7FF4E6",
    x"BF7FF4C8",
    x"BF7FF4AA",
    x"BF7FF48C",
    x"BF7FF46E",
    x"BF7FF450",
    x"BF7FF431",
    x"BF7FF413",
    x"BF7FF3F4",
    x"BF7FF3D5",
    x"BF7FF3B6",
    x"BF7FF397",
    x"BF7FF377",
    x"BF7FF358",
    x"BF7FF338",
    x"BF7FF318",
    x"BF7FF2F8",
    x"BF7FF2D8",
    x"BF7FF2B8",
    x"BF7FF297",
    x"BF7FF277",
    x"BF7FF256",
    x"BF7FF235",
    x"BF7FF214",
    x"BF7FF1F3",
    x"BF7FF1D1",
    x"BF7FF1B0",
    x"BF7FF18E",
    x"BF7FF16C",
    x"BF7FF14A",
    x"BF7FF128",
    x"BF7FF106",
    x"BF7FF0E3",
    x"BF7FF0C1",
    x"BF7FF09E",
    x"BF7FF07B",
    x"BF7FF058",
    x"BF7FF035",
    x"BF7FF011",
    x"BF7FEFEE",
    x"BF7FEFCA",
    x"BF7FEFA6",
    x"BF7FEF82",
    x"BF7FEF5E",
    x"BF7FEF3A",
    x"BF7FEF15",
    x"BF7FEEF1",
    x"BF7FEECC",
    x"BF7FEEA7",
    x"BF7FEE82",
    x"BF7FEE5D",
    x"BF7FEE37",
    x"BF7FEE12",
    x"BF7FEDEC",
    x"BF7FEDC6",
    x"BF7FEDA0",
    x"BF7FED7A",
    x"BF7FED54",
    x"BF7FED2D",
    x"BF7FED06",
    x"BF7FECE0",
    x"BF7FECB9",
    x"BF7FEC92",
    x"BF7FEC6A",
    x"BF7FEC43",
    x"BF7FEC1B",
    x"BF7FEBF4",
    x"BF7FEBCC",
    x"BF7FEBA4",
    x"BF7FEB7C",
    x"BF7FEB53",
    x"BF7FEB2B",
    x"BF7FEB02",
    x"BF7FEADA",
    x"BF7FEAB1",
    x"BF7FEA87",
    x"BF7FEA5E",
    x"BF7FEA35",
    x"BF7FEA0B",
    x"BF7FE9E2",
    x"BF7FE9B8",
    x"BF7FE98E",
    x"BF7FE964",
    x"BF7FE939",
    x"BF7FE90F",
    x"BF7FE8E4",
    x"BF7FE8B9",
    x"BF7FE88E",
    x"BF7FE863",
    x"BF7FE838",
    x"BF7FE80D",
    x"BF7FE7E1",
    x"BF7FE7B5",
    x"BF7FE789",
    x"BF7FE75D",
    x"BF7FE731",
    x"BF7FE705",
    x"BF7FE6D8",
    x"BF7FE6AC",
    x"BF7FE67F",
    x"BF7FE652",
    x"BF7FE625",
    x"BF7FE5F8",
    x"BF7FE5CA",
    x"BF7FE59D",
    x"BF7FE56F",
    x"BF7FE541",
    x"BF7FE513",
    x"BF7FE4E5",
    x"BF7FE4B7",
    x"BF7FE488",
    x"BF7FE459",
    x"BF7FE42B",
    x"BF7FE3FC",
    x"BF7FE3CD",
    x"BF7FE39D",
    x"BF7FE36E",
    x"BF7FE33E",
    x"BF7FE30F",
    x"BF7FE2DF",
    x"BF7FE2AF",
    x"BF7FE27F",
    x"BF7FE24E",
    x"BF7FE21E",
    x"BF7FE1ED",
    x"BF7FE1BC",
    x"BF7FE18B",
    x"BF7FE15A",
    x"BF7FE129",
    x"BF7FE0F8",
    x"BF7FE0C6",
    x"BF7FE094",
    x"BF7FE062",
    x"BF7FE030",
    x"BF7FDFFE",
    x"BF7FDFCC",
    x"BF7FDF99",
    x"BF7FDF67",
    x"BF7FDF34",
    x"BF7FDF01",
    x"BF7FDECE",
    x"BF7FDE9A",
    x"BF7FDE67",
    x"BF7FDE33",
    x"BF7FDE00",
    x"BF7FDDCC",
    x"BF7FDD98",
    x"BF7FDD64",
    x"BF7FDD2F",
    x"BF7FDCFB",
    x"BF7FDCC6",
    x"BF7FDC91",
    x"BF7FDC5C",
    x"BF7FDC27",
    x"BF7FDBF2",
    x"BF7FDBBD",
    x"BF7FDB87",
    x"BF7FDB51",
    x"BF7FDB1B",
    x"BF7FDAE5",
    x"BF7FDAAF",
    x"BF7FDA79",
    x"BF7FDA42",
    x"BF7FDA0C",
    x"BF7FD9D5",
    x"BF7FD99E",
    x"BF7FD967",
    x"BF7FD92F",
    x"BF7FD8F8",
    x"BF7FD8C0",
    x"BF7FD889",
    x"BF7FD851",
    x"BF7FD819",
    x"BF7FD7E1",
    x"BF7FD7A8",
    x"BF7FD770",
    x"BF7FD737",
    x"BF7FD6FE",
    x"BF7FD6C5",
    x"BF7FD68C",
    x"BF7FD653",
    x"BF7FD619",
    x"BF7FD5E0",
    x"BF7FD5A6",
    x"BF7FD56C",
    x"BF7FD532",
    x"BF7FD4F8",
    x"BF7FD4BE",
    x"BF7FD483",
    x"BF7FD448",
    x"BF7FD40E",
    x"BF7FD3D3",
    x"BF7FD397",
    x"BF7FD35C",
    x"BF7FD321",
    x"BF7FD2E5",
    x"BF7FD2A9",
    x"BF7FD26E",
    x"BF7FD232",
    x"BF7FD1F5",
    x"BF7FD1B9",
    x"BF7FD17C",
    x"BF7FD140",
    x"BF7FD103",
    x"BF7FD0C6",
    x"BF7FD089",
    x"BF7FD04C",
    x"BF7FD00E",
    x"BF7FCFD1",
    x"BF7FCF93",
    x"BF7FCF55",
    x"BF7FCF17",
    x"BF7FCED9",
    x"BF7FCE9A",
    x"BF7FCE5C",
    x"BF7FCE1D",
    x"BF7FCDDE",
    x"BF7FCD9F",
    x"BF7FCD60",
    x"BF7FCD21",
    x"BF7FCCE1",
    x"BF7FCCA2",
    x"BF7FCC62",
    x"BF7FCC22",
    x"BF7FCBE2",
    x"BF7FCBA2",
    x"BF7FCB61",
    x"BF7FCB21",
    x"BF7FCAE0",
    x"BF7FCA9F",
    x"BF7FCA5E",
    x"BF7FCA1D",
    x"BF7FC9DC",
    x"BF7FC99B",
    x"BF7FC959",
    x"BF7FC917",
    x"BF7FC8D5",
    x"BF7FC893",
    x"BF7FC851",
    x"BF7FC80F",
    x"BF7FC7CC",
    x"BF7FC789",
    x"BF7FC747",
    x"BF7FC704",
    x"BF7FC6C1",
    x"BF7FC67D",
    x"BF7FC63A",
    x"BF7FC5F6",
    x"BF7FC5B2",
    x"BF7FC56F",
    x"BF7FC52A",
    x"BF7FC4E6",
    x"BF7FC4A2",
    x"BF7FC45D",
    x"BF7FC419",
    x"BF7FC3D4",
    x"BF7FC38F",
    x"BF7FC34A",
    x"BF7FC304",
    x"BF7FC2BF",
    x"BF7FC279",
    x"BF7FC234",
    x"BF7FC1EE",
    x"BF7FC1A8",
    x"BF7FC161",
    x"BF7FC11B",
    x"BF7FC0D4",
    x"BF7FC08E",
    x"BF7FC047",
    x"BF7FC000",
    x"BF7FBFB9",
    x"BF7FBF72",
    x"BF7FBF2A",
    x"BF7FBEE2",
    x"BF7FBE9B",
    x"BF7FBE53",
    x"BF7FBE0B",
    x"BF7FBDC2",
    x"BF7FBD7A",
    x"BF7FBD32",
    x"BF7FBCE9",
    x"BF7FBCA0",
    x"BF7FBC57",
    x"BF7FBC0E",
    x"BF7FBBC5",
    x"BF7FBB7B",
    x"BF7FBB32",
    x"BF7FBAE8",
    x"BF7FBA9E",
    x"BF7FBA54",
    x"BF7FBA0A",
    x"BF7FB9BF",
    x"BF7FB975",
    x"BF7FB92A",
    x"BF7FB8DF",
    x"BF7FB894",
    x"BF7FB849",
    x"BF7FB7FE",
    x"BF7FB7B2",
    x"BF7FB767",
    x"BF7FB71B",
    x"BF7FB6CF",
    x"BF7FB683",
    x"BF7FB637",
    x"BF7FB5EA",
    x"BF7FB59E",
    x"BF7FB551",
    x"BF7FB504",
    x"BF7FB4B7",
    x"BF7FB46A",
    x"BF7FB41D",
    x"BF7FB3CF",
    x"BF7FB382",
    x"BF7FB334",
    x"BF7FB2E6",
    x"BF7FB298",
    x"BF7FB24A",
    x"BF7FB1FB",
    x"BF7FB1AD",
    x"BF7FB15E",
    x"BF7FB10F",
    x"BF7FB0C0",
    x"BF7FB071",
    x"BF7FB022",
    x"BF7FAFD2",
    x"BF7FAF83",
    x"BF7FAF33",
    x"BF7FAEE3",
    x"BF7FAE93",
    x"BF7FAE43",
    x"BF7FADF2",
    x"BF7FADA2",
    x"BF7FAD51",
    x"BF7FAD00",
    x"BF7FACAF",
    x"BF7FAC5E",
    x"BF7FAC0D",
    x"BF7FABBB",
    x"BF7FAB6A",
    x"BF7FAB18",
    x"BF7FAAC6",
    x"BF7FAA74",
    x"BF7FAA21",
    x"BF7FA9CF",
    x"BF7FA97D",
    x"BF7FA92A",
    x"BF7FA8D7",
    x"BF7FA884",
    x"BF7FA831",
    x"BF7FA7DE",
    x"BF7FA78A",
    x"BF7FA736",
    x"BF7FA6E3",
    x"BF7FA68F",
    x"BF7FA63B",
    x"BF7FA5E6",
    x"BF7FA592",
    x"BF7FA53D",
    x"BF7FA4E9",
    x"BF7FA494",
    x"BF7FA43F",
    x"BF7FA3EA",
    x"BF7FA394",
    x"BF7FA33F",
    x"BF7FA2E9",
    x"BF7FA294",
    x"BF7FA23E",
    x"BF7FA1E8",
    x"BF7FA191",
    x"BF7FA13B",
    x"BF7FA0E4",
    x"BF7FA08E",
    x"BF7FA037",
    x"BF7F9FE0",
    x"BF7F9F89",
    x"BF7F9F31",
    x"BF7F9EDA",
    x"BF7F9E82",
    x"BF7F9E2A",
    x"BF7F9DD2",
    x"BF7F9D7A",
    x"BF7F9D22",
    x"BF7F9CCA",
    x"BF7F9C71",
    x"BF7F9C18",
    x"BF7F9BC0",
    x"BF7F9B67",
    x"BF7F9B0D",
    x"BF7F9AB4",
    x"BF7F9A5B",
    x"BF7F9A01",
    x"BF7F99A7",
    x"BF7F994D",
    x"BF7F98F3",
    x"BF7F9899",
    x"BF7F983F",
    x"BF7F97E4",
    x"BF7F9789",
    x"BF7F972E",
    x"BF7F96D3",
    x"BF7F9678",
    x"BF7F961D",
    x"BF7F95C1",
    x"BF7F9566",
    x"BF7F950A",
    x"BF7F94AE",
    x"BF7F9452",
    x"BF7F93F6",
    x"BF7F9399",
    x"BF7F933D",
    x"BF7F92E0",
    x"BF7F9283",
    x"BF7F9226",
    x"BF7F91C9",
    x"BF7F916C",
    x"BF7F910E",
    x"BF7F90B1",
    x"BF7F9053",
    x"BF7F8FF5",
    x"BF7F8F97",
    x"BF7F8F39",
    x"BF7F8EDA",
    x"BF7F8E7C",
    x"BF7F8E1D",
    x"BF7F8DBE",
    x"BF7F8D5F",
    x"BF7F8D00",
    x"BF7F8CA1",
    x"BF7F8C41",
    x"BF7F8BE1",
    x"BF7F8B82",
    x"BF7F8B22",
    x"BF7F8AC2",
    x"BF7F8A61",
    x"BF7F8A01",
    x"BF7F89A0",
    x"BF7F8940",
    x"BF7F88DF",
    x"BF7F887E",
    x"BF7F881D",
    x"BF7F87BB",
    x"BF7F875A",
    x"BF7F86F8",
    x"BF7F8696",
    x"BF7F8634",
    x"BF7F85D2",
    x"BF7F8570",
    x"BF7F850E",
    x"BF7F84AB",
    x"BF7F8448",
    x"BF7F83E6",
    x"BF7F8383",
    x"BF7F831F",
    x"BF7F82BC",
    x"BF7F8259",
    x"BF7F81F5",
    x"BF7F8191",
    x"BF7F812D",
    x"BF7F80C9",
    x"BF7F8065",
    x"BF7F8000",
    x"BF7F7F9C",
    x"BF7F7F37",
    x"BF7F7ED2",
    x"BF7F7E6D",
    x"BF7F7E08",
    x"BF7F7DA3",
    x"BF7F7D3D",
    x"BF7F7CD8",
    x"BF7F7C72",
    x"BF7F7C0C",
    x"BF7F7BA6",
    x"BF7F7B40",
    x"BF7F7AD9",
    x"BF7F7A73",
    x"BF7F7A0C",
    x"BF7F79A5",
    x"BF7F793E",
    x"BF7F78D7",
    x"BF7F7870",
    x"BF7F7808",
    x"BF7F77A0",
    x"BF7F7739",
    x"BF7F76D1",
    x"BF7F7669",
    x"BF7F7600",
    x"BF7F7598",
    x"BF7F752F",
    x"BF7F74C7",
    x"BF7F745E",
    x"BF7F73F5",
    x"BF7F738C",
    x"BF7F7322",
    x"BF7F72B9",
    x"BF7F724F",
    x"BF7F71E5",
    x"BF7F717B",
    x"BF7F7111",
    x"BF7F70A7",
    x"BF7F703D",
    x"BF7F6FD2",
    x"BF7F6F67",
    x"BF7F6EFD",
    x"BF7F6E92",
    x"BF7F6E26",
    x"BF7F6DBB",
    x"BF7F6D50",
    x"BF7F6CE4",
    x"BF7F6C78",
    x"BF7F6C0C",
    x"BF7F6BA0",
    x"BF7F6B34",
    x"BF7F6AC7",
    x"BF7F6A5B",
    x"BF7F69EE",
    x"BF7F6981",
    x"BF7F6914",
    x"BF7F68A7",
    x"BF7F683A",
    x"BF7F67CC",
    x"BF7F675F",
    x"BF7F66F1",
    x"BF7F6683",
    x"BF7F6615",
    x"BF7F65A7",
    x"BF7F6538",
    x"BF7F64CA",
    x"BF7F645B",
    x"BF7F63EC",
    x"BF7F637D",
    x"BF7F630E",
    x"BF7F629E",
    x"BF7F622F",
    x"BF7F61BF",
    x"BF7F6150",
    x"BF7F60E0",
    x"BF7F606F",
    x"BF7F5FFF",
    x"BF7F5F8F",
    x"BF7F5F1E",
    x"BF7F5EAE",
    x"BF7F5E3D",
    x"BF7F5DCC",
    x"BF7F5D5A",
    x"BF7F5CE9",
    x"BF7F5C78",
    x"BF7F5C06",
    x"BF7F5B94",
    x"BF7F5B22",
    x"BF7F5AB0",
    x"BF7F5A3E",
    x"BF7F59CC",
    x"BF7F5959",
    x"BF7F58E6",
    x"BF7F5873",
    x"BF7F5800",
    x"BF7F578D",
    x"BF7F571A",
    x"BF7F56A6",
    x"BF7F5633",
    x"BF7F55BF",
    x"BF7F554B",
    x"BF7F54D7",
    x"BF7F5463",
    x"BF7F53EE",
    x"BF7F537A",
    x"BF7F5305",
    x"BF7F5290",
    x"BF7F521B",
    x"BF7F51A6",
    x"BF7F5131",
    x"BF7F50BB",
    x"BF7F5045",
    x"BF7F4FD0",
    x"BF7F4F5A",
    x"BF7F4EE4",
    x"BF7F4E6D",
    x"BF7F4DF7",
    x"BF7F4D80",
    x"BF7F4D0A",
    x"BF7F4C93",
    x"BF7F4C1C",
    x"BF7F4BA5",
    x"BF7F4B2D",
    x"BF7F4AB6",
    x"BF7F4A3E",
    x"BF7F49C6",
    x"BF7F494E",
    x"BF7F48D6",
    x"BF7F485E",
    x"BF7F47E6",
    x"BF7F476D",
    x"BF7F46F4",
    x"BF7F467C",
    x"BF7F4603",
    x"BF7F4589",
    x"BF7F4510",
    x"BF7F4497",
    x"BF7F441D",
    x"BF7F43A3",
    x"BF7F4329",
    x"BF7F42AF",
    x"BF7F4235",
    x"BF7F41BA",
    x"BF7F4140",
    x"BF7F40C5",
    x"BF7F404A",
    x"BF7F3FCF",
    x"BF7F3F54",
    x"BF7F3ED9",
    x"BF7F3E5D",
    x"BF7F3DE2",
    x"BF7F3D66",
    x"BF7F3CEA",
    x"BF7F3C6E",
    x"BF7F3BF2",
    x"BF7F3B75",
    x"BF7F3AF9",
    x"BF7F3A7C",
    x"BF7F39FF",
    x"BF7F3982",
    x"BF7F3905",
    x"BF7F3888",
    x"BF7F380A",
    x"BF7F378C",
    x"BF7F370F",
    x"BF7F3691",
    x"BF7F3613",
    x"BF7F3594",
    x"BF7F3516",
    x"BF7F3497",
    x"BF7F3419",
    x"BF7F339A",
    x"BF7F331B",
    x"BF7F329C",
    x"BF7F321C",
    x"BF7F319D",
    x"BF7F311D",
    x"BF7F309E",
    x"BF7F301E",
    x"BF7F2F9D",
    x"BF7F2F1D",
    x"BF7F2E9D",
    x"BF7F2E1C",
    x"BF7F2D9C",
    x"BF7F2D1B",
    x"BF7F2C9A",
    x"BF7F2C19",
    x"BF7F2B97",
    x"BF7F2B16",
    x"BF7F2A94",
    x"BF7F2A12",
    x"BF7F2990",
    x"BF7F290E",
    x"BF7F288C",
    x"BF7F280A",
    x"BF7F2787",
    x"BF7F2704",
    x"BF7F2682",
    x"BF7F25FF",
    x"BF7F257B",
    x"BF7F24F8",
    x"BF7F2475",
    x"BF7F23F1",
    x"BF7F236D",
    x"BF7F22E9",
    x"BF7F2265",
    x"BF7F21E1",
    x"BF7F215C",
    x"BF7F20D8",
    x"BF7F2053",
    x"BF7F1FCE",
    x"BF7F1F49",
    x"BF7F1EC4",
    x"BF7F1E3F",
    x"BF7F1DB9",
    x"BF7F1D34",
    x"BF7F1CAE",
    x"BF7F1C28",
    x"BF7F1BA2",
    x"BF7F1B1C",
    x"BF7F1A95",
    x"BF7F1A0F",
    x"BF7F1988",
    x"BF7F1901",
    x"BF7F187A",
    x"BF7F17F3",
    x"BF7F176C",
    x"BF7F16E4",
    x"BF7F165D",
    x"BF7F15D5",
    x"BF7F154D",
    x"BF7F14C5",
    x"BF7F143D",
    x"BF7F13B4",
    x"BF7F132C",
    x"BF7F12A3",
    x"BF7F121A",
    x"BF7F1191",
    x"BF7F1108",
    x"BF7F107F",
    x"BF7F0FF5",
    x"BF7F0F6C",
    x"BF7F0EE2",
    x"BF7F0E58",
    x"BF7F0DCE",
    x"BF7F0D44",
    x"BF7F0CB9",
    x"BF7F0C2F",
    x"BF7F0BA4",
    x"BF7F0B19",
    x"BF7F0A8E",
    x"BF7F0A03",
    x"BF7F0978",
    x"BF7F08EC",
    x"BF7F0861",
    x"BF7F07D5",
    x"BF7F0749",
    x"BF7F06BD",
    x"BF7F0631",
    x"BF7F05A4",
    x"BF7F0518",
    x"BF7F048B",
    x"BF7F03FE",
    x"BF7F0371",
    x"BF7F02E4",
    x"BF7F0257",
    x"BF7F01C9",
    x"BF7F013C",
    x"BF7F00AE",
    x"BF7F0020",
    x"BF7EFF92",
    x"BF7EFF04",
    x"BF7EFE75",
    x"BF7EFDE7",
    x"BF7EFD58",
    x"BF7EFCC9",
    x"BF7EFC3A",
    x"BF7EFBAB",
    x"BF7EFB1C",
    x"BF7EFA8C",
    x"BF7EF9FD",
    x"BF7EF96D",
    x"BF7EF8DD",
    x"BF7EF84D",
    x"BF7EF7BD",
    x"BF7EF72C",
    x"BF7EF69C",
    x"BF7EF60B",
    x"BF7EF57A",
    x"BF7EF4E9",
    x"BF7EF458",
    x"BF7EF3C7",
    x"BF7EF335",
    x"BF7EF2A4",
    x"BF7EF212",
    x"BF7EF180",
    x"BF7EF0EE",
    x"BF7EF05C",
    x"BF7EEFC9",
    x"BF7EEF37",
    x"BF7EEEA4",
    x"BF7EEE11",
    x"BF7EED7E",
    x"BF7EECEB",
    x"BF7EEC58",
    x"BF7EEBC4",
    x"BF7EEB31",
    x"BF7EEA9D",
    x"BF7EEA09",
    x"BF7EE975",
    x"BF7EE8E1",
    x"BF7EE84C",
    x"BF7EE7B8",
    x"BF7EE723",
    x"BF7EE68E",
    x"BF7EE5F9",
    x"BF7EE564",
    x"BF7EE4CF",
    x"BF7EE43A",
    x"BF7EE3A4",
    x"BF7EE30E",
    x"BF7EE278",
    x"BF7EE1E2",
    x"BF7EE14C",
    x"BF7EE0B6",
    x"BF7EE01F",
    x"BF7EDF88",
    x"BF7EDEF2",
    x"BF7EDE5B",
    x"BF7EDDC3",
    x"BF7EDD2C",
    x"BF7EDC95",
    x"BF7EDBFD",
    x"BF7EDB65",
    x"BF7EDACD",
    x"BF7EDA35",
    x"BF7ED99D",
    x"BF7ED905",
    x"BF7ED86C",
    x"BF7ED7D4",
    x"BF7ED73B",
    x"BF7ED6A2",
    x"BF7ED609",
    x"BF7ED56F",
    x"BF7ED4D6",
    x"BF7ED43C",
    x"BF7ED3A3",
    x"BF7ED309",
    x"BF7ED26F",
    x"BF7ED1D4",
    x"BF7ED13A",
    x"BF7ED0A0",
    x"BF7ED005",
    x"BF7ECF6A",
    x"BF7ECECF",
    x"BF7ECE34",
    x"BF7ECD99",
    x"BF7ECCFD",
    x"BF7ECC62",
    x"BF7ECBC6",
    x"BF7ECB2A",
    x"BF7ECA8E",
    x"BF7EC9F2",
    x"BF7EC955",
    x"BF7EC8B9",
    x"BF7EC81C",
    x"BF7EC780",
    x"BF7EC6E3",
    x"BF7EC645",
    x"BF7EC5A8",
    x"BF7EC50B",
    x"BF7EC46D",
    x"BF7EC3CF",
    x"BF7EC331",
    x"BF7EC293",
    x"BF7EC1F5",
    x"BF7EC157",
    x"BF7EC0B8",
    x"BF7EC01A",
    x"BF7EBF7B",
    x"BF7EBEDC",
    x"BF7EBE3D",
    x"BF7EBD9E",
    x"BF7EBCFE",
    x"BF7EBC5F",
    x"BF7EBBBF",
    x"BF7EBB1F",
    x"BF7EBA7F",
    x"BF7EB9DF",
    x"BF7EB93E",
    x"BF7EB89E",
    x"BF7EB7FD",
    x"BF7EB75C",
    x"BF7EB6BB",
    x"BF7EB61A",
    x"BF7EB579",
    x"BF7EB4D8",
    x"BF7EB436",
    x"BF7EB394",
    x"BF7EB2F2",
    x"BF7EB250",
    x"BF7EB1AE",
    x"BF7EB10C",
    x"BF7EB069",
    x"BF7EAFC7",
    x"BF7EAF24",
    x"BF7EAE81",
    x"BF7EADDE",
    x"BF7EAD3B",
    x"BF7EAC97",
    x"BF7EABF4",
    x"BF7EAB50",
    x"BF7EAAAC",
    x"BF7EAA08",
    x"BF7EA964",
    x"BF7EA8C0",
    x"BF7EA81B",
    x"BF7EA776",
    x"BF7EA6D2",
    x"BF7EA62D",
    x"BF7EA588",
    x"BF7EA4E2",
    x"BF7EA43D",
    x"BF7EA397",
    x"BF7EA2F2",
    x"BF7EA24C",
    x"BF7EA1A6",
    x"BF7EA100",
    x"BF7EA059",
    x"BF7E9FB3",
    x"BF7E9F0C",
    x"BF7E9E65",
    x"BF7E9DBE",
    x"BF7E9D17",
    x"BF7E9C70",
    x"BF7E9BC9",
    x"BF7E9B21",
    x"BF7E9A79",
    x"BF7E99D2",
    x"BF7E9929",
    x"BF7E9881",
    x"BF7E97D9",
    x"BF7E9731",
    x"BF7E9688",
    x"BF7E95DF",
    x"BF7E9536",
    x"BF7E948D",
    x"BF7E93E4",
    x"BF7E933A",
    x"BF7E9291",
    x"BF7E91E7",
    x"BF7E913D",
    x"BF7E9093",
    x"BF7E8FE9",
    x"BF7E8F3F",
    x"BF7E8E94",
    x"BF7E8DEA",
    x"BF7E8D3F",
    x"BF7E8C94",
    x"BF7E8BE9",
    x"BF7E8B3E",
    x"BF7E8A92",
    x"BF7E89E7",
    x"BF7E893B",
    x"BF7E888F",
    x"BF7E87E3",
    x"BF7E8737",
    x"BF7E868B",
    x"BF7E85DE",
    x"BF7E8532",
    x"BF7E8485",
    x"BF7E83D8",
    x"BF7E832B",
    x"BF7E827E",
    x"BF7E81D0",
    x"BF7E8123",
    x"BF7E8075",
    x"BF7E7FC7",
    x"BF7E7F19",
    x"BF7E7E6B",
    x"BF7E7DBD",
    x"BF7E7D0E",
    x"BF7E7C60",
    x"BF7E7BB1",
    x"BF7E7B02",
    x"BF7E7A53",
    x"BF7E79A4",
    x"BF7E78F4",
    x"BF7E7845",
    x"BF7E7795",
    x"BF7E76E5",
    x"BF7E7635",
    x"BF7E7585",
    x"BF7E74D5",
    x"BF7E7424",
    x"BF7E7374",
    x"BF7E72C3",
    x"BF7E7212",
    x"BF7E7161",
    x"BF7E70B0",
    x"BF7E6FFF",
    x"BF7E6F4D",
    x"BF7E6E9B",
    x"BF7E6DEA",
    x"BF7E6D38",
    x"BF7E6C85",
    x"BF7E6BD3",
    x"BF7E6B21",
    x"BF7E6A6E",
    x"BF7E69BB",
    x"BF7E6908",
    x"BF7E6855",
    x"BF7E67A2",
    x"BF7E66EF",
    x"BF7E663B",
    x"BF7E6588",
    x"BF7E64D4",
    x"BF7E6420",
    x"BF7E636C",
    x"BF7E62B7",
    x"BF7E6203",
    x"BF7E614E",
    x"BF7E609A",
    x"BF7E5FE5",
    x"BF7E5F30",
    x"BF7E5E7B",
    x"BF7E5DC5",
    x"BF7E5D10",
    x"BF7E5C5A",
    x"BF7E5BA4",
    x"BF7E5AEE",
    x"BF7E5A38",
    x"BF7E5982",
    x"BF7E58CB",
    x"BF7E5815",
    x"BF7E575E",
    x"BF7E56A7",
    x"BF7E55F0",
    x"BF7E5539",
    x"BF7E5482",
    x"BF7E53CA",
    x"BF7E5312",
    x"BF7E525B",
    x"BF7E51A3",
    x"BF7E50EB",
    x"BF7E5032",
    x"BF7E4F7A",
    x"BF7E4EC1",
    x"BF7E4E09",
    x"BF7E4D50",
    x"BF7E4C97",
    x"BF7E4BDE",
    x"BF7E4B24",
    x"BF7E4A6B",
    x"BF7E49B1",
    x"BF7E48F7",
    x"BF7E483D",
    x"BF7E4783",
    x"BF7E46C9",
    x"BF7E460F",
    x"BF7E4554",
    x"BF7E4499",
    x"BF7E43DE",
    x"BF7E4323",
    x"BF7E4268",
    x"BF7E41AD",
    x"BF7E40F1",
    x"BF7E4036",
    x"BF7E3F7A",
    x"BF7E3EBE",
    x"BF7E3E02",
    x"BF7E3D46",
    x"BF7E3C89",
    x"BF7E3BCD",
    x"BF7E3B10",
    x"BF7E3A53",
    x"BF7E3996",
    x"BF7E38D9",
    x"BF7E381C",
    x"BF7E375E",
    x"BF7E36A1",
    x"BF7E35E3",
    x"BF7E3525",
    x"BF7E3467",
    x"BF7E33A9",
    x"BF7E32EA",
    x"BF7E322C",
    x"BF7E316D",
    x"BF7E30AE",
    x"BF7E2FEF",
    x"BF7E2F30",
    x"BF7E2E71",
    x"BF7E2DB1",
    x"BF7E2CF2",
    x"BF7E2C32",
    x"BF7E2B72",
    x"BF7E2AB2",
    x"BF7E29F2",
    x"BF7E2931",
    x"BF7E2871",
    x"BF7E27B0",
    x"BF7E26EF",
    x"BF7E262E",
    x"BF7E256D",
    x"BF7E24AC",
    x"BF7E23EA",
    x"BF7E2329",
    x"BF7E2267",
    x"BF7E21A5",
    x"BF7E20E3",
    x"BF7E2021",
    x"BF7E1F5E",
    x"BF7E1E9C",
    x"BF7E1DD9",
    x"BF7E1D16",
    x"BF7E1C53",
    x"BF7E1B90",
    x"BF7E1ACD",
    x"BF7E1A09",
    x"BF7E1946",
    x"BF7E1882",
    x"BF7E17BE",
    x"BF7E16FA",
    x"BF7E1636",
    x"BF7E1572",
    x"BF7E14AD",
    x"BF7E13E8",
    x"BF7E1324",
    x"BF7E125F",
    x"BF7E1199",
    x"BF7E10D4",
    x"BF7E100F",
    x"BF7E0F49",
    x"BF7E0E83",
    x"BF7E0DBD",
    x"BF7E0CF7",
    x"BF7E0C31",
    x"BF7E0B6B",
    x"BF7E0AA4",
    x"BF7E09DE",
    x"BF7E0917",
    x"BF7E0850",
    x"BF7E0789",
    x"BF7E06C2",
    x"BF7E05FA",
    x"BF7E0533",
    x"BF7E046B",
    x"BF7E03A3",
    x"BF7E02DB",
    x"BF7E0213",
    x"BF7E014A",
    x"BF7E0082",
    x"BF7DFFB9",
    x"BF7DFEF0",
    x"BF7DFE28",
    x"BF7DFD5E",
    x"BF7DFC95",
    x"BF7DFBCC",
    x"BF7DFB02",
    x"BF7DFA38",
    x"BF7DF96F",
    x"BF7DF8A5",
    x"BF7DF7DA",
    x"BF7DF710",
    x"BF7DF646",
    x"BF7DF57B",
    x"BF7DF4B0",
    x"BF7DF3E5",
    x"BF7DF31A",
    x"BF7DF24F",
    x"BF7DF183",
    x"BF7DF0B8",
    x"BF7DEFEC",
    x"BF7DEF20",
    x"BF7DEE54",
    x"BF7DED88",
    x"BF7DECBC",
    x"BF7DEBEF",
    x"BF7DEB23",
    x"BF7DEA56",
    x"BF7DE989",
    x"BF7DE8BC",
    x"BF7DE7EF",
    x"BF7DE721",
    x"BF7DE654",
    x"BF7DE586",
    x"BF7DE4B8",
    x"BF7DE3EA",
    x"BF7DE31C",
    x"BF7DE24E",
    x"BF7DE17F",
    x"BF7DE0B1",
    x"BF7DDFE2",
    x"BF7DDF13",
    x"BF7DDE44",
    x"BF7DDD75",
    x"BF7DDCA5",
    x"BF7DDBD6",
    x"BF7DDB06",
    x"BF7DDA36",
    x"BF7DD966",
    x"BF7DD896",
    x"BF7DD7C6",
    x"BF7DD6F5",
    x"BF7DD625",
    x"BF7DD554",
    x"BF7DD483",
    x"BF7DD3B2",
    x"BF7DD2E1",
    x"BF7DD210",
    x"BF7DD13E",
    x"BF7DD06C",
    x"BF7DCF9B",
    x"BF7DCEC9",
    x"BF7DCDF6",
    x"BF7DCD24",
    x"BF7DCC52",
    x"BF7DCB7F",
    x"BF7DCAAC",
    x"BF7DC9DA",
    x"BF7DC906",
    x"BF7DC833",
    x"BF7DC760",
    x"BF7DC68C",
    x"BF7DC5B9",
    x"BF7DC4E5",
    x"BF7DC411",
    x"BF7DC33D",
    x"BF7DC269",
    x"BF7DC194",
    x"BF7DC0C0",
    x"BF7DBFEB",
    x"BF7DBF16",
    x"BF7DBE41",
    x"BF7DBD6C",
    x"BF7DBC96",
    x"BF7DBBC1",
    x"BF7DBAEB",
    x"BF7DBA15",
    x"BF7DB940",
    x"BF7DB869",
    x"BF7DB793",
    x"BF7DB6BD",
    x"BF7DB5E6",
    x"BF7DB510",
    x"BF7DB439",
    x"BF7DB362",
    x"BF7DB28A",
    x"BF7DB1B3",
    x"BF7DB0DC",
    x"BF7DB004",
    x"BF7DAF2C",
    x"BF7DAE54",
    x"BF7DAD7C",
    x"BF7DACA4",
    x"BF7DABCC",
    x"BF7DAAF3",
    x"BF7DAA1A",
    x"BF7DA941",
    x"BF7DA868",
    x"BF7DA78F",
    x"BF7DA6B6",
    x"BF7DA5DC",
    x"BF7DA503",
    x"BF7DA429",
    x"BF7DA34F",
    x"BF7DA275",
    x"BF7DA19B",
    x"BF7DA0C0",
    x"BF7D9FE6",
    x"BF7D9F0B",
    x"BF7D9E30",
    x"BF7D9D55",
    x"BF7D9C7A",
    x"BF7D9B9F",
    x"BF7D9AC4",
    x"BF7D99E8",
    x"BF7D990C",
    x"BF7D9830",
    x"BF7D9754",
    x"BF7D9678",
    x"BF7D959C",
    x"BF7D94BF",
    x"BF7D93E2",
    x"BF7D9306",
    x"BF7D9229",
    x"BF7D914B",
    x"BF7D906E",
    x"BF7D8F91",
    x"BF7D8EB3",
    x"BF7D8DD5",
    x"BF7D8CF8",
    x"BF7D8C19",
    x"BF7D8B3B",
    x"BF7D8A5D",
    x"BF7D897E",
    x"BF7D88A0",
    x"BF7D87C1",
    x"BF7D86E2",
    x"BF7D8603",
    x"BF7D8524",
    x"BF7D8444",
    x"BF7D8365",
    x"BF7D8285",
    x"BF7D81A5",
    x"BF7D80C5",
    x"BF7D7FE5",
    x"BF7D7F04",
    x"BF7D7E24",
    x"BF7D7D43",
    x"BF7D7C62",
    x"BF7D7B82",
    x"BF7D7AA0",
    x"BF7D79BF",
    x"BF7D78DE",
    x"BF7D77FC",
    x"BF7D771B",
    x"BF7D7639",
    x"BF7D7557",
    x"BF7D7474",
    x"BF7D7392",
    x"BF7D72B0",
    x"BF7D71CD",
    x"BF7D70EA",
    x"BF7D7007",
    x"BF7D6F24",
    x"BF7D6E41",
    x"BF7D6D5E",
    x"BF7D6C7A",
    x"BF7D6B96",
    x"BF7D6AB2",
    x"BF7D69CE",
    x"BF7D68EA",
    x"BF7D6806",
    x"BF7D6722",
    x"BF7D663D",
    x"BF7D6558",
    x"BF7D6473",
    x"BF7D638E",
    x"BF7D62A9",
    x"BF7D61C4",
    x"BF7D60DE",
    x"BF7D5FF8",
    x"BF7D5F13",
    x"BF7D5E2D",
    x"BF7D5D46",
    x"BF7D5C60",
    x"BF7D5B7A",
    x"BF7D5A93",
    x"BF7D59AC",
    x"BF7D58C5",
    x"BF7D57DE",
    x"BF7D56F7",
    x"BF7D5610",
    x"BF7D5528",
    x"BF7D5441",
    x"BF7D5359",
    x"BF7D5271",
    x"BF7D5189",
    x"BF7D50A0",
    x"BF7D4FB8",
    x"BF7D4ECF",
    x"BF7D4DE7",
    x"BF7D4CFE",
    x"BF7D4C15",
    x"BF7D4B2C",
    x"BF7D4A42",
    x"BF7D4959",
    x"BF7D486F",
    x"BF7D4785",
    x"BF7D469B",
    x"BF7D45B1",
    x"BF7D44C7",
    x"BF7D43DC",
    x"BF7D42F2",
    x"BF7D4207",
    x"BF7D411C",
    x"BF7D4031",
    x"BF7D3F46",
    x"BF7D3E5B",
    x"BF7D3D6F",
    x"BF7D3C84",
    x"BF7D3B98",
    x"BF7D3AAC",
    x"BF7D39C0",
    x"BF7D38D4",
    x"BF7D37E7",
    x"BF7D36FB",
    x"BF7D360E",
    x"BF7D3521",
    x"BF7D3434",
    x"BF7D3347",
    x"BF7D325A",
    x"BF7D316C",
    x"BF7D307F",
    x"BF7D2F91",
    x"BF7D2EA3",
    x"BF7D2DB5",
    x"BF7D2CC7",
    x"BF7D2BD8",
    x"BF7D2AEA",
    x"BF7D29FB",
    x"BF7D290C",
    x"BF7D281D",
    x"BF7D272E",
    x"BF7D263F",
    x"BF7D254F",
    x"BF7D2460",
    x"BF7D2370",
    x"BF7D2280",
    x"BF7D2190",
    x"BF7D20A0",
    x"BF7D1FAF",
    x"BF7D1EBF",
    x"BF7D1DCE",
    x"BF7D1CDD",
    x"BF7D1BEC",
    x"BF7D1AFB",
    x"BF7D1A0A",
    x"BF7D1919",
    x"BF7D1827",
    x"BF7D1735",
    x"BF7D1643",
    x"BF7D1551",
    x"BF7D145F",
    x"BF7D136D",
    x"BF7D127A",
    x"BF7D1188",
    x"BF7D1095",
    x"BF7D0FA2",
    x"BF7D0EAF",
    x"BF7D0DBC",
    x"BF7D0CC8",
    x"BF7D0BD5",
    x"BF7D0AE1",
    x"BF7D09ED",
    x"BF7D08F9",
    x"BF7D0805",
    x"BF7D0710",
    x"BF7D061C",
    x"BF7D0527",
    x"BF7D0433",
    x"BF7D033E",
    x"BF7D0249",
    x"BF7D0153",
    x"BF7D005E",
    x"BF7CFF68",
    x"BF7CFE73",
    x"BF7CFD7D",
    x"BF7CFC87",
    x"BF7CFB91",
    x"BF7CFA9A",
    x"BF7CF9A4",
    x"BF7CF8AD",
    x"BF7CF7B7",
    x"BF7CF6C0",
    x"BF7CF5C9",
    x"BF7CF4D1",
    x"BF7CF3DA",
    x"BF7CF2E2",
    x"BF7CF1EB",
    x"BF7CF0F3",
    x"BF7CEFFB",
    x"BF7CEF03",
    x"BF7CEE0B",
    x"BF7CED12",
    x"BF7CEC19",
    x"BF7CEB21",
    x"BF7CEA28",
    x"BF7CE92F",
    x"BF7CE836",
    x"BF7CE73C",
    x"BF7CE643",
    x"BF7CE549",
    x"BF7CE44F",
    x"BF7CE355",
    x"BF7CE25B",
    x"BF7CE161",
    x"BF7CE066",
    x"BF7CDF6C",
    x"BF7CDE71",
    x"BF7CDD76",
    x"BF7CDC7B",
    x"BF7CDB80",
    x"BF7CDA85",
    x"BF7CD989",
    x"BF7CD88E",
    x"BF7CD792",
    x"BF7CD696",
    x"BF7CD59A",
    x"BF7CD49E",
    x"BF7CD3A1",
    x"BF7CD2A5",
    x"BF7CD1A8",
    x"BF7CD0AB",
    x"BF7CCFAE",
    x"BF7CCEB1",
    x"BF7CCDB4",
    x"BF7CCCB6",
    x"BF7CCBB8",
    x"BF7CCABB",
    x"BF7CC9BD",
    x"BF7CC8BF",
    x"BF7CC7C0",
    x"BF7CC6C2",
    x"BF7CC5C4",
    x"BF7CC4C5",
    x"BF7CC3C6",
    x"BF7CC2C7",
    x"BF7CC1C8",
    x"BF7CC0C9",
    x"BF7CBFC9",
    x"BF7CBECA",
    x"BF7CBDCA",
    x"BF7CBCCA",
    x"BF7CBBCA",
    x"BF7CBACA",
    x"BF7CB9C9",
    x"BF7CB8C9",
    x"BF7CB7C8",
    x"BF7CB6C7",
    x"BF7CB5C6",
    x"BF7CB4C5",
    x"BF7CB3C4",
    x"BF7CB2C2",
    x"BF7CB1C1",
    x"BF7CB0BF",
    x"BF7CAFBD",
    x"BF7CAEBB",
    x"BF7CADB9",
    x"BF7CACB7",
    x"BF7CABB4",
    x"BF7CAAB2",
    x"BF7CA9AF",
    x"BF7CA8AC",
    x"BF7CA7A9",
    x"BF7CA6A6",
    x"BF7CA5A2",
    x"BF7CA49F",
    x"BF7CA39B",
    x"BF7CA297",
    x"BF7CA193",
    x"BF7CA08F",
    x"BF7C9F8A",
    x"BF7C9E86",
    x"BF7C9D81",
    x"BF7C9C7D",
    x"BF7C9B78",
    x"BF7C9A73",
    x"BF7C996D",
    x"BF7C9868",
    x"BF7C9762",
    x"BF7C965D",
    x"BF7C9557",
    x"BF7C9451",
    x"BF7C934B",
    x"BF7C9245",
    x"BF7C913E",
    x"BF7C9037",
    x"BF7C8F31",
    x"BF7C8E2A",
    x"BF7C8D23",
    x"BF7C8C1C",
    x"BF7C8B14",
    x"BF7C8A0D",
    x"BF7C8905",
    x"BF7C87FD",
    x"BF7C86F5",
    x"BF7C85ED",
    x"BF7C84E5",
    x"BF7C83DC",
    x"BF7C82D4",
    x"BF7C81CB",
    x"BF7C80C2",
    x"BF7C7FB9",
    x"BF7C7EB0",
    x"BF7C7DA7",
    x"BF7C7C9D",
    x"BF7C7B94",
    x"BF7C7A8A",
    x"BF7C7980",
    x"BF7C7876",
    x"BF7C776B",
    x"BF7C7661",
    x"BF7C7556",
    x"BF7C744C",
    x"BF7C7341",
    x"BF7C7236",
    x"BF7C712B",
    x"BF7C701F",
    x"BF7C6F14",
    x"BF7C6E08",
    x"BF7C6CFD",
    x"BF7C6BF1",
    x"BF7C6AE5",
    x"BF7C69D8",
    x"BF7C68CC",
    x"BF7C67BF",
    x"BF7C66B3",
    x"BF7C65A6",
    x"BF7C6499",
    x"BF7C638C",
    x"BF7C627E",
    x"BF7C6171",
    x"BF7C6063",
    x"BF7C5F56",
    x"BF7C5E48",
    x"BF7C5D3A",
    x"BF7C5C2C",
    x"BF7C5B1D",
    x"BF7C5A0F",
    x"BF7C5900",
    x"BF7C57F1",
    x"BF7C56E2",
    x"BF7C55D3",
    x"BF7C54C4",
    x"BF7C53B4",
    x"BF7C52A5",
    x"BF7C5195",
    x"BF7C5085",
    x"BF7C4F75",
    x"BF7C4E65",
    x"BF7C4D55",
    x"BF7C4C44",
    x"BF7C4B34",
    x"BF7C4A23",
    x"BF7C4912",
    x"BF7C4801",
    x"BF7C46F0",
    x"BF7C45DE",
    x"BF7C44CD",
    x"BF7C43BB",
    x"BF7C42A9",
    x"BF7C4197",
    x"BF7C4085",
    x"BF7C3F73",
    x"BF7C3E60",
    x"BF7C3D4E",
    x"BF7C3C3B",
    x"BF7C3B28",
    x"BF7C3A15",
    x"BF7C3902",
    x"BF7C37EE",
    x"BF7C36DB",
    x"BF7C35C7",
    x"BF7C34B3",
    x"BF7C339F",
    x"BF7C328B",
    x"BF7C3177",
    x"BF7C3062",
    x"BF7C2F4E",
    x"BF7C2E39",
    x"BF7C2D24",
    x"BF7C2C0F",
    x"BF7C2AFA",
    x"BF7C29E5",
    x"BF7C28CF",
    x"BF7C27B9",
    x"BF7C26A4",
    x"BF7C258E",
    x"BF7C2478",
    x"BF7C2361",
    x"BF7C224B",
    x"BF7C2134",
    x"BF7C201E",
    x"BF7C1F07",
    x"BF7C1DF0",
    x"BF7C1CD9",
    x"BF7C1BC1",
    x"BF7C1AAA",
    x"BF7C1992",
    x"BF7C187A",
    x"BF7C1762",
    x"BF7C164A",
    x"BF7C1532",
    x"BF7C141A",
    x"BF7C1301",
    x"BF7C11E8",
    x"BF7C10D0",
    x"BF7C0FB7",
    x"BF7C0E9D",
    x"BF7C0D84",
    x"BF7C0C6B",
    x"BF7C0B51",
    x"BF7C0A37",
    x"BF7C091E",
    x"BF7C0803",
    x"BF7C06E9",
    x"BF7C05CF",
    x"BF7C04B4",
    x"BF7C039A",
    x"BF7C027F",
    x"BF7C0164",
    x"BF7C0049",
    x"BF7BFF2E",
    x"BF7BFE12",
    x"BF7BFCF7",
    x"BF7BFBDB",
    x"BF7BFABF",
    x"BF7BF9A3",
    x"BF7BF887",
    x"BF7BF76A",
    x"BF7BF64E",
    x"BF7BF531",
    x"BF7BF415",
    x"BF7BF2F8",
    x"BF7BF1DA",
    x"BF7BF0BD",
    x"BF7BEFA0",
    x"BF7BEE82",
    x"BF7BED65",
    x"BF7BEC47",
    x"BF7BEB29",
    x"BF7BEA0B",
    x"BF7BE8EC",
    x"BF7BE7CE",
    x"BF7BE6AF",
    x"BF7BE590",
    x"BF7BE472",
    x"BF7BE353",
    x"BF7BE233",
    x"BF7BE114",
    x"BF7BDFF4",
    x"BF7BDED5",
    x"BF7BDDB5",
    x"BF7BDC95",
    x"BF7BDB75",
    x"BF7BDA55",
    x"BF7BD934",
    x"BF7BD814",
    x"BF7BD6F3",
    x"BF7BD5D2",
    x"BF7BD4B1",
    x"BF7BD390",
    x"BF7BD26E",
    x"BF7BD14D",
    x"BF7BD02B",
    x"BF7BCF09",
    x"BF7BCDE7",
    x"BF7BCCC5",
    x"BF7BCBA3",
    x"BF7BCA81",
    x"BF7BC95E",
    x"BF7BC83B",
    x"BF7BC719",
    x"BF7BC5F6",
    x"BF7BC4D2",
    x"BF7BC3AF",
    x"BF7BC28C",
    x"BF7BC168",
    x"BF7BC044",
    x"BF7BBF20",
    x"BF7BBDFC",
    x"BF7BBCD8",
    x"BF7BBBB4",
    x"BF7BBA8F",
    x"BF7BB96B",
    x"BF7BB846",
    x"BF7BB721",
    x"BF7BB5FC",
    x"BF7BB4D6",
    x"BF7BB3B1",
    x"BF7BB28B",
    x"BF7BB166",
    x"BF7BB040",
    x"BF7BAF1A",
    x"BF7BADF3",
    x"BF7BACCD",
    x"BF7BABA7",
    x"BF7BAA80",
    x"BF7BA959",
    x"BF7BA832",
    x"BF7BA70B",
    x"BF7BA5E4",
    x"BF7BA4BC",
    x"BF7BA395",
    x"BF7BA26D",
    x"BF7BA145",
    x"BF7BA01D",
    x"BF7B9EF5",
    x"BF7B9DCD",
    x"BF7B9CA4",
    x"BF7B9B7C",
    x"BF7B9A53",
    x"BF7B992A",
    x"BF7B9801",
    x"BF7B96D8",
    x"BF7B95AE",
    x"BF7B9485",
    x"BF7B935B",
    x"BF7B9231",
    x"BF7B9107",
    x"BF7B8FDD",
    x"BF7B8EB3",
    x"BF7B8D89",
    x"BF7B8C5E",
    x"BF7B8B33",
    x"BF7B8A08",
    x"BF7B88DD",
    x"BF7B87B2",
    x"BF7B8687",
    x"BF7B855B",
    x"BF7B8430",
    x"BF7B8304",
    x"BF7B81D8",
    x"BF7B80AC",
    x"BF7B7F80",
    x"BF7B7E53",
    x"BF7B7D27",
    x"BF7B7BFA",
    x"BF7B7ACD",
    x"BF7B79A0",
    x"BF7B7873",
    x"BF7B7745",
    x"BF7B7618",
    x"BF7B74EA",
    x"BF7B73BD",
    x"BF7B728F",
    x"BF7B7161",
    x"BF7B7032",
    x"BF7B6F04",
    x"BF7B6DD6",
    x"BF7B6CA7",
    x"BF7B6B78",
    x"BF7B6A49",
    x"BF7B691A",
    x"BF7B67EB",
    x"BF7B66BB",
    x"BF7B658C",
    x"BF7B645C",
    x"BF7B632C",
    x"BF7B61FC",
    x"BF7B60CC",
    x"BF7B5F9B",
    x"BF7B5E6B",
    x"BF7B5D3A",
    x"BF7B5C09",
    x"BF7B5AD9",
    x"BF7B59A7",
    x"BF7B5876",
    x"BF7B5745",
    x"BF7B5613",
    x"BF7B54E1",
    x"BF7B53B0",
    x"BF7B527E",
    x"BF7B514B",
    x"BF7B5019",
    x"BF7B4EE7",
    x"BF7B4DB4",
    x"BF7B4C81",
    x"BF7B4B4E",
    x"BF7B4A1B",
    x"BF7B48E8",
    x"BF7B47B5",
    x"BF7B4681",
    x"BF7B454E",
    x"BF7B441A",
    x"BF7B42E6",
    x"BF7B41B2",
    x"BF7B407D",
    x"BF7B3F49",
    x"BF7B3E14",
    x"BF7B3CE0",
    x"BF7B3BAB",
    x"BF7B3A76",
    x"BF7B3940",
    x"BF7B380B",
    x"BF7B36D6",
    x"BF7B35A0",
    x"BF7B346A",
    x"BF7B3334",
    x"BF7B31FE",
    x"BF7B30C8",
    x"BF7B2F92",
    x"BF7B2E5B",
    x"BF7B2D24",
    x"BF7B2BED",
    x"BF7B2AB6",
    x"BF7B297F",
    x"BF7B2848",
    x"BF7B2711",
    x"BF7B25D9",
    x"BF7B24A1",
    x"BF7B2369",
    x"BF7B2231",
    x"BF7B20F9",
    x"BF7B1FC1",
    x"BF7B1E88",
    x"BF7B1D4F",
    x"BF7B1C17",
    x"BF7B1ADE",
    x"BF7B19A4",
    x"BF7B186B",
    x"BF7B1732",
    x"BF7B15F8",
    x"BF7B14BE",
    x"BF7B1385",
    x"BF7B124B",
    x"BF7B1110",
    x"BF7B0FD6",
    x"BF7B0E9C",
    x"BF7B0D61",
    x"BF7B0C26",
    x"BF7B0AEB",
    x"BF7B09B0",
    x"BF7B0875",
    x"BF7B073A",
    x"BF7B05FE",
    x"BF7B04C2",
    x"BF7B0386",
    x"BF7B024A",
    x"BF7B010E",
    x"BF7AFFD2",
    x"BF7AFE96",
    x"BF7AFD59",
    x"BF7AFC1C",
    x"BF7AFADF",
    x"BF7AF9A2",
    x"BF7AF865",
    x"BF7AF728",
    x"BF7AF5EA",
    x"BF7AF4AD",
    x"BF7AF36F",
    x"BF7AF231",
    x"BF7AF0F3",
    x"BF7AEFB4",
    x"BF7AEE76",
    x"BF7AED37",
    x"BF7AEBF9",
    x"BF7AEABA",
    x"BF7AE97B",
    x"BF7AE83C",
    x"BF7AE6FC",
    x"BF7AE5BD",
    x"BF7AE47D",
    x"BF7AE33D",
    x"BF7AE1FE",
    x"BF7AE0BD",
    x"BF7ADF7D",
    x"BF7ADE3D",
    x"BF7ADCFC",
    x"BF7ADBBC",
    x"BF7ADA7B",
    x"BF7AD93A",
    x"BF7AD7F9",
    x"BF7AD6B7",
    x"BF7AD576",
    x"BF7AD434",
    x"BF7AD2F3",
    x"BF7AD1B1",
    x"BF7AD06F",
    x"BF7ACF2D",
    x"BF7ACDEA",
    x"BF7ACCA8",
    x"BF7ACB65",
    x"BF7ACA22",
    x"BF7AC8DF",
    x"BF7AC79C",
    x"BF7AC659",
    x"BF7AC516",
    x"BF7AC3D2",
    x"BF7AC28E",
    x"BF7AC14A",
    x"BF7AC006",
    x"BF7ABEC2",
    x"BF7ABD7E",
    x"BF7ABC3A",
    x"BF7ABAF5",
    x"BF7AB9B0",
    x"BF7AB86B",
    x"BF7AB726",
    x"BF7AB5E1",
    x"BF7AB49C",
    x"BF7AB356",
    x"BF7AB210",
    x"BF7AB0CB",
    x"BF7AAF85",
    x"BF7AAE3F",
    x"BF7AACF8",
    x"BF7AABB2",
    x"BF7AAA6B",
    x"BF7AA925",
    x"BF7AA7DE",
    x"BF7AA697",
    x"BF7AA54F",
    x"BF7AA408",
    x"BF7AA2C1",
    x"BF7AA179",
    x"BF7AA031",
    x"BF7A9EE9",
    x"BF7A9DA1",
    x"BF7A9C59",
    x"BF7A9B11",
    x"BF7A99C8",
    x"BF7A987F",
    x"BF7A9737",
    x"BF7A95EE",
    x"BF7A94A4",
    x"BF7A935B",
    x"BF7A9212",
    x"BF7A90C8",
    x"BF7A8F7E",
    x"BF7A8E34",
    x"BF7A8CEA",
    x"BF7A8BA0",
    x"BF7A8A56",
    x"BF7A890B",
    x"BF7A87C1",
    x"BF7A8676",
    x"BF7A852B",
    x"BF7A83E0",
    x"BF7A8295",
    x"BF7A8149",
    x"BF7A7FFE",
    x"BF7A7EB2",
    x"BF7A7D66",
    x"BF7A7C1A",
    x"BF7A7ACE",
    x"BF7A7982",
    x"BF7A7835",
    x"BF7A76E9",
    x"BF7A759C",
    x"BF7A744F",
    x"BF7A7302",
    x"BF7A71B5",
    x"BF7A7067",
    x"BF7A6F1A",
    x"BF7A6DCC",
    x"BF7A6C7E",
    x"BF7A6B30",
    x"BF7A69E2",
    x"BF7A6894",
    x"BF7A6745",
    x"BF7A65F7",
    x"BF7A64A8",
    x"BF7A6359",
    x"BF7A620A",
    x"BF7A60BB",
    x"BF7A5F6C",
    x"BF7A5E1C",
    x"BF7A5CCD",
    x"BF7A5B7D",
    x"BF7A5A2D",
    x"BF7A58DD",
    x"BF7A578D",
    x"BF7A563C",
    x"BF7A54EC",
    x"BF7A539B",
    x"BF7A524A",
    x"BF7A50F9",
    x"BF7A4FA8",
    x"BF7A4E57",
    x"BF7A4D05",
    x"BF7A4BB4",
    x"BF7A4A62",
    x"BF7A4910",
    x"BF7A47BE",
    x"BF7A466C",
    x"BF7A451A",
    x"BF7A43C7",
    x"BF7A4275",
    x"BF7A4122",
    x"BF7A3FCF",
    x"BF7A3E7C",
    x"BF7A3D28",
    x"BF7A3BD5",
    x"BF7A3A81",
    x"BF7A392E",
    x"BF7A37DA",
    x"BF7A3686",
    x"BF7A3532",
    x"BF7A33DD",
    x"BF7A3289",
    x"BF7A3134",
    x"BF7A2FE0",
    x"BF7A2E8B",
    x"BF7A2D36",
    x"BF7A2BE1",
    x"BF7A2A8B",
    x"BF7A2936",
    x"BF7A27E0",
    x"BF7A268A",
    x"BF7A2534",
    x"BF7A23DE",
    x"BF7A2288",
    x"BF7A2131",
    x"BF7A1FDB",
    x"BF7A1E84",
    x"BF7A1D2D",
    x"BF7A1BD6",
    x"BF7A1A7F",
    x"BF7A1928",
    x"BF7A17D0",
    x"BF7A1679",
    x"BF7A1521",
    x"BF7A13C9",
    x"BF7A1271",
    x"BF7A1119",
    x"BF7A0FC0",
    x"BF7A0E68",
    x"BF7A0D0F",
    x"BF7A0BB6",
    x"BF7A0A5D",
    x"BF7A0904",
    x"BF7A07AB",
    x"BF7A0652",
    x"BF7A04F8",
    x"BF7A039E",
    x"BF7A0244",
    x"BF7A00EA",
    x"BF79FF90",
    x"BF79FE36",
    x"BF79FCDB",
    x"BF79FB81",
    x"BF79FA26",
    x"BF79F8CB",
    x"BF79F770",
    x"BF79F615",
    x"BF79F4B9",
    x"BF79F35E",
    x"BF79F202",
    x"BF79F0A6",
    x"BF79EF4A",
    x"BF79EDEE",
    x"BF79EC92",
    x"BF79EB36",
    x"BF79E9D9",
    x"BF79E87C",
    x"BF79E71F",
    x"BF79E5C2",
    x"BF79E465",
    x"BF79E308",
    x"BF79E1AA",
    x"BF79E04D",
    x"BF79DEEF",
    x"BF79DD91",
    x"BF79DC33",
    x"BF79DAD5",
    x"BF79D976",
    x"BF79D818",
    x"BF79D6B9",
    x"BF79D55A",
    x"BF79D3FB",
    x"BF79D29C",
    x"BF79D13D",
    x"BF79CFDD",
    x"BF79CE7E",
    x"BF79CD1E",
    x"BF79CBBE",
    x"BF79CA5E",
    x"BF79C8FE",
    x"BF79C79D",
    x"BF79C63D",
    x"BF79C4DC",
    x"BF79C37B",
    x"BF79C21A",
    x"BF79C0B9",
    x"BF79BF58",
    x"BF79BDF7",
    x"BF79BC95",
    x"BF79BB33",
    x"BF79B9D2",
    x"BF79B870",
    x"BF79B70D",
    x"BF79B5AB",
    x"BF79B449",
    x"BF79B2E6",
    x"BF79B183",
    x"BF79B020",
    x"BF79AEBD",
    x"BF79AD5A",
    x"BF79ABF7",
    x"BF79AA93",
    x"BF79A930",
    x"BF79A7CC",
    x"BF79A668",
    x"BF79A504",
    x"BF79A3A0",
    x"BF79A23B",
    x"BF79A0D7",
    x"BF799F72",
    x"BF799E0D",
    x"BF799CA8",
    x"BF799B43",
    x"BF7999DE",
    x"BF799878",
    x"BF799712",
    x"BF7995AD",
    x"BF799447",
    x"BF7992E1",
    x"BF79917A",
    x"BF799014",
    x"BF798EAE",
    x"BF798D47",
    x"BF798BE0",
    x"BF798A79",
    x"BF798912",
    x"BF7987AB",
    x"BF798643",
    x"BF7984DC",
    x"BF798374",
    x"BF79820C",
    x"BF7980A4",
    x"BF797F3C",
    x"BF797DD4",
    x"BF797C6B",
    x"BF797B03",
    x"BF79799A",
    x"BF797831",
    x"BF7976C8",
    x"BF79755F",
    x"BF7973F5",
    x"BF79728C",
    x"BF797122",
    x"BF796FB8",
    x"BF796E4E",
    x"BF796CE4",
    x"BF796B7A",
    x"BF796A0F",
    x"BF7968A5",
    x"BF79673A",
    x"BF7965CF",
    x"BF796464",
    x"BF7962F9",
    x"BF79618E",
    x"BF796022",
    x"BF795EB7",
    x"BF795D4B",
    x"BF795BDF",
    x"BF795A73",
    x"BF795907",
    x"BF79579A",
    x"BF79562E",
    x"BF7954C1",
    x"BF795354",
    x"BF7951E7",
    x"BF79507A",
    x"BF794F0D",
    x"BF794D9F",
    x"BF794C32",
    x"BF794AC4",
    x"BF794956",
    x"BF7947E8",
    x"BF79467A",
    x"BF79450C",
    x"BF79439D",
    x"BF79422F",
    x"BF7940C0",
    x"BF793F51",
    x"BF793DE2",
    x"BF793C73",
    x"BF793B03",
    x"BF793994",
    x"BF793824",
    x"BF7936B4",
    x"BF793544",
    x"BF7933D4",
    x"BF793264",
    x"BF7930F3",
    x"BF792F83",
    x"BF792E12",
    x"BF792CA1",
    x"BF792B30",
    x"BF7929BF",
    x"BF79284E",
    x"BF7926DC",
    x"BF79256B",
    x"BF7923F9",
    x"BF792287",
    x"BF792115",
    x"BF791FA3",
    x"BF791E30",
    x"BF791CBE",
    x"BF791B4B",
    x"BF7919D8",
    x"BF791865",
    x"BF7916F2",
    x"BF79157F",
    x"BF79140B",
    x"BF791298",
    x"BF791124",
    x"BF790FB0",
    x"BF790E3C",
    x"BF790CC8",
    x"BF790B54",
    x"BF7909DF",
    x"BF79086A",
    x"BF7906F6",
    x"BF790581",
    x"BF79040C",
    x"BF790296",
    x"BF790121",
    x"BF78FFAC",
    x"BF78FE36",
    x"BF78FCC0",
    x"BF78FB4A",
    x"BF78F9D4",
    x"BF78F85E",
    x"BF78F6E7",
    x"BF78F571",
    x"BF78F3FA",
    x"BF78F283",
    x"BF78F10C",
    x"BF78EF95",
    x"BF78EE1D",
    x"BF78ECA6",
    x"BF78EB2E",
    x"BF78E9B7",
    x"BF78E83F",
    x"BF78E6C7",
    x"BF78E54E",
    x"BF78E3D6",
    x"BF78E25D",
    x"BF78E0E5",
    x"BF78DF6C",
    x"BF78DDF3",
    x"BF78DC7A",
    x"BF78DB01",
    x"BF78D987",
    x"BF78D80E",
    x"BF78D694",
    x"BF78D51A",
    x"BF78D3A0",
    x"BF78D226",
    x"BF78D0AB",
    x"BF78CF31",
    x"BF78CDB6",
    x"BF78CC3B",
    x"BF78CAC1",
    x"BF78C945",
    x"BF78C7CA",
    x"BF78C64F",
    x"BF78C4D3",
    x"BF78C358",
    x"BF78C1DC",
    x"BF78C060",
    x"BF78BEE4",
    x"BF78BD67",
    x"BF78BBEB",
    x"BF78BA6E",
    x"BF78B8F2",
    x"BF78B775",
    x"BF78B5F8",
    x"BF78B47B",
    x"BF78B2FD",
    x"BF78B180",
    x"BF78B002",
    x"BF78AE84",
    x"BF78AD06",
    x"BF78AB88",
    x"BF78AA0A",
    x"BF78A88C",
    x"BF78A70D",
    x"BF78A58F",
    x"BF78A410",
    x"BF78A291",
    x"BF78A112",
    x"BF789F92",
    x"BF789E13",
    x"BF789C93",
    x"BF789B14",
    x"BF789994",
    x"BF789814",
    x"BF789694",
    x"BF789513",
    x"BF789393",
    x"BF789212",
    x"BF789091",
    x"BF788F11",
    x"BF788D8F",
    x"BF788C0E",
    x"BF788A8D",
    x"BF78890B",
    x"BF78878A",
    x"BF788608",
    x"BF788486",
    x"BF788304",
    x"BF788182",
    x"BF787FFF",
    x"BF787E7D",
    x"BF787CFA",
    x"BF787B77",
    x"BF7879F4",
    x"BF787871",
    x"BF7876ED",
    x"BF78756A",
    x"BF7873E6",
    x"BF787263",
    x"BF7870DF",
    x"BF786F5B",
    x"BF786DD6",
    x"BF786C52",
    x"BF786ACE",
    x"BF786949",
    x"BF7867C4",
    x"BF78663F",
    x"BF7864BA",
    x"BF786335",
    x"BF7861AF",
    x"BF78602A",
    x"BF785EA4",
    x"BF785D1E",
    x"BF785B98",
    x"BF785A12",
    x"BF78588C",
    x"BF785705",
    x"BF78557F",
    x"BF7853F8",
    x"BF785271",
    x"BF7850EA",
    x"BF784F63",
    x"BF784DDB",
    x"BF784C54",
    x"BF784ACC",
    x"BF784944",
    x"BF7847BC",
    x"BF784634",
    x"BF7844AC",
    x"BF784324",
    x"BF78419B",
    x"BF784012",
    x"BF783E8A",
    x"BF783D01",
    x"BF783B77",
    x"BF7839EE",
    x"BF783865",
    x"BF7836DB",
    x"BF783551",
    x"BF7833C7",
    x"BF78323D",
    x"BF7830B3",
    x"BF782F29",
    x"BF782D9E",
    x"BF782C14",
    x"BF782A89",
    x"BF7828FE",
    x"BF782773",
    x"BF7825E8",
    x"BF78245C",
    x"BF7822D1",
    x"BF782145",
    x"BF781FB9",
    x"BF781E2D",
    x"BF781CA1",
    x"BF781B15",
    x"BF781988",
    x"BF7817FC",
    x"BF78166F",
    x"BF7814E2",
    x"BF781355",
    x"BF7811C8",
    x"BF78103A",
    x"BF780EAD",
    x"BF780D1F",
    x"BF780B92",
    x"BF780A04",
    x"BF780876",
    x"BF7806E7",
    x"BF780559",
    x"BF7803CA",
    x"BF78023C",
    x"BF7800AD",
    x"BF77FF1E",
    x"BF77FD8F",
    x"BF77FC00",
    x"BF77FA70",
    x"BF77F8E1",
    x"BF77F751",
    x"BF77F5C1",
    x"BF77F431",
    x"BF77F2A1",
    x"BF77F110",
    x"BF77EF80",
    x"BF77EDEF",
    x"BF77EC5F",
    x"BF77EACE",
    x"BF77E93D",
    x"BF77E7AB",
    x"BF77E61A",
    x"BF77E488",
    x"BF77E2F7",
    x"BF77E165",
    x"BF77DFD3",
    x"BF77DE41",
    x"BF77DCAF",
    x"BF77DB1C",
    x"BF77D98A",
    x"BF77D7F7",
    x"BF77D664",
    x"BF77D4D1",
    x"BF77D33E",
    x"BF77D1AB",
    x"BF77D017",
    x"BF77CE83",
    x"BF77CCF0",
    x"BF77CB5C",
    x"BF77C9C8",
    x"BF77C834",
    x"BF77C69F",
    x"BF77C50B",
    x"BF77C376",
    x"BF77C1E1",
    x"BF77C04C",
    x"BF77BEB7",
    x"BF77BD22",
    x"BF77BB8D",
    x"BF77B9F7",
    x"BF77B861",
    x"BF77B6CB",
    x"BF77B535",
    x"BF77B39F",
    x"BF77B209",
    x"BF77B073",
    x"BF77AEDC",
    x"BF77AD45",
    x"BF77ABAE",
    x"BF77AA17",
    x"BF77A880",
    x"BF77A6E9",
    x"BF77A551",
    x"BF77A3BA",
    x"BF77A222",
    x"BF77A08A",
    x"BF779EF2",
    x"BF779D5A",
    x"BF779BC1",
    x"BF779A29",
    x"BF779890",
    x"BF7796F7",
    x"BF77955E",
    x"BF7793C5",
    x"BF77922C",
    x"BF779092",
    x"BF778EF9",
    x"BF778D5F",
    x"BF778BC5",
    x"BF778A2B",
    x"BF778891",
    x"BF7786F7",
    x"BF77855C",
    x"BF7783C2",
    x"BF778227",
    x"BF77808C",
    x"BF777EF1",
    x"BF777D56",
    x"BF777BBA",
    x"BF777A1F",
    x"BF777883",
    x"BF7776E7",
    x"BF77754B",
    x"BF7773AF",
    x"BF777213",
    x"BF777076",
    x"BF776EDA",
    x"BF776D3D",
    x"BF776BA0",
    x"BF776A03",
    x"BF776866",
    x"BF7766C9",
    x"BF77652B",
    x"BF77638E",
    x"BF7761F0",
    x"BF776052",
    x"BF775EB4",
    x"BF775D16",
    x"BF775B78",
    x"BF7759D9",
    x"BF77583A",
    x"BF77569C",
    x"BF7754FD",
    x"BF77535E",
    x"BF7751BE",
    x"BF77501F",
    x"BF774E7F",
    x"BF774CE0",
    x"BF774B40",
    x"BF7749A0",
    x"BF774800",
    x"BF77465F",
    x"BF7744BF",
    x"BF77431E",
    x"BF77417E",
    x"BF773FDD",
    x"BF773E3C",
    x"BF773C9B",
    x"BF773AF9",
    x"BF773958",
    x"BF7737B6",
    x"BF773614",
    x"BF773472",
    x"BF7732D0",
    x"BF77312E",
    x"BF772F8C",
    x"BF772DE9",
    x"BF772C47",
    x"BF772AA4",
    x"BF772901",
    x"BF77275E",
    x"BF7725BA",
    x"BF772417",
    x"BF772274",
    x"BF7720D0",
    x"BF771F2C",
    x"BF771D88",
    x"BF771BE4",
    x"BF771A3F",
    x"BF77189B",
    x"BF7716F6",
    x"BF771552",
    x"BF7713AD",
    x"BF771208",
    x"BF771063",
    x"BF770EBD",
    x"BF770D18",
    x"BF770B72",
    x"BF7709CC",
    x"BF770826",
    x"BF770680",
    x"BF7704DA",
    x"BF770334",
    x"BF77018D",
    x"BF76FFE6",
    x"BF76FE40",
    x"BF76FC99",
    x"BF76FAF1",
    x"BF76F94A",
    x"BF76F7A3",
    x"BF76F5FB",
    x"BF76F453",
    x"BF76F2AC",
    x"BF76F103",
    x"BF76EF5B",
    x"BF76EDB3",
    x"BF76EC0B",
    x"BF76EA62",
    x"BF76E8B9",
    x"BF76E710",
    x"BF76E567",
    x"BF76E3BE",
    x"BF76E215",
    x"BF76E06B",
    x"BF76DEC1",
    x"BF76DD18",
    x"BF76DB6E",
    x"BF76D9C4",
    x"BF76D819",
    x"BF76D66F",
    x"BF76D4C4",
    x"BF76D31A",
    x"BF76D16F",
    x"BF76CFC4",
    x"BF76CE19",
    x"BF76CC6D",
    x"BF76CAC2",
    x"BF76C916",
    x"BF76C76B",
    x"BF76C5BF",
    x"BF76C413",
    x"BF76C266",
    x"BF76C0BA",
    x"BF76BF0E",
    x"BF76BD61",
    x"BF76BBB4",
    x"BF76BA07",
    x"BF76B85A",
    x"BF76B6AD",
    x"BF76B500",
    x"BF76B352",
    x"BF76B1A4",
    x"BF76AFF7",
    x"BF76AE49",
    x"BF76AC9A",
    x"BF76AAEC",
    x"BF76A93E",
    x"BF76A78F",
    x"BF76A5E0",
    x"BF76A432",
    x"BF76A283",
    x"BF76A0D3",
    x"BF769F24",
    x"BF769D75",
    x"BF769BC5",
    x"BF769A15",
    x"BF769865",
    x"BF7696B5",
    x"BF769505",
    x"BF769355",
    x"BF7691A4",
    x"BF768FF4",
    x"BF768E43",
    x"BF768C92",
    x"BF768AE1",
    x"BF768930",
    x"BF76877E",
    x"BF7685CD",
    x"BF76841B",
    x"BF768269",
    x"BF7680B7",
    x"BF767F05",
    x"BF767D53",
    x"BF767BA0",
    x"BF7679EE",
    x"BF76783B",
    x"BF767688",
    x"BF7674D5",
    x"BF767322",
    x"BF76716F",
    x"BF766FBB",
    x"BF766E08",
    x"BF766C54",
    x"BF766AA0",
    x"BF7668EC",
    x"BF766738",
    x"BF766583",
    x"BF7663CF",
    x"BF76621A",
    x"BF766065",
    x"BF765EB0",
    x"BF765CFB",
    x"BF765B46",
    x"BF765991",
    x"BF7657DB",
    x"BF765625",
    x"BF76546F",
    x"BF7652B9",
    x"BF765103",
    x"BF764F4D",
    x"BF764D97",
    x"BF764BE0",
    x"BF764A29",
    x"BF764872",
    x"BF7646BB",
    x"BF764504",
    x"BF76434D",
    x"BF764195",
    x"BF763FDE",
    x"BF763E26",
    x"BF763C6E",
    x"BF763AB6",
    x"BF7638FE",
    x"BF763745",
    x"BF76358D",
    x"BF7633D4",
    x"BF76321B",
    x"BF763063",
    x"BF762EA9",
    x"BF762CF0",
    x"BF762B37",
    x"BF76297D",
    x"BF7627C3",
    x"BF76260A",
    x"BF762450",
    x"BF762296",
    x"BF7620DB",
    x"BF761F21",
    x"BF761D66",
    x"BF761BAB",
    x"BF7619F1",
    x"BF761836",
    x"BF76167A",
    x"BF7614BF",
    x"BF761304",
    x"BF761148",
    x"BF760F8C",
    x"BF760DD0",
    x"BF760C14",
    x"BF760A58",
    x"BF76089C",
    x"BF7606DF",
    x"BF760522",
    x"BF760366",
    x"BF7601A9",
    x"BF75FFEB",
    x"BF75FE2E",
    x"BF75FC71",
    x"BF75FAB3",
    x"BF75F8F6",
    x"BF75F738",
    x"BF75F57A",
    x"BF75F3BC",
    x"BF75F1FD",
    x"BF75F03F",
    x"BF75EE80",
    x"BF75ECC2",
    x"BF75EB03",
    x"BF75E944",
    x"BF75E784",
    x"BF75E5C5",
    x"BF75E406",
    x"BF75E246",
    x"BF75E086",
    x"BF75DEC6",
    x"BF75DD06",
    x"BF75DB46",
    x"BF75D986",
    x"BF75D7C5",
    x"BF75D604",
    x"BF75D444",
    x"BF75D283",
    x"BF75D0C2",
    x"BF75CF00",
    x"BF75CD3F",
    x"BF75CB7D",
    x"BF75C9BC",
    x"BF75C7FA",
    x"BF75C638",
    x"BF75C476",
    x"BF75C2B3",
    x"BF75C0F1",
    x"BF75BF2E",
    x"BF75BD6C",
    x"BF75BBA9",
    x"BF75B9E6",
    x"BF75B822",
    x"BF75B65F",
    x"BF75B49C",
    x"BF75B2D8",
    x"BF75B114",
    x"BF75AF50",
    x"BF75AD8C",
    x"BF75ABC8",
    x"BF75AA04",
    x"BF75A83F",
    x"BF75A67B",
    x"BF75A4B6",
    x"BF75A2F1",
    x"BF75A12C",
    x"BF759F66",
    x"BF759DA1",
    x"BF759BDB",
    x"BF759A16",
    x"BF759850",
    x"BF75968A",
    x"BF7594C4",
    x"BF7592FE",
    x"BF759137",
    x"BF758F70",
    x"BF758DAA",
    x"BF758BE3",
    x"BF758A1C",
    x"BF758855",
    x"BF75868D",
    x"BF7584C6",
    x"BF7582FE",
    x"BF758136",
    x"BF757F6F",
    x"BF757DA7",
    x"BF757BDE",
    x"BF757A16",
    x"BF75784D",
    x"BF757685",
    x"BF7574BC",
    x"BF7572F3",
    x"BF75712A",
    x"BF756F61",
    x"BF756D97",
    x"BF756BCE",
    x"BF756A04",
    x"BF75683A",
    x"BF756670",
    x"BF7564A6",
    x"BF7562DC",
    x"BF756111",
    x"BF755F47",
    x"BF755D7C",
    x"BF755BB1",
    x"BF7559E6",
    x"BF75581B",
    x"BF755650",
    x"BF755484",
    x"BF7552B9",
    x"BF7550ED",
    x"BF754F21",
    x"BF754D55",
    x"BF754B89",
    x"BF7549BC",
    x"BF7547F0",
    x"BF754623",
    x"BF754456",
    x"BF754289",
    x"BF7540BC",
    x"BF753EEF",
    x"BF753D22",
    x"BF753B54",
    x"BF753987",
    x"BF7537B9",
    x"BF7535EB",
    x"BF75341D",
    x"BF75324E",
    x"BF753080",
    x"BF752EB1",
    x"BF752CE3",
    x"BF752B14",
    x"BF752945",
    x"BF752776",
    x"BF7525A6",
    x"BF7523D7",
    x"BF752207",
    x"BF752038",
    x"BF751E68",
    x"BF751C98",
    x"BF751AC7",
    x"BF7518F7",
    x"BF751727",
    x"BF751556",
    x"BF751385",
    x"BF7511B4",
    x"BF750FE3",
    x"BF750E12",
    x"BF750C41",
    x"BF750A6F",
    x"BF75089D",
    x"BF7506CC",
    x"BF7504FA",
    x"BF750327",
    x"BF750155",
    x"BF74FF83",
    x"BF74FDB0",
    x"BF74FBDE",
    x"BF74FA0B",
    x"BF74F838",
    x"BF74F665",
    x"BF74F491",
    x"BF74F2BE",
    x"BF74F0EA",
    x"BF74EF17",
    x"BF74ED43",
    x"BF74EB6F",
    x"BF74E99A",
    x"BF74E7C6",
    x"BF74E5F2",
    x"BF74E41D",
    x"BF74E248",
    x"BF74E073",
    x"BF74DE9E",
    x"BF74DCC9",
    x"BF74DAF4",
    x"BF74D91E",
    x"BF74D749",
    x"BF74D573",
    x"BF74D39D",
    x"BF74D1C7",
    x"BF74CFF0",
    x"BF74CE1A",
    x"BF74CC44",
    x"BF74CA6D",
    x"BF74C896",
    x"BF74C6BF",
    x"BF74C4E8",
    x"BF74C311",
    x"BF74C139",
    x"BF74BF62",
    x"BF74BD8A",
    x"BF74BBB2",
    x"BF74B9DA",
    x"BF74B802",
    x"BF74B62A",
    x"BF74B451",
    x"BF74B279",
    x"BF74B0A0",
    x"BF74AEC7",
    x"BF74ACEE",
    x"BF74AB15",
    x"BF74A93B",
    x"BF74A762",
    x"BF74A588",
    x"BF74A3AE",
    x"BF74A1D5",
    x"BF749FFA",
    x"BF749E20",
    x"BF749C46",
    x"BF749A6B",
    x"BF749891",
    x"BF7496B6",
    x"BF7494DB",
    x"BF749300",
    x"BF749125",
    x"BF748F49",
    x"BF748D6E",
    x"BF748B92",
    x"BF7489B6",
    x"BF7487DA",
    x"BF7485FE",
    x"BF748422",
    x"BF748245",
    x"BF748069",
    x"BF747E8C",
    x"BF747CAF",
    x"BF747AD2",
    x"BF7478F5",
    x"BF747718",
    x"BF74753A",
    x"BF74735D",
    x"BF74717F",
    x"BF746FA1",
    x"BF746DC3",
    x"BF746BE5",
    x"BF746A06",
    x"BF746828",
    x"BF746649",
    x"BF74646A",
    x"BF74628B",
    x"BF7460AC",
    x"BF745ECD",
    x"BF745CEE",
    x"BF745B0E",
    x"BF74592F",
    x"BF74574F",
    x"BF74556F",
    x"BF74538F",
    x"BF7451AE",
    x"BF744FCE",
    x"BF744DED",
    x"BF744C0D",
    x"BF744A2C",
    x"BF74484B",
    x"BF74466A",
    x"BF744488",
    x"BF7442A7",
    x"BF7440C5",
    x"BF743EE4",
    x"BF743D02",
    x"BF743B20",
    x"BF74393E",
    x"BF74375B",
    x"BF743579",
    x"BF743396",
    x"BF7431B3",
    x"BF742FD1",
    x"BF742DED",
    x"BF742C0A",
    x"BF742A27",
    x"BF742843",
    x"BF742660",
    x"BF74247C",
    x"BF742298",
    x"BF7420B4",
    x"BF741ED0",
    x"BF741CEB",
    x"BF741B07",
    x"BF741922",
    x"BF74173D",
    x"BF741558",
    x"BF741373",
    x"BF74118E",
    x"BF740FA9",
    x"BF740DC3",
    x"BF740BDD",
    x"BF7409F8",
    x"BF740812",
    x"BF74062B",
    x"BF740445",
    x"BF74025F",
    x"BF740078",
    x"BF73FE91",
    x"BF73FCAA",
    x"BF73FAC3",
    x"BF73F8DC",
    x"BF73F6F5",
    x"BF73F50D",
    x"BF73F326",
    x"BF73F13E",
    x"BF73EF56",
    x"BF73ED6E",
    x"BF73EB86",
    x"BF73E99E",
    x"BF73E7B5",
    x"BF73E5CC",
    x"BF73E3E4",
    x"BF73E1FB",
    x"BF73E012",
    x"BF73DE28",
    x"BF73DC3F",
    x"BF73DA56",
    x"BF73D86C",
    x"BF73D682",
    x"BF73D498",
    x"BF73D2AE",
    x"BF73D0C4",
    x"BF73CED9",
    x"BF73CCEF",
    x"BF73CB04",
    x"BF73C919",
    x"BF73C72E",
    x"BF73C543",
    x"BF73C358",
    x"BF73C16C",
    x"BF73BF81",
    x"BF73BD95",
    x"BF73BBA9",
    x"BF73B9BD",
    x"BF73B7D1",
    x"BF73B5E5",
    x"BF73B3F8",
    x"BF73B20C",
    x"BF73B01F",
    x"BF73AE32",
    x"BF73AC45",
    x"BF73AA58",
    x"BF73A86A",
    x"BF73A67D",
    x"BF73A48F",
    x"BF73A2A1",
    x"BF73A0B4",
    x"BF739EC5",
    x"BF739CD7",
    x"BF739AE9",
    x"BF7398FA",
    x"BF73970C",
    x"BF73951D",
    x"BF73932E",
    x"BF73913F",
    x"BF738F50",
    x"BF738D60",
    x"BF738B71",
    x"BF738981",
    x"BF738791",
    x"BF7385A1",
    x"BF7383B1",
    x"BF7381C1",
    x"BF737FD0",
    x"BF737DE0",
    x"BF737BEF",
    x"BF7379FE",
    x"BF73780D",
    x"BF73761C",
    x"BF73742B",
    x"BF737239",
    x"BF737048",
    x"BF736E56",
    x"BF736C64",
    x"BF736A72",
    x"BF736880",
    x"BF73668E",
    x"BF73649B",
    x"BF7362A8",
    x"BF7360B6",
    x"BF735EC3",
    x"BF735CD0",
    x"BF735ADC",
    x"BF7358E9",
    x"BF7356F6",
    x"BF735502",
    x"BF73530E",
    x"BF73511A",
    x"BF734F26",
    x"BF734D32",
    x"BF734B3E",
    x"BF734949",
    x"BF734754",
    x"BF734560",
    x"BF73436B",
    x"BF734175",
    x"BF733F80",
    x"BF733D8B",
    x"BF733B95",
    x"BF7339A0",
    x"BF7337AA",
    x"BF7335B4",
    x"BF7333BE",
    x"BF7331C7",
    x"BF732FD1",
    x"BF732DDA",
    x"BF732BE4",
    x"BF7329ED",
    x"BF7327F6",
    x"BF7325FE",
    x"BF732407",
    x"BF732210",
    x"BF732018",
    x"BF731E20",
    x"BF731C28",
    x"BF731A30",
    x"BF731838",
    x"BF731640",
    x"BF731447",
    x"BF73124F",
    x"BF731056",
    x"BF730E5D",
    x"BF730C64",
    x"BF730A6B",
    x"BF730871",
    x"BF730678",
    x"BF73047E",
    x"BF730284",
    x"BF73008B",
    x"BF72FE90",
    x"BF72FC96",
    x"BF72FA9C",
    x"BF72F8A1",
    x"BF72F6A7",
    x"BF72F4AC",
    x"BF72F2B1",
    x"BF72F0B6",
    x"BF72EEBA",
    x"BF72ECBF",
    x"BF72EAC3",
    x"BF72E8C8",
    x"BF72E6CC",
    x"BF72E4D0",
    x"BF72E2D4",
    x"BF72E0D7",
    x"BF72DEDB",
    x"BF72DCDE",
    x"BF72DAE2",
    x"BF72D8E5",
    x"BF72D6E8",
    x"BF72D4EB",
    x"BF72D2ED",
    x"BF72D0F0",
    x"BF72CEF2",
    x"BF72CCF5",
    x"BF72CAF7",
    x"BF72C8F9",
    x"BF72C6FA",
    x"BF72C4FC",
    x"BF72C2FE",
    x"BF72C0FF",
    x"BF72BF00",
    x"BF72BD01",
    x"BF72BB02",
    x"BF72B903",
    x"BF72B704",
    x"BF72B504",
    x"BF72B304",
    x"BF72B105",
    x"BF72AF05",
    x"BF72AD05",
    x"BF72AB04",
    x"BF72A904",
    x"BF72A703",
    x"BF72A503",
    x"BF72A302",
    x"BF72A101",
    x"BF729F00",
    x"BF729CFF",
    x"BF729AFD",
    x"BF7298FC",
    x"BF7296FA",
    x"BF7294F8",
    x"BF7292F6",
    x"BF7290F4",
    x"BF728EF2",
    x"BF728CEF",
    x"BF728AED",
    x"BF7288EA",
    x"BF7286E7",
    x"BF7284E4",
    x"BF7282E1",
    x"BF7280DE",
    x"BF727EDA",
    x"BF727CD7",
    x"BF727AD3",
    x"BF7278CF",
    x"BF7276CB",
    x"BF7274C7",
    x"BF7272C2",
    x"BF7270BE",
    x"BF726EB9",
    x"BF726CB5",
    x"BF726AB0",
    x"BF7268AB",
    x"BF7266A5",
    x"BF7264A0",
    x"BF72629B",
    x"BF726095",
    x"BF725E8F",
    x"BF725C89",
    x"BF725A83",
    x"BF72587D",
    x"BF725677",
    x"BF725470",
    x"BF725269",
    x"BF725063",
    x"BF724E5C",
    x"BF724C54",
    x"BF724A4D",
    x"BF724846",
    x"BF72463E",
    x"BF724437",
    x"BF72422F",
    x"BF724027",
    x"BF723E1F",
    x"BF723C16",
    x"BF723A0E",
    x"BF723805",
    x"BF7235FD",
    x"BF7233F4",
    x"BF7231EB",
    x"BF722FE2",
    x"BF722DD8",
    x"BF722BCF",
    x"BF7229C5",
    x"BF7227BC",
    x"BF7225B2",
    x"BF7223A8",
    x"BF72219E",
    x"BF721F93",
    x"BF721D89",
    x"BF721B7E",
    x"BF721973",
    x"BF721769",
    x"BF72155E",
    x"BF721352",
    x"BF721147",
    x"BF720F3C",
    x"BF720D30",
    x"BF720B24",
    x"BF720918",
    x"BF72070C",
    x"BF720500",
    x"BF7202F4",
    x"BF7200E7",
    x"BF71FEDA",
    x"BF71FCCE",
    x"BF71FAC1",
    x"BF71F8B4",
    x"BF71F6A6",
    x"BF71F499",
    x"BF71F28C",
    x"BF71F07E",
    x"BF71EE70",
    x"BF71EC62",
    x"BF71EA54",
    x"BF71E846",
    x"BF71E637",
    x"BF71E429",
    x"BF71E21A",
    x"BF71E00B",
    x"BF71DDFC",
    x"BF71DBED",
    x"BF71D9DE",
    x"BF71D7CF",
    x"BF71D5BF",
    x"BF71D3AF",
    x"BF71D19F",
    x"BF71CF8F",
    x"BF71CD7F",
    x"BF71CB6F",
    x"BF71C95F",
    x"BF71C74E",
    x"BF71C53D",
    x"BF71C32C",
    x"BF71C11B",
    x"BF71BF0A",
    x"BF71BCF9",
    x"BF71BAE7",
    x"BF71B8D6",
    x"BF71B6C4",
    x"BF71B4B2",
    x"BF71B2A0",
    x"BF71B08E",
    x"BF71AE7C",
    x"BF71AC69",
    x"BF71AA57",
    x"BF71A844",
    x"BF71A631",
    x"BF71A41E",
    x"BF71A20B",
    x"BF719FF7",
    x"BF719DE4",
    x"BF719BD0",
    x"BF7199BC",
    x"BF7197A8",
    x"BF719594",
    x"BF719380",
    x"BF71916C",
    x"BF718F57",
    x"BF718D43",
    x"BF718B2E",
    x"BF718919",
    x"BF718704",
    x"BF7184EF",
    x"BF7182D9",
    x"BF7180C4",
    x"BF717EAE",
    x"BF717C98",
    x"BF717A82",
    x"BF71786C",
    x"BF717656",
    x"BF71743F",
    x"BF717229",
    x"BF717012",
    x"BF716DFB",
    x"BF716BE4",
    x"BF7169CD",
    x"BF7167B6",
    x"BF71659F",
    x"BF716387",
    x"BF71616F",
    x"BF715F57",
    x"BF715D3F",
    x"BF715B27",
    x"BF71590F",
    x"BF7156F6",
    x"BF7154DE",
    x"BF7152C5",
    x"BF7150AC",
    x"BF714E93",
    x"BF714C7A",
    x"BF714A61",
    x"BF714847",
    x"BF71462E",
    x"BF714414",
    x"BF7141FA",
    x"BF713FE0",
    x"BF713DC6",
    x"BF713BAC",
    x"BF713991",
    x"BF713776",
    x"BF71355C",
    x"BF713341",
    x"BF713126",
    x"BF712F0B",
    x"BF712CEF",
    x"BF712AD4",
    x"BF7128B8",
    x"BF71269C",
    x"BF712480",
    x"BF712264",
    x"BF712048",
    x"BF711E2C",
    x"BF711C0F",
    x"BF7119F3",
    x"BF7117D6",
    x"BF7115B9",
    x"BF71139C",
    x"BF71117F",
    x"BF710F61",
    x"BF710D44",
    x"BF710B26",
    x"BF710908",
    x"BF7106EA",
    x"BF7104CC",
    x"BF7102AE",
    x"BF71008F",
    x"BF70FE71",
    x"BF70FC52",
    x"BF70FA33",
    x"BF70F814",
    x"BF70F5F5",
    x"BF70F3D6",
    x"BF70F1B7",
    x"BF70EF97",
    x"BF70ED77",
    x"BF70EB58",
    x"BF70E938",
    x"BF70E717",
    x"BF70E4F7",
    x"BF70E2D7",
    x"BF70E0B6",
    x"BF70DE95",
    x"BF70DC75",
    x"BF70DA54",
    x"BF70D832",
    x"BF70D611",
    x"BF70D3F0",
    x"BF70D1CE",
    x"BF70CFAC",
    x"BF70CD8A",
    x"BF70CB68",
    x"BF70C946",
    x"BF70C724",
    x"BF70C501",
    x"BF70C2DF",
    x"BF70C0BC",
    x"BF70BE99",
    x"BF70BC76",
    x"BF70BA53",
    x"BF70B830",
    x"BF70B60C",
    x"BF70B3E9",
    x"BF70B1C5",
    x"BF70AFA1",
    x"BF70AD7D",
    x"BF70AB59",
    x"BF70A934",
    x"BF70A710",
    x"BF70A4EB",
    x"BF70A2C6",
    x"BF70A0A2",
    x"BF709E7C",
    x"BF709C57",
    x"BF709A32",
    x"BF70980C",
    x"BF7095E7",
    x"BF7093C1",
    x"BF70919B",
    x"BF708F75",
    x"BF708D4F",
    x"BF708B28",
    x"BF708902",
    x"BF7086DB",
    x"BF7084B4",
    x"BF70828D",
    x"BF708066",
    x"BF707E3F",
    x"BF707C18",
    x"BF7079F0",
    x"BF7077C8",
    x"BF7075A1",
    x"BF707379",
    x"BF707151",
    x"BF706F28",
    x"BF706D00",
    x"BF706AD7",
    x"BF7068AF",
    x"BF706686",
    x"BF70645D",
    x"BF706234",
    x"BF70600A",
    x"BF705DE1",
    x"BF705BB8",
    x"BF70598E",
    x"BF705764",
    x"BF70553A",
    x"BF705310",
    x"BF7050E6",
    x"BF704EBB",
    x"BF704C91",
    x"BF704A66",
    x"BF70483B",
    x"BF704610",
    x"BF7043E5",
    x"BF7041BA",
    x"BF703F8E",
    x"BF703D63",
    x"BF703B37",
    x"BF70390B",
    x"BF7036DF",
    x"BF7034B3",
    x"BF703286",
    x"BF70305A",
    x"BF702E2D",
    x"BF702C01",
    x"BF7029D4",
    x"BF7027A7",
    x"BF70257A",
    x"BF70234C",
    x"BF70211F",
    x"BF701EF1",
    x"BF701CC3",
    x"BF701A95",
    x"BF701867",
    x"BF701639",
    x"BF70140B",
    x"BF7011DC",
    x"BF700FAE",
    x"BF700D7F",
    x"BF700B50",
    x"BF700921",
    x"BF7006F2",
    x"BF7004C3",
    x"BF700293",
    x"BF700063",
    x"BF6FFE34",
    x"BF6FFC04",
    x"BF6FF9D4",
    x"BF6FF7A3",
    x"BF6FF573",
    x"BF6FF343",
    x"BF6FF112",
    x"BF6FEEE1",
    x"BF6FECB0",
    x"BF6FEA7F",
    x"BF6FE84E",
    x"BF6FE61D",
    x"BF6FE3EB",
    x"BF6FE1B9",
    x"BF6FDF88",
    x"BF6FDD56",
    x"BF6FDB24",
    x"BF6FD8F1",
    x"BF6FD6BF",
    x"BF6FD48C",
    x"BF6FD25A",
    x"BF6FD027",
    x"BF6FCDF4",
    x"BF6FCBC1",
    x"BF6FC98E",
    x"BF6FC75A",
    x"BF6FC527",
    x"BF6FC2F3",
    x"BF6FC0BF",
    x"BF6FBE8B",
    x"BF6FBC57",
    x"BF6FBA23",
    x"BF6FB7EE",
    x"BF6FB5BA",
    x"BF6FB385",
    x"BF6FB150",
    x"BF6FAF1B",
    x"BF6FACE6",
    x"BF6FAAB1",
    x"BF6FA87C",
    x"BF6FA646",
    x"BF6FA410",
    x"BF6FA1DA",
    x"BF6F9FA4",
    x"BF6F9D6E",
    x"BF6F9B38",
    x"BF6F9902",
    x"BF6F96CB",
    x"BF6F9494",
    x"BF6F925D",
    x"BF6F9026",
    x"BF6F8DEF",
    x"BF6F8BB8",
    x"BF6F8981",
    x"BF6F8749",
    x"BF6F8511",
    x"BF6F82D9",
    x"BF6F80A1",
    x"BF6F7E69",
    x"BF6F7C31",
    x"BF6F79F8",
    x"BF6F77C0",
    x"BF6F7587",
    x"BF6F734E",
    x"BF6F7115",
    x"BF6F6EDC",
    x"BF6F6CA3",
    x"BF6F6A69",
    x"BF6F6830",
    x"BF6F65F6",
    x"BF6F63BC",
    x"BF6F6182",
    x"BF6F5F48",
    x"BF6F5D0E",
    x"BF6F5AD3",
    x"BF6F5899",
    x"BF6F565E",
    x"BF6F5423",
    x"BF6F51E8",
    x"BF6F4FAD",
    x"BF6F4D71",
    x"BF6F4B36",
    x"BF6F48FA",
    x"BF6F46BE",
    x"BF6F4483",
    x"BF6F4247",
    x"BF6F400A",
    x"BF6F3DCE",
    x"BF6F3B92",
    x"BF6F3955",
    x"BF6F3718",
    x"BF6F34DB",
    x"BF6F329E",
    x"BF6F3061",
    x"BF6F2E24",
    x"BF6F2BE6",
    x"BF6F29A8",
    x"BF6F276B",
    x"BF6F252D",
    x"BF6F22EF",
    x"BF6F20B0",
    x"BF6F1E72",
    x"BF6F1C34",
    x"BF6F19F5",
    x"BF6F17B6",
    x"BF6F1577",
    x"BF6F1338",
    x"BF6F10F9",
    x"BF6F0EBA",
    x"BF6F0C7A",
    x"BF6F0A3A",
    x"BF6F07FB",
    x"BF6F05BB",
    x"BF6F037B",
    x"BF6F013A",
    x"BF6EFEFA",
    x"BF6EFCBA",
    x"BF6EFA79",
    x"BF6EF838",
    x"BF6EF5F7",
    x"BF6EF3B6",
    x"BF6EF175",
    x"BF6EEF33",
    x"BF6EECF2",
    x"BF6EEAB0",
    x"BF6EE86E",
    x"BF6EE62C",
    x"BF6EE3EA",
    x"BF6EE1A8",
    x"BF6EDF66",
    x"BF6EDD23",
    x"BF6EDAE1",
    x"BF6ED89E",
    x"BF6ED65B",
    x"BF6ED418",
    x"BF6ED1D4",
    x"BF6ECF91",
    x"BF6ECD4D",
    x"BF6ECB0A",
    x"BF6EC8C6",
    x"BF6EC682",
    x"BF6EC43E",
    x"BF6EC1FA",
    x"BF6EBFB5",
    x"BF6EBD71",
    x"BF6EBB2C",
    x"BF6EB8E7",
    x"BF6EB6A2",
    x"BF6EB45D",
    x"BF6EB218",
    x"BF6EAFD2",
    x"BF6EAD8D",
    x"BF6EAB47",
    x"BF6EA901",
    x"BF6EA6BB",
    x"BF6EA475",
    x"BF6EA22F",
    x"BF6E9FE9",
    x"BF6E9DA2",
    x"BF6E9B5B",
    x"BF6E9914",
    x"BF6E96CD",
    x"BF6E9486",
    x"BF6E923F",
    x"BF6E8FF8",
    x"BF6E8DB0",
    x"BF6E8B68",
    x"BF6E8920",
    x"BF6E86D8",
    x"BF6E8490",
    x"BF6E8248",
    x"BF6E8000",
    x"BF6E7DB7",
    x"BF6E7B6E",
    x"BF6E7926",
    x"BF6E76DD",
    x"BF6E7493",
    x"BF6E724A",
    x"BF6E7001",
    x"BF6E6DB7",
    x"BF6E6B6D",
    x"BF6E6924",
    x"BF6E66D9",
    x"BF6E648F",
    x"BF6E6245",
    x"BF6E5FFB",
    x"BF6E5DB0",
    x"BF6E5B65",
    x"BF6E591A",
    x"BF6E56CF",
    x"BF6E5484",
    x"BF6E5239",
    x"BF6E4FEE",
    x"BF6E4DA2",
    x"BF6E4B56",
    x"BF6E490A",
    x"BF6E46BE",
    x"BF6E4472",
    x"BF6E4226",
    x"BF6E3FD9",
    x"BF6E3D8D",
    x"BF6E3B40",
    x"BF6E38F3",
    x"BF6E36A6",
    x"BF6E3459",
    x"BF6E320C",
    x"BF6E2FBE",
    x"BF6E2D71",
    x"BF6E2B23",
    x"BF6E28D5",
    x"BF6E2687",
    x"BF6E2439",
    x"BF6E21EB",
    x"BF6E1F9C",
    x"BF6E1D4E",
    x"BF6E1AFF",
    x"BF6E18B0",
    x"BF6E1661",
    x"BF6E1412",
    x"BF6E11C2",
    x"BF6E0F73",
    x"BF6E0D23",
    x"BF6E0AD4",
    x"BF6E0884",
    x"BF6E0634",
    x"BF6E03E3",
    x"BF6E0193",
    x"BF6DFF43",
    x"BF6DFCF2",
    x"BF6DFAA1",
    x"BF6DF850",
    x"BF6DF5FF",
    x"BF6DF3AE",
    x"BF6DF15D",
    x"BF6DEF0B",
    x"BF6DECBA",
    x"BF6DEA68",
    x"BF6DE816",
    x"BF6DE5C4",
    x"BF6DE372",
    x"BF6DE120",
    x"BF6DDECD",
    x"BF6DDC7B",
    x"BF6DDA28",
    x"BF6DD7D5",
    x"BF6DD582",
    x"BF6DD32F",
    x"BF6DD0DB",
    x"BF6DCE88",
    x"BF6DCC34",
    x"BF6DC9E1",
    x"BF6DC78D",
    x"BF6DC539",
    x"BF6DC2E4",
    x"BF6DC090",
    x"BF6DBE3C",
    x"BF6DBBE7",
    x"BF6DB992",
    x"BF6DB73D",
    x"BF6DB4E8",
    x"BF6DB293",
    x"BF6DB03E",
    x"BF6DADE8",
    x"BF6DAB93",
    x"BF6DA93D",
    x"BF6DA6E7",
    x"BF6DA491",
    x"BF6DA23B",
    x"BF6D9FE4",
    x"BF6D9D8E",
    x"BF6D9B37",
    x"BF6D98E1",
    x"BF6D968A",
    x"BF6D9433",
    x"BF6D91DB",
    x"BF6D8F84",
    x"BF6D8D2D",
    x"BF6D8AD5",
    x"BF6D887D",
    x"BF6D8625",
    x"BF6D83CD",
    x"BF6D8175",
    x"BF6D7F1D",
    x"BF6D7CC4",
    x"BF6D7A6C",
    x"BF6D7813",
    x"BF6D75BA",
    x"BF6D7361",
    x"BF6D7108",
    x"BF6D6EAE",
    x"BF6D6C55",
    x"BF6D69FB",
    x"BF6D67A1",
    x"BF6D6547",
    x"BF6D62ED",
    x"BF6D6093",
    x"BF6D5E39",
    x"BF6D5BDE",
    x"BF6D5984",
    x"BF6D5729",
    x"BF6D54CE",
    x"BF6D5273",
    x"BF6D5018",
    x"BF6D4DBC",
    x"BF6D4B61",
    x"BF6D4905",
    x"BF6D46AA",
    x"BF6D444E",
    x"BF6D41F2",
    x"BF6D3F95",
    x"BF6D3D39",
    x"BF6D3ADD",
    x"BF6D3880",
    x"BF6D3623",
    x"BF6D33C6",
    x"BF6D3169",
    x"BF6D2F0C",
    x"BF6D2CAF",
    x"BF6D2A51",
    x"BF6D27F4",
    x"BF6D2596",
    x"BF6D2338",
    x"BF6D20DA",
    x"BF6D1E7C",
    x"BF6D1C1D",
    x"BF6D19BF",
    x"BF6D1760",
    x"BF6D1501",
    x"BF6D12A2",
    x"BF6D1043",
    x"BF6D0DE4",
    x"BF6D0B85",
    x"BF6D0925",
    x"BF6D06C6",
    x"BF6D0466",
    x"BF6D0206",
    x"BF6CFFA6",
    x"BF6CFD46",
    x"BF6CFAE5",
    x"BF6CF885",
    x"BF6CF624",
    x"BF6CF3C4",
    x"BF6CF163",
    x"BF6CEF02",
    x"BF6CECA0",
    x"BF6CEA3F",
    x"BF6CE7DE",
    x"BF6CE57C",
    x"BF6CE31A",
    x"BF6CE0B8",
    x"BF6CDE56",
    x"BF6CDBF4",
    x"BF6CD992",
    x"BF6CD72F",
    x"BF6CD4CD",
    x"BF6CD26A",
    x"BF6CD007",
    x"BF6CCDA4",
    x"BF6CCB41",
    x"BF6CC8DD",
    x"BF6CC67A",
    x"BF6CC416",
    x"BF6CC1B2",
    x"BF6CBF4F",
    x"BF6CBCEA",
    x"BF6CBA86",
    x"BF6CB822",
    x"BF6CB5BD",
    x"BF6CB359",
    x"BF6CB0F4",
    x"BF6CAE8F",
    x"BF6CAC2A",
    x"BF6CA9C5",
    x"BF6CA760",
    x"BF6CA4FA",
    x"BF6CA295",
    x"BF6CA02F",
    x"BF6C9DC9",
    x"BF6C9B63",
    x"BF6C98FD",
    x"BF6C9696",
    x"BF6C9430",
    x"BF6C91C9",
    x"BF6C8F62",
    x"BF6C8CFC",
    x"BF6C8A94",
    x"BF6C882D",
    x"BF6C85C6",
    x"BF6C835E",
    x"BF6C80F7",
    x"BF6C7E8F",
    x"BF6C7C27",
    x"BF6C79BF",
    x"BF6C7757",
    x"BF6C74EF",
    x"BF6C7286",
    x"BF6C701E",
    x"BF6C6DB5",
    x"BF6C6B4C",
    x"BF6C68E3",
    x"BF6C667A",
    x"BF6C6410",
    x"BF6C61A7",
    x"BF6C5F3D",
    x"BF6C5CD4",
    x"BF6C5A6A",
    x"BF6C5800",
    x"BF6C5595",
    x"BF6C532B",
    x"BF6C50C1",
    x"BF6C4E56",
    x"BF6C4BEB",
    x"BF6C4980",
    x"BF6C4715",
    x"BF6C44AA",
    x"BF6C423F",
    x"BF6C3FD3",
    x"BF6C3D68",
    x"BF6C3AFC",
    x"BF6C3890",
    x"BF6C3624",
    x"BF6C33B8",
    x"BF6C314C",
    x"BF6C2EDF",
    x"BF6C2C73",
    x"BF6C2A06",
    x"BF6C2799",
    x"BF6C252C",
    x"BF6C22BF",
    x"BF6C2051",
    x"BF6C1DE4",
    x"BF6C1B76",
    x"BF6C1909",
    x"BF6C169B",
    x"BF6C142D",
    x"BF6C11BF",
    x"BF6C0F50",
    x"BF6C0CE2",
    x"BF6C0A73",
    x"BF6C0805",
    x"BF6C0596",
    x"BF6C0327",
    x"BF6C00B7",
    x"BF6BFE48",
    x"BF6BFBD9",
    x"BF6BF969",
    x"BF6BF6F9",
    x"BF6BF48A",
    x"BF6BF21A",
    x"BF6BEFA9",
    x"BF6BED39",
    x"BF6BEAC9",
    x"BF6BE858",
    x"BF6BE5E7",
    x"BF6BE376",
    x"BF6BE105",
    x"BF6BDE94",
    x"BF6BDC23",
    x"BF6BD9B2",
    x"BF6BD740",
    x"BF6BD4CE",
    x"BF6BD25C",
    x"BF6BCFEA",
    x"BF6BCD78",
    x"BF6BCB06",
    x"BF6BC894",
    x"BF6BC621",
    x"BF6BC3AE",
    x"BF6BC13B",
    x"BF6BBEC8",
    x"BF6BBC55",
    x"BF6BB9E2",
    x"BF6BB76F",
    x"BF6BB4FB",
    x"BF6BB287",
    x"BF6BB014",
    x"BF6BADA0",
    x"BF6BAB2B",
    x"BF6BA8B7",
    x"BF6BA643",
    x"BF6BA3CE",
    x"BF6BA159",
    x"BF6B9EE5",
    x"BF6B9C70",
    x"BF6B99FB",
    x"BF6B9785",
    x"BF6B9510",
    x"BF6B929A",
    x"BF6B9025",
    x"BF6B8DAF",
    x"BF6B8B39",
    x"BF6B88C3",
    x"BF6B864C",
    x"BF6B83D6",
    x"BF6B815F",
    x"BF6B7EE9",
    x"BF6B7C72",
    x"BF6B79FB",
    x"BF6B7784",
    x"BF6B750D",
    x"BF6B7295",
    x"BF6B701E",
    x"BF6B6DA6",
    x"BF6B6B2E",
    x"BF6B68B6",
    x"BF6B663E",
    x"BF6B63C6",
    x"BF6B614D",
    x"BF6B5ED5",
    x"BF6B5C5C",
    x"BF6B59E3",
    x"BF6B576B",
    x"BF6B54F1",
    x"BF6B5278",
    x"BF6B4FFF",
    x"BF6B4D85",
    x"BF6B4B0C",
    x"BF6B4892",
    x"BF6B4618",
    x"BF6B439E",
    x"BF6B4124",
    x"BF6B3EA9",
    x"BF6B3C2F",
    x"BF6B39B4",
    x"BF6B3739",
    x"BF6B34BE",
    x"BF6B3243",
    x"BF6B2FC8",
    x"BF6B2D4D",
    x"BF6B2AD1",
    x"BF6B2855",
    x"BF6B25DA",
    x"BF6B235E",
    x"BF6B20E2",
    x"BF6B1E65",
    x"BF6B1BE9",
    x"BF6B196D",
    x"BF6B16F0",
    x"BF6B1473",
    x"BF6B11F6",
    x"BF6B0F79",
    x"BF6B0CFC",
    x"BF6B0A7F",
    x"BF6B0801",
    x"BF6B0584",
    x"BF6B0306",
    x"BF6B0088",
    x"BF6AFE0A",
    x"BF6AFB8C",
    x"BF6AF90D",
    x"BF6AF68F",
    x"BF6AF410",
    x"BF6AF191",
    x"BF6AEF12",
    x"BF6AEC93",
    x"BF6AEA14",
    x"BF6AE795",
    x"BF6AE515",
    x"BF6AE296",
    x"BF6AE016",
    x"BF6ADD96",
    x"BF6ADB16",
    x"BF6AD896",
    x"BF6AD616",
    x"BF6AD395",
    x"BF6AD115",
    x"BF6ACE94",
    x"BF6ACC13",
    x"BF6AC992",
    x"BF6AC711",
    x"BF6AC48F",
    x"BF6AC20E",
    x"BF6ABF8C",
    x"BF6ABD0B",
    x"BF6ABA89",
    x"BF6AB807",
    x"BF6AB585",
    x"BF6AB302",
    x"BF6AB080",
    x"BF6AADFD",
    x"BF6AAB7B",
    x"BF6AA8F8",
    x"BF6AA675",
    x"BF6AA3F2",
    x"BF6AA16E",
    x"BF6A9EEB",
    x"BF6A9C67",
    x"BF6A99E4",
    x"BF6A9760",
    x"BF6A94DC",
    x"BF6A9258",
    x"BF6A8FD3",
    x"BF6A8D4F",
    x"BF6A8ACA",
    x"BF6A8846",
    x"BF6A85C1",
    x"BF6A833C",
    x"BF6A80B7",
    x"BF6A7E31",
    x"BF6A7BAC",
    x"BF6A7926",
    x"BF6A76A1",
    x"BF6A741B",
    x"BF6A7195",
    x"BF6A6F0F",
    x"BF6A6C89",
    x"BF6A6A02",
    x"BF6A677C",
    x"BF6A64F5",
    x"BF6A626E",
    x"BF6A5FE7",
    x"BF6A5D60",
    x"BF6A5AD9",
    x"BF6A5851",
    x"BF6A55CA",
    x"BF6A5342",
    x"BF6A50BA",
    x"BF6A4E33",
    x"BF6A4BAA",
    x"BF6A4922",
    x"BF6A469A",
    x"BF6A4411",
    x"BF6A4189",
    x"BF6A3F00",
    x"BF6A3C77",
    x"BF6A39EE",
    x"BF6A3765",
    x"BF6A34DB",
    x"BF6A3252",
    x"BF6A2FC8",
    x"BF6A2D3E",
    x"BF6A2AB4",
    x"BF6A282A",
    x"BF6A25A0",
    x"BF6A2316",
    x"BF6A208B",
    x"BF6A1E01",
    x"BF6A1B76",
    x"BF6A18EB",
    x"BF6A1660",
    x"BF6A13D5",
    x"BF6A1149",
    x"BF6A0EBE",
    x"BF6A0C32",
    x"BF6A09A7",
    x"BF6A071B",
    x"BF6A048F",
    x"BF6A0202",
    x"BF69FF76",
    x"BF69FCEA",
    x"BF69FA5D",
    x"BF69F7D0",
    x"BF69F543",
    x"BF69F2B6",
    x"BF69F029",
    x"BF69ED9C",
    x"BF69EB0E",
    x"BF69E881",
    x"BF69E5F3",
    x"BF69E365",
    x"BF69E0D7",
    x"BF69DE49",
    x"BF69DBBB",
    x"BF69D92C",
    x"BF69D69E",
    x"BF69D40F",
    x"BF69D180",
    x"BF69CEF1",
    x"BF69CC62",
    x"BF69C9D3",
    x"BF69C743",
    x"BF69C4B4",
    x"BF69C224",
    x"BF69BF94",
    x"BF69BD04",
    x"BF69BA74",
    x"BF69B7E4",
    x"BF69B553",
    x"BF69B2C3",
    x"BF69B032",
    x"BF69ADA1",
    x"BF69AB10",
    x"BF69A87F",
    x"BF69A5EE",
    x"BF69A35D",
    x"BF69A0CB",
    x"BF699E39",
    x"BF699BA8",
    x"BF699916",
    x"BF699684",
    x"BF6993F1",
    x"BF69915F",
    x"BF698ECC",
    x"BF698C3A",
    x"BF6989A7",
    x"BF698714",
    x"BF698481",
    x"BF6981EE",
    x"BF697F5A",
    x"BF697CC7",
    x"BF697A33",
    x"BF69779F",
    x"BF69750C",
    x"BF697277",
    x"BF696FE3",
    x"BF696D4F",
    x"BF696ABA",
    x"BF696826",
    x"BF696591",
    x"BF6962FC",
    x"BF696067",
    x"BF695DD2",
    x"BF695B3D",
    x"BF6958A7",
    x"BF695611",
    x"BF69537C",
    x"BF6950E6",
    x"BF694E50",
    x"BF694BBA",
    x"BF694923",
    x"BF69468D",
    x"BF6943F6",
    x"BF694160",
    x"BF693EC9",
    x"BF693C32",
    x"BF69399A",
    x"BF693703",
    x"BF69346C",
    x"BF6931D4",
    x"BF692F3C",
    x"BF692CA5",
    x"BF692A0D",
    x"BF692774",
    x"BF6924DC",
    x"BF692244",
    x"BF691FAB",
    x"BF691D12",
    x"BF691A7A",
    x"BF6917E1",
    x"BF691547",
    x"BF6912AE",
    x"BF691015",
    x"BF690D7B",
    x"BF690AE2",
    x"BF690848",
    x"BF6905AE",
    x"BF690314",
    x"BF690079",
    x"BF68FDDF",
    x"BF68FB45",
    x"BF68F8AA",
    x"BF68F60F",
    x"BF68F374",
    x"BF68F0D9",
    x"BF68EE3E",
    x"BF68EBA2",
    x"BF68E907",
    x"BF68E66B",
    x"BF68E3CF",
    x"BF68E134",
    x"BF68DE97",
    x"BF68DBFB",
    x"BF68D95F",
    x"BF68D6C2",
    x"BF68D426",
    x"BF68D189",
    x"BF68CEEC",
    x"BF68CC4F",
    x"BF68C9B2",
    x"BF68C714",
    x"BF68C477",
    x"BF68C1D9",
    x"BF68BF3C",
    x"BF68BC9E",
    x"BF68BA00",
    x"BF68B762",
    x"BF68B4C3",
    x"BF68B225",
    x"BF68AF86",
    x"BF68ACE7",
    x"BF68AA49",
    x"BF68A7AA",
    x"BF68A50A",
    x"BF68A26B",
    x"BF689FCC",
    x"BF689D2C",
    x"BF689A8C",
    x"BF6897EC",
    x"BF68954C",
    x"BF6892AC",
    x"BF68900C",
    x"BF688D6C",
    x"BF688ACB",
    x"BF68882A",
    x"BF68858A",
    x"BF6882E9",
    x"BF688047",
    x"BF687DA6",
    x"BF687B05",
    x"BF687863",
    x"BF6875C2",
    x"BF687320",
    x"BF68707E",
    x"BF686DDC",
    x"BF686B39",
    x"BF686897",
    x"BF6865F5",
    x"BF686352",
    x"BF6860AF",
    x"BF685E0C",
    x"BF685B69",
    x"BF6858C6",
    x"BF685623",
    x"BF68537F",
    x"BF6850DB",
    x"BF684E38",
    x"BF684B94",
    x"BF6848F0",
    x"BF68464B",
    x"BF6843A7",
    x"BF684103",
    x"BF683E5E",
    x"BF683BB9",
    x"BF683914",
    x"BF68366F",
    x"BF6833CA",
    x"BF683125",
    x"BF682E7F",
    x"BF682BDA",
    x"BF682934",
    x"BF68268E",
    x"BF6823E8",
    x"BF682142",
    x"BF681E9C",
    x"BF681BF5",
    x"BF68194F",
    x"BF6816A8",
    x"BF681401",
    x"BF68115A",
    x"BF680EB3",
    x"BF680C0C",
    x"BF680964",
    x"BF6806BD",
    x"BF680415",
    x"BF68016D",
    x"BF67FEC5",
    x"BF67FC1D",
    x"BF67F975",
    x"BF67F6CC",
    x"BF67F424",
    x"BF67F17B",
    x"BF67EED2",
    x"BF67EC29",
    x"BF67E980",
    x"BF67E6D7",
    x"BF67E42E",
    x"BF67E184",
    x"BF67DEDB",
    x"BF67DC31",
    x"BF67D987",
    x"BF67D6DD",
    x"BF67D433",
    x"BF67D188",
    x"BF67CEDE",
    x"BF67CC33",
    x"BF67C988",
    x"BF67C6DE",
    x"BF67C432",
    x"BF67C187",
    x"BF67BEDC",
    x"BF67BC30",
    x"BF67B985",
    x"BF67B6D9",
    x"BF67B42D",
    x"BF67B181",
    x"BF67AED5",
    x"BF67AC29",
    x"BF67A97C",
    x"BF67A6D0",
    x"BF67A423",
    x"BF67A176",
    x"BF679EC9",
    x"BF679C1C",
    x"BF67996F",
    x"BF6796C1",
    x"BF679414",
    x"BF679166",
    x"BF678EB8",
    x"BF678C0A",
    x"BF67895C",
    x"BF6786AE",
    x"BF6783FF",
    x"BF678151",
    x"BF677EA2",
    x"BF677BF3",
    x"BF677944",
    x"BF677695",
    x"BF6773E6",
    x"BF677137",
    x"BF676E87",
    x"BF676BD8",
    x"BF676928",
    x"BF676678",
    x"BF6763C8",
    x"BF676118",
    x"BF675E67",
    x"BF675BB7",
    x"BF675906",
    x"BF675655",
    x"BF6753A5",
    x"BF6750F3",
    x"BF674E42",
    x"BF674B91",
    x"BF6748DF",
    x"BF67462E",
    x"BF67437C",
    x"BF6740CA",
    x"BF673E18",
    x"BF673B66",
    x"BF6738B4",
    x"BF673601",
    x"BF67334F",
    x"BF67309C",
    x"BF672DE9",
    x"BF672B36",
    x"BF672883",
    x"BF6725D0",
    x"BF67231C",
    x"BF672069",
    x"BF671DB5",
    x"BF671B01",
    x"BF67184D",
    x"BF671599",
    x"BF6712E5",
    x"BF671031",
    x"BF670D7C",
    x"BF670AC7",
    x"BF670813",
    x"BF67055E",
    x"BF6702A9",
    x"BF66FFF3",
    x"BF66FD3E",
    x"BF66FA88",
    x"BF66F7D3",
    x"BF66F51D",
    x"BF66F267",
    x"BF66EFB1",
    x"BF66ECFB",
    x"BF66EA45",
    x"BF66E78E",
    x"BF66E4D7",
    x"BF66E221",
    x"BF66DF6A",
    x"BF66DCB3",
    x"BF66D9FC",
    x"BF66D744",
    x"BF66D48D",
    x"BF66D1D5",
    x"BF66CF1E",
    x"BF66CC66",
    x"BF66C9AE",
    x"BF66C6F6",
    x"BF66C43D",
    x"BF66C185",
    x"BF66BECC",
    x"BF66BC14",
    x"BF66B95B",
    x"BF66B6A2",
    x"BF66B3E9",
    x"BF66B12F",
    x"BF66AE76",
    x"BF66ABBC",
    x"BF66A903",
    x"BF66A649",
    x"BF66A38F",
    x"BF66A0D5",
    x"BF669E1B",
    x"BF669B60",
    x"BF6698A6",
    x"BF6695EB",
    x"BF669330",
    x"BF669076",
    x"BF668DBA",
    x"BF668AFF",
    x"BF668844",
    x"BF668588",
    x"BF6682CD",
    x"BF668011",
    x"BF667D55",
    x"BF667A99",
    x"BF6677DD",
    x"BF667521",
    x"BF667264",
    x"BF666FA8",
    x"BF666CEB",
    x"BF666A2E",
    x"BF666771",
    x"BF6664B4",
    x"BF6661F7",
    x"BF665F39",
    x"BF665C7C",
    x"BF6659BE",
    x"BF665700",
    x"BF665442",
    x"BF665184",
    x"BF664EC6",
    x"BF664C07",
    x"BF664949",
    x"BF66468A",
    x"BF6643CB",
    x"BF66410C",
    x"BF663E4D",
    x"BF663B8E",
    x"BF6638CF",
    x"BF66360F",
    x"BF663350",
    x"BF663090",
    x"BF662DD0",
    x"BF662B10",
    x"BF662850",
    x"BF66258F",
    x"BF6622CF",
    x"BF66200E",
    x"BF661D4D",
    x"BF661A8D",
    x"BF6617CC",
    x"BF66150A",
    x"BF661249",
    x"BF660F88",
    x"BF660CC6",
    x"BF660A04",
    x"BF660742",
    x"BF660480",
    x"BF6601BE",
    x"BF65FEFC",
    x"BF65FC3A",
    x"BF65F977",
    x"BF65F6B4",
    x"BF65F3F2",
    x"BF65F12F",
    x"BF65EE6C",
    x"BF65EBA8",
    x"BF65E8E5",
    x"BF65E621",
    x"BF65E35E",
    x"BF65E09A",
    x"BF65DDD6",
    x"BF65DB12",
    x"BF65D84E",
    x"BF65D589",
    x"BF65D2C5",
    x"BF65D000",
    x"BF65CD3B",
    x"BF65CA77",
    x"BF65C7B1",
    x"BF65C4EC",
    x"BF65C227",
    x"BF65BF62",
    x"BF65BC9C",
    x"BF65B9D6",
    x"BF65B710",
    x"BF65B44A",
    x"BF65B184",
    x"BF65AEBE",
    x"BF65ABF7",
    x"BF65A931",
    x"BF65A66A",
    x"BF65A3A3",
    x"BF65A0DC",
    x"BF659E15",
    x"BF659B4E",
    x"BF659887",
    x"BF6595BF",
    x"BF6592F7",
    x"BF659030",
    x"BF658D68",
    x"BF658AA0",
    x"BF6587D7",
    x"BF65850F",
    x"BF658246",
    x"BF657F7E",
    x"BF657CB5",
    x"BF6579EC",
    x"BF657723",
    x"BF65745A",
    x"BF657190",
    x"BF656EC7",
    x"BF656BFD",
    x"BF656934",
    x"BF65666A",
    x"BF6563A0",
    x"BF6560D6",
    x"BF655E0B",
    x"BF655B41",
    x"BF655876",
    x"BF6555AC",
    x"BF6552E1",
    x"BF655016",
    x"BF654D4B",
    x"BF654A7F",
    x"BF6547B4",
    x"BF6544E8",
    x"BF65421D",
    x"BF653F51",
    x"BF653C85",
    x"BF6539B9",
    x"BF6536ED",
    x"BF653420",
    x"BF653154",
    x"BF652E87",
    x"BF652BBA",
    x"BF6528ED",
    x"BF652620",
    x"BF652353",
    x"BF652086",
    x"BF651DB8",
    x"BF651AEB",
    x"BF65181D",
    x"BF65154F",
    x"BF651281",
    x"BF650FB3",
    x"BF650CE5",
    x"BF650A16",
    x"BF650748",
    x"BF650479",
    x"BF6501AA",
    x"BF64FEDB",
    x"BF64FC0C",
    x"BF64F93D",
    x"BF64F66D",
    x"BF64F39E",
    x"BF64F0CE",
    x"BF64EDFE",
    x"BF64EB2E",
    x"BF64E85E",
    x"BF64E58E",
    x"BF64E2BD",
    x"BF64DFED",
    x"BF64DD1C",
    x"BF64DA4B",
    x"BF64D77B",
    x"BF64D4AA",
    x"BF64D1D8",
    x"BF64CF07",
    x"BF64CC35",
    x"BF64C964",
    x"BF64C692",
    x"BF64C3C0",
    x"BF64C0EE",
    x"BF64BE1C",
    x"BF64BB4A",
    x"BF64B877",
    x"BF64B5A5",
    x"BF64B2D2",
    x"BF64AFFF",
    x"BF64AD2C",
    x"BF64AA59",
    x"BF64A786",
    x"BF64A4B2",
    x"BF64A1DF",
    x"BF649F0B",
    x"BF649C37",
    x"BF649963",
    x"BF64968F",
    x"BF6493BB",
    x"BF6490E7",
    x"BF648E12",
    x"BF648B3E",
    x"BF648869",
    x"BF648594",
    x"BF6482BF",
    x"BF647FEA",
    x"BF647D14",
    x"BF647A3F",
    x"BF647769",
    x"BF647493",
    x"BF6471BE",
    x"BF646EE8",
    x"BF646C11",
    x"BF64693B",
    x"BF646665",
    x"BF64638E",
    x"BF6460B7",
    x"BF645DE1",
    x"BF645B0A",
    x"BF645832",
    x"BF64555B",
    x"BF645284",
    x"BF644FAC",
    x"BF644CD5",
    x"BF6449FD",
    x"BF644725",
    x"BF64444D",
    x"BF644174",
    x"BF643E9C",
    x"BF643BC4",
    x"BF6438EB",
    x"BF643612",
    x"BF643339",
    x"BF643060",
    x"BF642D87",
    x"BF642AAE",
    x"BF6427D4",
    x"BF6424FB",
    x"BF642221",
    x"BF641F47",
    x"BF641C6D",
    x"BF641993",
    x"BF6416B9",
    x"BF6413DE",
    x"BF641104",
    x"BF640E29",
    x"BF640B4E",
    x"BF640873",
    x"BF640598",
    x"BF6402BD",
    x"BF63FFE1",
    x"BF63FD06",
    x"BF63FA2A",
    x"BF63F74E",
    x"BF63F473",
    x"BF63F196",
    x"BF63EEBA",
    x"BF63EBDE",
    x"BF63E901",
    x"BF63E625",
    x"BF63E348",
    x"BF63E06B",
    x"BF63DD8E",
    x"BF63DAB1",
    x"BF63D7D4",
    x"BF63D4F6",
    x"BF63D219",
    x"BF63CF3B",
    x"BF63CC5D",
    x"BF63C97F",
    x"BF63C6A1",
    x"BF63C3C3",
    x"BF63C0E4",
    x"BF63BE06",
    x"BF63BB27",
    x"BF63B848",
    x"BF63B569",
    x"BF63B28A",
    x"BF63AFAB",
    x"BF63ACCC",
    x"BF63A9EC",
    x"BF63A70D",
    x"BF63A42D",
    x"BF63A14D",
    x"BF639E6D",
    x"BF639B8D",
    x"BF6398AC",
    x"BF6395CC",
    x"BF6392EB",
    x"BF63900B",
    x"BF638D2A",
    x"BF638A49",
    x"BF638767",
    x"BF638486",
    x"BF6381A5",
    x"BF637EC3",
    x"BF637BE2",
    x"BF637900",
    x"BF63761E",
    x"BF63733C",
    x"BF637059",
    x"BF636D77",
    x"BF636A95",
    x"BF6367B2",
    x"BF6364CF",
    x"BF6361EC",
    x"BF635F09",
    x"BF635C26",
    x"BF635943",
    x"BF63565F",
    x"BF63537B",
    x"BF635098",
    x"BF634DB4",
    x"BF634AD0",
    x"BF6347EC",
    x"BF634507",
    x"BF634223",
    x"BF633F3E",
    x"BF633C5A",
    x"BF633975",
    x"BF633690",
    x"BF6333AB",
    x"BF6330C5",
    x"BF632DE0",
    x"BF632AFB",
    x"BF632815",
    x"BF63252F",
    x"BF632249",
    x"BF631F63",
    x"BF631C7D",
    x"BF631996",
    x"BF6316B0",
    x"BF6313C9",
    x"BF6310E3",
    x"BF630DFC",
    x"BF630B15",
    x"BF63082E",
    x"BF630546",
    x"BF63025F",
    x"BF62FF77",
    x"BF62FC8F",
    x"BF62F9A8",
    x"BF62F6C0",
    x"BF62F3D8",
    x"BF62F0EF",
    x"BF62EE07",
    x"BF62EB1E",
    x"BF62E836",
    x"BF62E54D",
    x"BF62E264",
    x"BF62DF7B",
    x"BF62DC92",
    x"BF62D9A8",
    x"BF62D6BF",
    x"BF62D3D5",
    x"BF62D0EB",
    x"BF62CE01",
    x"BF62CB17",
    x"BF62C82D",
    x"BF62C543",
    x"BF62C258",
    x"BF62BF6E",
    x"BF62BC83",
    x"BF62B998",
    x"BF62B6AD",
    x"BF62B3C2",
    x"BF62B0D7",
    x"BF62ADEB",
    x"BF62AB00",
    x"BF62A814",
    x"BF62A528",
    x"BF62A23D",
    x"BF629F50",
    x"BF629C64",
    x"BF629978",
    x"BF62968B",
    x"BF62939F",
    x"BF6290B2",
    x"BF628DC5",
    x"BF628AD8",
    x"BF6287EB",
    x"BF6284FD",
    x"BF628210",
    x"BF627F22",
    x"BF627C35",
    x"BF627947",
    x"BF627659",
    x"BF62736B",
    x"BF62707C",
    x"BF626D8E",
    x"BF626AA0",
    x"BF6267B1",
    x"BF6264C2",
    x"BF6261D3",
    x"BF625EE4",
    x"BF625BF5",
    x"BF625905",
    x"BF625616",
    x"BF625326",
    x"BF625036",
    x"BF624D47",
    x"BF624A57",
    x"BF624766",
    x"BF624476",
    x"BF624186",
    x"BF623E95",
    x"BF623BA4",
    x"BF6238B3",
    x"BF6235C2",
    x"BF6232D1",
    x"BF622FE0",
    x"BF622CEF",
    x"BF6229FD",
    x"BF62270B",
    x"BF62241A",
    x"BF622128",
    x"BF621E35",
    x"BF621B43",
    x"BF621851",
    x"BF62155E",
    x"BF62126C",
    x"BF620F79",
    x"BF620C86",
    x"BF620993",
    x"BF6206A0",
    x"BF6203AD",
    x"BF6200B9",
    x"BF61FDC6",
    x"BF61FAD2",
    x"BF61F7DE",
    x"BF61F4EA",
    x"BF61F1F6",
    x"BF61EF02",
    x"BF61EC0D",
    x"BF61E919",
    x"BF61E624",
    x"BF61E32F",
    x"BF61E03A",
    x"BF61DD45",
    x"BF61DA50",
    x"BF61D75B",
    x"BF61D465",
    x"BF61D16F",
    x"BF61CE7A",
    x"BF61CB84",
    x"BF61C88E",
    x"BF61C598",
    x"BF61C2A1",
    x"BF61BFAB",
    x"BF61BCB4",
    x"BF61B9BE",
    x"BF61B6C7",
    x"BF61B3D0",
    x"BF61B0D9",
    x"BF61ADE1",
    x"BF61AAEA",
    x"BF61A7F2",
    x"BF61A4FB",
    x"BF61A203",
    x"BF619F0B",
    x"BF619C13",
    x"BF61991B",
    x"BF619622",
    x"BF61932A",
    x"BF619031",
    x"BF618D38",
    x"BF618A40",
    x"BF618747",
    x"BF61844D",
    x"BF618154",
    x"BF617E5B",
    x"BF617B61",
    x"BF617867",
    x"BF61756E",
    x"BF617274",
    x"BF616F79",
    x"BF616C7F",
    x"BF616985",
    x"BF61668A",
    x"BF616390",
    x"BF616095",
    x"BF615D9A",
    x"BF615A9F",
    x"BF6157A4",
    x"BF6154A8",
    x"BF6151AD",
    x"BF614EB1",
    x"BF614BB5",
    x"BF6148BA",
    x"BF6145BE",
    x"BF6142C1",
    x"BF613FC5",
    x"BF613CC9",
    x"BF6139CC",
    x"BF6136D0",
    x"BF6133D3",
    x"BF6130D6",
    x"BF612DD9",
    x"BF612ADB",
    x"BF6127DE",
    x"BF6124E1",
    x"BF6121E3",
    x"BF611EE5",
    x"BF611BE7",
    x"BF6118E9",
    x"BF6115EB",
    x"BF6112ED",
    x"BF610FEE",
    x"BF610CF0",
    x"BF6109F1",
    x"BF6106F2",
    x"BF6103F3",
    x"BF6100F4",
    x"BF60FDF5",
    x"BF60FAF5",
    x"BF60F7F6",
    x"BF60F4F6",
    x"BF60F1F6",
    x"BF60EEF6",
    x"BF60EBF6",
    x"BF60E8F6",
    x"BF60E5F6",
    x"BF60E2F5",
    x"BF60DFF4",
    x"BF60DCF4",
    x"BF60D9F3",
    x"BF60D6F2",
    x"BF60D3F1",
    x"BF60D0EF",
    x"BF60CDEE",
    x"BF60CAEC",
    x"BF60C7EB",
    x"BF60C4E9",
    x"BF60C1E7",
    x"BF60BEE5",
    x"BF60BBE2",
    x"BF60B8E0",
    x"BF60B5DE",
    x"BF60B2DB",
    x"BF60AFD8",
    x"BF60ACD5",
    x"BF60A9D2",
    x"BF60A6CF",
    x"BF60A3CC",
    x"BF60A0C8",
    x"BF609DC4",
    x"BF609AC1",
    x"BF6097BD",
    x"BF6094B9",
    x"BF6091B5",
    x"BF608EB0",
    x"BF608BAC",
    x"BF6088A7",
    x"BF6085A3",
    x"BF60829E",
    x"BF607F99",
    x"BF607C94",
    x"BF60798F",
    x"BF607689",
    x"BF607384",
    x"BF60707E",
    x"BF606D78",
    x"BF606A73",
    x"BF60676D",
    x"BF606466",
    x"BF606160",
    x"BF605E5A",
    x"BF605B53",
    x"BF60584C",
    x"BF605545",
    x"BF60523E",
    x"BF604F37",
    x"BF604C30",
    x"BF604929",
    x"BF604621",
    x"BF60431A",
    x"BF604012",
    x"BF603D0A",
    x"BF603A02",
    x"BF6036FA",
    x"BF6033F1",
    x"BF6030E9",
    x"BF602DE0",
    x"BF602AD7",
    x"BF6027CF",
    x"BF6024C6",
    x"BF6021BC",
    x"BF601EB3",
    x"BF601BAA",
    x"BF6018A0",
    x"BF601596",
    x"BF60128D",
    x"BF600F83",
    x"BF600C79",
    x"BF60096E",
    x"BF600664",
    x"BF60035A",
    x"BF60004F",
    x"BF5FFD44",
    x"BF5FFA39",
    x"BF5FF72E",
    x"BF5FF423",
    x"BF5FF118",
    x"BF5FEE0C",
    x"BF5FEB01",
    x"BF5FE7F5",
    x"BF5FE4E9",
    x"BF5FE1DD",
    x"BF5FDED1",
    x"BF5FDBC5",
    x"BF5FD8B8",
    x"BF5FD5AC",
    x"BF5FD29F",
    x"BF5FCF93",
    x"BF5FCC86",
    x"BF5FC979",
    x"BF5FC66B",
    x"BF5FC35E",
    x"BF5FC051",
    x"BF5FBD43",
    x"BF5FBA35",
    x"BF5FB727",
    x"BF5FB419",
    x"BF5FB10B",
    x"BF5FADFD",
    x"BF5FAAEF",
    x"BF5FA7E0",
    x"BF5FA4D1",
    x"BF5FA1C3",
    x"BF5F9EB4",
    x"BF5F9BA5",
    x"BF5F9895",
    x"BF5F9586",
    x"BF5F9276",
    x"BF5F8F67",
    x"BF5F8C57",
    x"BF5F8947",
    x"BF5F8637",
    x"BF5F8327",
    x"BF5F8017",
    x"BF5F7D06",
    x"BF5F79F6",
    x"BF5F76E5",
    x"BF5F73D4",
    x"BF5F70C3",
    x"BF5F6DB2",
    x"BF5F6AA1",
    x"BF5F6790",
    x"BF5F647E",
    x"BF5F616C",
    x"BF5F5E5B",
    x"BF5F5B49",
    x"BF5F5837",
    x"BF5F5525",
    x"BF5F5212",
    x"BF5F4F00",
    x"BF5F4BED",
    x"BF5F48DB",
    x"BF5F45C8",
    x"BF5F42B5",
    x"BF5F3FA2",
    x"BF5F3C8E",
    x"BF5F397B",
    x"BF5F3667",
    x"BF5F3354",
    x"BF5F3040",
    x"BF5F2D2C",
    x"BF5F2A18",
    x"BF5F2704",
    x"BF5F23EF",
    x"BF5F20DB",
    x"BF5F1DC6",
    x"BF5F1AB2",
    x"BF5F179D",
    x"BF5F1488",
    x"BF5F1173",
    x"BF5F0E5D",
    x"BF5F0B48",
    x"BF5F0833",
    x"BF5F051D",
    x"BF5F0207",
    x"BF5EFEF1",
    x"BF5EFBDB",
    x"BF5EF8C5",
    x"BF5EF5AE",
    x"BF5EF298",
    x"BF5EEF81",
    x"BF5EEC6B",
    x"BF5EE954",
    x"BF5EE63D",
    x"BF5EE326",
    x"BF5EE00E",
    x"BF5EDCF7",
    x"BF5ED9DF",
    x"BF5ED6C8",
    x"BF5ED3B0",
    x"BF5ED098",
    x"BF5ECD80",
    x"BF5ECA68",
    x"BF5EC74F",
    x"BF5EC437",
    x"BF5EC11E",
    x"BF5EBE05",
    x"BF5EBAEC",
    x"BF5EB7D3",
    x"BF5EB4BA",
    x"BF5EB1A1",
    x"BF5EAE88",
    x"BF5EAB6E",
    x"BF5EA854",
    x"BF5EA53A",
    x"BF5EA221",
    x"BF5E9F06",
    x"BF5E9BEC",
    x"BF5E98D2",
    x"BF5E95B7",
    x"BF5E929D",
    x"BF5E8F82",
    x"BF5E8C67",
    x"BF5E894C",
    x"BF5E8631",
    x"BF5E8316",
    x"BF5E7FFA",
    x"BF5E7CDE",
    x"BF5E79C3",
    x"BF5E76A7",
    x"BF5E738B",
    x"BF5E706F",
    x"BF5E6D53",
    x"BF5E6A36",
    x"BF5E671A",
    x"BF5E63FD",
    x"BF5E60E0",
    x"BF5E5DC3",
    x"BF5E5AA6",
    x"BF5E5789",
    x"BF5E546C",
    x"BF5E514E",
    x"BF5E4E31",
    x"BF5E4B13",
    x"BF5E47F5",
    x"BF5E44D7",
    x"BF5E41B9",
    x"BF5E3E9B",
    x"BF5E3B7D",
    x"BF5E385E",
    x"BF5E353F",
    x"BF5E3221",
    x"BF5E2F02",
    x"BF5E2BE3",
    x"BF5E28C3",
    x"BF5E25A4",
    x"BF5E2285",
    x"BF5E1F65",
    x"BF5E1C45",
    x"BF5E1925",
    x"BF5E1605",
    x"BF5E12E5",
    x"BF5E0FC5",
    x"BF5E0CA5",
    x"BF5E0984",
    x"BF5E0663",
    x"BF5E0343",
    x"BF5E0022",
    x"BF5DFD01",
    x"BF5DF9DF",
    x"BF5DF6BE",
    x"BF5DF39D",
    x"BF5DF07B",
    x"BF5DED59",
    x"BF5DEA37",
    x"BF5DE715",
    x"BF5DE3F3",
    x"BF5DE0D1",
    x"BF5DDDAF",
    x"BF5DDA8C",
    x"BF5DD769",
    x"BF5DD447",
    x"BF5DD124",
    x"BF5DCE01",
    x"BF5DCADD",
    x"BF5DC7BA",
    x"BF5DC497",
    x"BF5DC173",
    x"BF5DBE4F",
    x"BF5DBB2B",
    x"BF5DB807",
    x"BF5DB4E3",
    x"BF5DB1BF",
    x"BF5DAE9B",
    x"BF5DAB76",
    x"BF5DA851",
    x"BF5DA52D",
    x"BF5DA208",
    x"BF5D9EE3",
    x"BF5D9BBD",
    x"BF5D9898",
    x"BF5D9573",
    x"BF5D924D",
    x"BF5D8F27",
    x"BF5D8C01",
    x"BF5D88DB",
    x"BF5D85B5",
    x"BF5D828F",
    x"BF5D7F69",
    x"BF5D7C42",
    x"BF5D791B",
    x"BF5D75F5",
    x"BF5D72CE",
    x"BF5D6FA7",
    x"BF5D6C7F",
    x"BF5D6958",
    x"BF5D6631",
    x"BF5D6309",
    x"BF5D5FE1",
    x"BF5D5CB9",
    x"BF5D5991",
    x"BF5D5669",
    x"BF5D5341",
    x"BF5D5018",
    x"BF5D4CF0",
    x"BF5D49C7",
    x"BF5D469E",
    x"BF5D4376",
    x"BF5D404C",
    x"BF5D3D23",
    x"BF5D39FA",
    x"BF5D36D0",
    x"BF5D33A7",
    x"BF5D307D",
    x"BF5D2D53",
    x"BF5D2A29",
    x"BF5D26FF",
    x"BF5D23D5",
    x"BF5D20AA",
    x"BF5D1D80",
    x"BF5D1A55",
    x"BF5D172A",
    x"BF5D13FF",
    x"BF5D10D4",
    x"BF5D0DA9",
    x"BF5D0A7E",
    x"BF5D0752",
    x"BF5D0427",
    x"BF5D00FB",
    x"BF5CFDCF",
    x"BF5CFAA3",
    x"BF5CF777",
    x"BF5CF44B",
    x"BF5CF11E",
    x"BF5CEDF2",
    x"BF5CEAC5",
    x"BF5CE798",
    x"BF5CE46B",
    x"BF5CE13E",
    x"BF5CDE11",
    x"BF5CDAE4",
    x"BF5CD7B6",
    x"BF5CD489",
    x"BF5CD15B",
    x"BF5CCE2D",
    x"BF5CCAFF",
    x"BF5CC7D1",
    x"BF5CC4A3",
    x"BF5CC174",
    x"BF5CBE46",
    x"BF5CBB17",
    x"BF5CB7E8",
    x"BF5CB4B9",
    x"BF5CB18A",
    x"BF5CAE5B",
    x"BF5CAB2C",
    x"BF5CA7FC",
    x"BF5CA4CD",
    x"BF5CA19D",
    x"BF5C9E6D",
    x"BF5C9B3D",
    x"BF5C980D",
    x"BF5C94DD",
    x"BF5C91AC",
    x"BF5C8E7C",
    x"BF5C8B4B",
    x"BF5C881A",
    x"BF5C84EA",
    x"BF5C81B8",
    x"BF5C7E87",
    x"BF5C7B56",
    x"BF5C7824",
    x"BF5C74F3",
    x"BF5C71C1",
    x"BF5C6E8F",
    x"BF5C6B5D",
    x"BF5C682B",
    x"BF5C64F9",
    x"BF5C61C7",
    x"BF5C5E94",
    x"BF5C5B61",
    x"BF5C582F",
    x"BF5C54FC",
    x"BF5C51C9",
    x"BF5C4E95",
    x"BF5C4B62",
    x"BF5C482F",
    x"BF5C44FB",
    x"BF5C41C7",
    x"BF5C3E94",
    x"BF5C3B60",
    x"BF5C382B",
    x"BF5C34F7",
    x"BF5C31C3",
    x"BF5C2E8E",
    x"BF5C2B5A",
    x"BF5C2825",
    x"BF5C24F0",
    x"BF5C21BB",
    x"BF5C1E86",
    x"BF5C1B51",
    x"BF5C181B",
    x"BF5C14E6",
    x"BF5C11B0",
    x"BF5C0E7A",
    x"BF5C0B44",
    x"BF5C080E",
    x"BF5C04D8",
    x"BF5C01A1",
    x"BF5BFE6B",
    x"BF5BFB34",
    x"BF5BF7FD",
    x"BF5BF4C7",
    x"BF5BF190",
    x"BF5BEE58",
    x"BF5BEB21",
    x"BF5BE7EA",
    x"BF5BE4B2",
    x"BF5BE17A",
    x"BF5BDE43",
    x"BF5BDB0B",
    x"BF5BD7D3",
    x"BF5BD49A",
    x"BF5BD162",
    x"BF5BCE29",
    x"BF5BCAF1",
    x"BF5BC7B8",
    x"BF5BC47F",
    x"BF5BC146",
    x"BF5BBE0D",
    x"BF5BBAD4",
    x"BF5BB79A",
    x"BF5BB461",
    x"BF5BB127",
    x"BF5BADED",
    x"BF5BAAB3",
    x"BF5BA779",
    x"BF5BA43F",
    x"BF5BA105",
    x"BF5B9DCA",
    x"BF5B9A90",
    x"BF5B9755",
    x"BF5B941A",
    x"BF5B90DF",
    x"BF5B8DA4",
    x"BF5B8A69",
    x"BF5B872D",
    x"BF5B83F2",
    x"BF5B80B6",
    x"BF5B7D7A",
    x"BF5B7A3E",
    x"BF5B7702",
    x"BF5B73C6",
    x"BF5B708A",
    x"BF5B6D4D",
    x"BF5B6A11",
    x"BF5B66D4",
    x"BF5B6397",
    x"BF5B605A",
    x"BF5B5D1D",
    x"BF5B59E0",
    x"BF5B56A3",
    x"BF5B5365",
    x"BF5B5027",
    x"BF5B4CEA",
    x"BF5B49AC",
    x"BF5B466E",
    x"BF5B4330",
    x"BF5B3FF1",
    x"BF5B3CB3",
    x"BF5B3974",
    x"BF5B3636",
    x"BF5B32F7",
    x"BF5B2FB8",
    x"BF5B2C79",
    x"BF5B2939",
    x"BF5B25FA",
    x"BF5B22BB",
    x"BF5B1F7B",
    x"BF5B1C3B",
    x"BF5B18FB",
    x"BF5B15BB",
    x"BF5B127B",
    x"BF5B0F3B",
    x"BF5B0BFA",
    x"BF5B08BA",
    x"BF5B0579",
    x"BF5B0238",
    x"BF5AFEF7",
    x"BF5AFBB6",
    x"BF5AF875",
    x"BF5AF534",
    x"BF5AF1F2",
    x"BF5AEEB1",
    x"BF5AEB6F",
    x"BF5AE82D",
    x"BF5AE4EB",
    x"BF5AE1A9",
    x"BF5ADE67",
    x"BF5ADB24",
    x"BF5AD7E2",
    x"BF5AD49F",
    x"BF5AD15C",
    x"BF5ACE1A",
    x"BF5ACAD6",
    x"BF5AC793",
    x"BF5AC450",
    x"BF5AC10D",
    x"BF5ABDC9",
    x"BF5ABA85",
    x"BF5AB741",
    x"BF5AB3FD",
    x"BF5AB0B9",
    x"BF5AAD75",
    x"BF5AAA31",
    x"BF5AA6EC",
    x"BF5AA3A8",
    x"BF5AA063",
    x"BF5A9D1E",
    x"BF5A99D9",
    x"BF5A9694",
    x"BF5A934E",
    x"BF5A9009",
    x"BF5A8CC3",
    x"BF5A897E",
    x"BF5A8638",
    x"BF5A82F2",
    x"BF5A7FAC",
    x"BF5A7C66",
    x"BF5A791F",
    x"BF5A75D9",
    x"BF5A7292",
    x"BF5A6F4C",
    x"BF5A6C05",
    x"BF5A68BE",
    x"BF5A6577",
    x"BF5A622F",
    x"BF5A5EE8",
    x"BF5A5BA0",
    x"BF5A5859",
    x"BF5A5511",
    x"BF5A51C9",
    x"BF5A4E81",
    x"BF5A4B39",
    x"BF5A47F0",
    x"BF5A44A8",
    x"BF5A415F",
    x"BF5A3E17",
    x"BF5A3ACE",
    x"BF5A3785",
    x"BF5A343C",
    x"BF5A30F2",
    x"BF5A2DA9",
    x"BF5A2A60",
    x"BF5A2716",
    x"BF5A23CC",
    x"BF5A2082",
    x"BF5A1D38",
    x"BF5A19EE",
    x"BF5A16A4",
    x"BF5A1359",
    x"BF5A100F",
    x"BF5A0CC4",
    x"BF5A0979",
    x"BF5A062E",
    x"BF5A02E3",
    x"BF59FF98",
    x"BF59FC4D",
    x"BF59F901",
    x"BF59F5B6",
    x"BF59F26A",
    x"BF59EF1E",
    x"BF59EBD2",
    x"BF59E886",
    x"BF59E53A",
    x"BF59E1ED",
    x"BF59DEA1",
    x"BF59DB54",
    x"BF59D807",
    x"BF59D4BA",
    x"BF59D16D",
    x"BF59CE20",
    x"BF59CAD3",
    x"BF59C785",
    x"BF59C438",
    x"BF59C0EA",
    x"BF59BD9C",
    x"BF59BA4E",
    x"BF59B700",
    x"BF59B3B2",
    x"BF59B064",
    x"BF59AD15",
    x"BF59A9C7",
    x"BF59A678",
    x"BF59A329",
    x"BF599FDA",
    x"BF599C8B",
    x"BF59993C",
    x"BF5995EC",
    x"BF59929D",
    x"BF598F4D",
    x"BF598BFD",
    x"BF5988AD",
    x"BF59855D",
    x"BF59820D",
    x"BF597EBD",
    x"BF597B6C",
    x"BF59781C",
    x"BF5974CB",
    x"BF59717A",
    x"BF596E29",
    x"BF596AD8",
    x"BF596787",
    x"BF596435",
    x"BF5960E4",
    x"BF595D92",
    x"BF595A40",
    x"BF5956EE",
    x"BF59539C",
    x"BF59504A",
    x"BF594CF8",
    x"BF5949A6",
    x"BF594653",
    x"BF594300",
    x"BF593FAE",
    x"BF593C5B",
    x"BF593908",
    x"BF5935B4",
    x"BF593261",
    x"BF592F0E",
    x"BF592BBA",
    x"BF592866",
    x"BF592512",
    x"BF5921BE",
    x"BF591E6A",
    x"BF591B16",
    x"BF5917C2",
    x"BF59146D",
    x"BF591118",
    x"BF590DC4",
    x"BF590A6F",
    x"BF59071A",
    x"BF5903C5",
    x"BF59006F",
    x"BF58FD1A",
    x"BF58F9C4",
    x"BF58F66F",
    x"BF58F319",
    x"BF58EFC3",
    x"BF58EC6D",
    x"BF58E916",
    x"BF58E5C0",
    x"BF58E26A",
    x"BF58DF13",
    x"BF58DBBC",
    x"BF58D865",
    x"BF58D50E",
    x"BF58D1B7",
    x"BF58CE60",
    x"BF58CB09",
    x"BF58C7B1",
    x"BF58C45A",
    x"BF58C102",
    x"BF58BDAA",
    x"BF58BA52",
    x"BF58B6FA",
    x"BF58B3A1",
    x"BF58B049",
    x"BF58ACF0",
    x"BF58A998",
    x"BF58A63F",
    x"BF58A2E6",
    x"BF589F8D",
    x"BF589C34",
    x"BF5898DA",
    x"BF589581",
    x"BF589227",
    x"BF588ECD",
    x"BF588B74",
    x"BF58881A",
    x"BF5884BF",
    x"BF588165",
    x"BF587E0B",
    x"BF587AB0",
    x"BF587756",
    x"BF5873FB",
    x"BF5870A0",
    x"BF586D45",
    x"BF5869EA",
    x"BF58668E",
    x"BF586333",
    x"BF585FD7",
    x"BF585C7C",
    x"BF585920",
    x"BF5855C4",
    x"BF585268",
    x"BF584F0C",
    x"BF584BAF",
    x"BF584853",
    x"BF5844F6",
    x"BF584199",
    x"BF583E3D",
    x"BF583AE0",
    x"BF583782",
    x"BF583425",
    x"BF5830C8",
    x"BF582D6A",
    x"BF582A0D",
    x"BF5826AF",
    x"BF582351",
    x"BF581FF3",
    x"BF581C95",
    x"BF581936",
    x"BF5815D8",
    x"BF581279",
    x"BF580F1B",
    x"BF580BBC",
    x"BF58085D",
    x"BF5804FE",
    x"BF58019F",
    x"BF57FE3F",
    x"BF57FAE0",
    x"BF57F780",
    x"BF57F421",
    x"BF57F0C1",
    x"BF57ED61",
    x"BF57EA01",
    x"BF57E6A0",
    x"BF57E340",
    x"BF57DFDF",
    x"BF57DC7F",
    x"BF57D91E",
    x"BF57D5BD",
    x"BF57D25C",
    x"BF57CEFB",
    x"BF57CB9A",
    x"BF57C838",
    x"BF57C4D7",
    x"BF57C175",
    x"BF57BE13",
    x"BF57BAB1",
    x"BF57B74F",
    x"BF57B3ED",
    x"BF57B08B",
    x"BF57AD28",
    x"BF57A9C6",
    x"BF57A663",
    x"BF57A300",
    x"BF579F9D",
    x"BF579C3A",
    x"BF5798D7",
    x"BF579573",
    x"BF579210",
    x"BF578EAC",
    x"BF578B48",
    x"BF5787E4",
    x"BF578480",
    x"BF57811C",
    x"BF577DB8",
    x"BF577A54",
    x"BF5776EF",
    x"BF57738A",
    x"BF577026",
    x"BF576CC1",
    x"BF57695C",
    x"BF5765F6",
    x"BF576291",
    x"BF575F2C",
    x"BF575BC6",
    x"BF575860",
    x"BF5754FB",
    x"BF575195",
    x"BF574E2F",
    x"BF574AC8",
    x"BF574762",
    x"BF5743FB",
    x"BF574095",
    x"BF573D2E",
    x"BF5739C7",
    x"BF573660",
    x"BF5732F9",
    x"BF572F92",
    x"BF572C2A",
    x"BF5728C3",
    x"BF57255B",
    x"BF5721F3",
    x"BF571E8C",
    x"BF571B24",
    x"BF5717BB",
    x"BF571453",
    x"BF5710EB",
    x"BF570D82",
    x"BF570A19",
    x"BF5706B1",
    x"BF570348",
    x"BF56FFDF",
    x"BF56FC75",
    x"BF56F90C",
    x"BF56F5A3",
    x"BF56F239",
    x"BF56EECF",
    x"BF56EB65",
    x"BF56E7FB",
    x"BF56E491",
    x"BF56E127",
    x"BF56DDBD",
    x"BF56DA52",
    x"BF56D6E8",
    x"BF56D37D",
    x"BF56D012",
    x"BF56CCA7",
    x"BF56C93C",
    x"BF56C5D0",
    x"BF56C265",
    x"BF56BEF9",
    x"BF56BB8E",
    x"BF56B822",
    x"BF56B4B6",
    x"BF56B14A",
    x"BF56ADDE",
    x"BF56AA72",
    x"BF56A705",
    x"BF56A399",
    x"BF56A02C",
    x"BF569CBF",
    x"BF569952",
    x"BF5695E5",
    x"BF569278",
    x"BF568F0A",
    x"BF568B9D",
    x"BF56882F",
    x"BF5684C2",
    x"BF568154",
    x"BF567DE6",
    x"BF567A78",
    x"BF567709",
    x"BF56739B",
    x"BF56702C",
    x"BF566CBE",
    x"BF56694F",
    x"BF5665E0",
    x"BF566271",
    x"BF565F02",
    x"BF565B93",
    x"BF565823",
    x"BF5654B4",
    x"BF565144",
    x"BF564DD4",
    x"BF564A64",
    x"BF5646F4",
    x"BF564384",
    x"BF564014",
    x"BF563CA3",
    x"BF563933",
    x"BF5635C2",
    x"BF563251",
    x"BF562EE0",
    x"BF562B6F",
    x"BF5627FE",
    x"BF56248D",
    x"BF56211B",
    x"BF561DA9",
    x"BF561A38",
    x"BF5616C6",
    x"BF561354",
    x"BF560FE2",
    x"BF560C70",
    x"BF5608FD",
    x"BF56058B",
    x"BF560218",
    x"BF55FEA5",
    x"BF55FB32",
    x"BF55F7BF",
    x"BF55F44C",
    x"BF55F0D9",
    x"BF55ED65",
    x"BF55E9F2",
    x"BF55E67E",
    x"BF55E30A",
    x"BF55DF96",
    x"BF55DC22",
    x"BF55D8AE",
    x"BF55D53A",
    x"BF55D1C5",
    x"BF55CE51",
    x"BF55CADC",
    x"BF55C767",
    x"BF55C3F2",
    x"BF55C07D",
    x"BF55BD08",
    x"BF55B993",
    x"BF55B61D",
    x"BF55B2A8",
    x"BF55AF32",
    x"BF55ABBC",
    x"BF55A846",
    x"BF55A4D0",
    x"BF55A15A",
    x"BF559DE3",
    x"BF559A6D",
    x"BF5596F6",
    x"BF55937F",
    x"BF559009",
    x"BF558C92",
    x"BF55891A",
    x"BF5585A3",
    x"BF55822C",
    x"BF557EB4",
    x"BF557B3D",
    x"BF5577C5",
    x"BF55744D",
    x"BF5570D5",
    x"BF556D5D",
    x"BF5569E4",
    x"BF55666C",
    x"BF5562F3",
    x"BF555F7B",
    x"BF555C02",
    x"BF555889",
    x"BF555510",
    x"BF555197",
    x"BF554E1D",
    x"BF554AA4",
    x"BF55472A",
    x"BF5543B1",
    x"BF554037",
    x"BF553CBD",
    x"BF553943",
    x"BF5535C8",
    x"BF55324E",
    x"BF552ED4",
    x"BF552B59",
    x"BF5527DE",
    x"BF552463",
    x"BF5520E8",
    x"BF551D6D",
    x"BF5519F2",
    x"BF551676",
    x"BF5512FB",
    x"BF550F7F",
    x"BF550C04",
    x"BF550888",
    x"BF55050C",
    x"BF55018F",
    x"BF54FE13",
    x"BF54FA97",
    x"BF54F71A",
    x"BF54F39E",
    x"BF54F021",
    x"BF54ECA4",
    x"BF54E927",
    x"BF54E5AA",
    x"BF54E22C",
    x"BF54DEAF",
    x"BF54DB31",
    x"BF54D7B4",
    x"BF54D436",
    x"BF54D0B8",
    x"BF54CD3A",
    x"BF54C9BC",
    x"BF54C63D",
    x"BF54C2BF",
    x"BF54BF40",
    x"BF54BBC1",
    x"BF54B843",
    x"BF54B4C4",
    x"BF54B144",
    x"BF54ADC5",
    x"BF54AA46",
    x"BF54A6C6",
    x"BF54A347",
    x"BF549FC7",
    x"BF549C47",
    x"BF5498C7",
    x"BF549547",
    x"BF5491C7",
    x"BF548E46",
    x"BF548AC6",
    x"BF548745",
    x"BF5483C4",
    x"BF548044",
    x"BF547CC3",
    x"BF547941",
    x"BF5475C0",
    x"BF54723F",
    x"BF546EBD",
    x"BF546B3B",
    x"BF5467BA",
    x"BF546438",
    x"BF5460B6",
    x"BF545D33",
    x"BF5459B1",
    x"BF54562F",
    x"BF5452AC",
    x"BF544F2A",
    x"BF544BA7",
    x"BF544824",
    x"BF5444A1",
    x"BF54411D",
    x"BF543D9A",
    x"BF543A17",
    x"BF543693",
    x"BF54330F",
    x"BF542F8C",
    x"BF542C08",
    x"BF542883",
    x"BF5424FF",
    x"BF54217B",
    x"BF541DF6",
    x"BF541A72",
    x"BF5416ED",
    x"BF541368",
    x"BF540FE3",
    x"BF540C5E",
    x"BF5408D9",
    x"BF540553",
    x"BF5401CE",
    x"BF53FE48",
    x"BF53FAC3",
    x"BF53F73D",
    x"BF53F3B7",
    x"BF53F031",
    x"BF53ECAA",
    x"BF53E924",
    x"BF53E59D",
    x"BF53E217",
    x"BF53DE90",
    x"BF53DB09",
    x"BF53D782",
    x"BF53D3FB",
    x"BF53D074",
    x"BF53CCEC",
    x"BF53C965",
    x"BF53C5DD",
    x"BF53C255",
    x"BF53BECD",
    x"BF53BB45",
    x"BF53B7BD",
    x"BF53B435",
    x"BF53B0AC",
    x"BF53AD24",
    x"BF53A99B",
    x"BF53A612",
    x"BF53A289",
    x"BF539F00",
    x"BF539B77",
    x"BF5397EE",
    x"BF539464",
    x"BF5390DB",
    x"BF538D51",
    x"BF5389C7",
    x"BF53863D",
    x"BF5382B3",
    x"BF537F29",
    x"BF537B9E",
    x"BF537814",
    x"BF537489",
    x"BF5370FF",
    x"BF536D74",
    x"BF5369E9",
    x"BF53665E",
    x"BF5362D2",
    x"BF535F47",
    x"BF535BBB",
    x"BF535830",
    x"BF5354A4",
    x"BF535118",
    x"BF534D8C",
    x"BF534A00",
    x"BF534674",
    x"BF5342E7",
    x"BF533F5B",
    x"BF533BCE",
    x"BF533841",
    x"BF5334B5",
    x"BF533128",
    x"BF532D9A",
    x"BF532A0D",
    x"BF532680",
    x"BF5322F2",
    x"BF531F65",
    x"BF531BD7",
    x"BF531849",
    x"BF5314BB",
    x"BF53112D",
    x"BF530D9E",
    x"BF530A10",
    x"BF530681",
    x"BF5302F3",
    x"BF52FF64",
    x"BF52FBD5",
    x"BF52F846",
    x"BF52F4B7",
    x"BF52F127",
    x"BF52ED98",
    x"BF52EA08",
    x"BF52E679",
    x"BF52E2E9",
    x"BF52DF59",
    x"BF52DBC9",
    x"BF52D839",
    x"BF52D4A8",
    x"BF52D118",
    x"BF52CD87",
    x"BF52C9F7",
    x"BF52C666",
    x"BF52C2D5",
    x"BF52BF44",
    x"BF52BBB2",
    x"BF52B821",
    x"BF52B490",
    x"BF52B0FE",
    x"BF52AD6C",
    x"BF52A9DA",
    x"BF52A649",
    x"BF52A2B6",
    x"BF529F24",
    x"BF529B92",
    x"BF5297FF",
    x"BF52946D",
    x"BF5290DA",
    x"BF528D47",
    x"BF5289B4",
    x"BF528621",
    x"BF52828E",
    x"BF527EFA",
    x"BF527B67",
    x"BF5277D3",
    x"BF52743F",
    x"BF5270AC",
    x"BF526D18",
    x"BF526983",
    x"BF5265EF",
    x"BF52625B",
    x"BF525EC6",
    x"BF525B32",
    x"BF52579D",
    x"BF525408",
    x"BF525073",
    x"BF524CDE",
    x"BF524949",
    x"BF5245B3",
    x"BF52421E",
    x"BF523E88",
    x"BF523AF2",
    x"BF52375C",
    x"BF5233C6",
    x"BF523030",
    x"BF522C9A",
    x"BF522903",
    x"BF52256D",
    x"BF5221D6",
    x"BF521E3F",
    x"BF521AA8",
    x"BF521711",
    x"BF52137A",
    x"BF520FE3",
    x"BF520C4C",
    x"BF5208B4",
    x"BF52051C",
    x"BF520184",
    x"BF51FDED",
    x"BF51FA54",
    x"BF51F6BC",
    x"BF51F324",
    x"BF51EF8C",
    x"BF51EBF3",
    x"BF51E85A",
    x"BF51E4C1",
    x"BF51E129",
    x"BF51DD8F",
    x"BF51D9F6",
    x"BF51D65D",
    x"BF51D2C3",
    x"BF51CF2A",
    x"BF51CB90",
    x"BF51C7F6",
    x"BF51C45C",
    x"BF51C0C2",
    x"BF51BD28",
    x"BF51B98E",
    x"BF51B5F3",
    x"BF51B259",
    x"BF51AEBE",
    x"BF51AB23",
    x"BF51A788",
    x"BF51A3ED",
    x"BF51A052",
    x"BF519CB7",
    x"BF51991B",
    x"BF51957F",
    x"BF5191E4",
    x"BF518E48",
    x"BF518AAC",
    x"BF518710",
    x"BF518374",
    x"BF517FD7",
    x"BF517C3B",
    x"BF51789E",
    x"BF517501",
    x"BF517165",
    x"BF516DC8",
    x"BF516A2A",
    x"BF51668D",
    x"BF5162F0",
    x"BF515F52",
    x"BF515BB5",
    x"BF515817",
    x"BF515479",
    x"BF5150DB",
    x"BF514D3D",
    x"BF51499F",
    x"BF514600",
    x"BF514262",
    x"BF513EC3",
    x"BF513B25",
    x"BF513786",
    x"BF5133E7",
    x"BF513047",
    x"BF512CA8",
    x"BF512909",
    x"BF512569",
    x"BF5121CA",
    x"BF511E2A",
    x"BF511A8A",
    x"BF5116EA",
    x"BF51134A",
    x"BF510FAA",
    x"BF510C09",
    x"BF510869",
    x"BF5104C8",
    x"BF510127",
    x"BF50FD86",
    x"BF50F9E5",
    x"BF50F644",
    x"BF50F2A3",
    x"BF50EF02",
    x"BF50EB60",
    x"BF50E7BE",
    x"BF50E41D",
    x"BF50E07B",
    x"BF50DCD9",
    x"BF50D937",
    x"BF50D594",
    x"BF50D1F2",
    x"BF50CE4F",
    x"BF50CAAD",
    x"BF50C70A",
    x"BF50C367",
    x"BF50BFC4",
    x"BF50BC21",
    x"BF50B87E",
    x"BF50B4DA",
    x"BF50B137",
    x"BF50AD93",
    x"BF50A9EF",
    x"BF50A64B",
    x"BF50A2A7",
    x"BF509F03",
    x"BF509B5F",
    x"BF5097BA",
    x"BF509416",
    x"BF509071",
    x"BF508CCC",
    x"BF508927",
    x"BF508582",
    x"BF5081DD",
    x"BF507E38",
    x"BF507A92",
    x"BF5076ED",
    x"BF507347",
    x"BF506FA1",
    x"BF506BFC",
    x"BF506856",
    x"BF5064AF",
    x"BF506109",
    x"BF505D63",
    x"BF5059BC",
    x"BF505615",
    x"BF50526F",
    x"BF504EC8",
    x"BF504B21",
    x"BF504779",
    x"BF5043D2",
    x"BF50402B",
    x"BF503C83",
    x"BF5038DB",
    x"BF503534",
    x"BF50318C",
    x"BF502DE4",
    x"BF502A3B",
    x"BF502693",
    x"BF5022EB",
    x"BF501F42",
    x"BF501B9A",
    x"BF5017F1",
    x"BF501448",
    x"BF50109F",
    x"BF500CF6",
    x"BF50094C",
    x"BF5005A3",
    x"BF5001F9",
    x"BF4FFE50",
    x"BF4FFAA6",
    x"BF4FF6FC",
    x"BF4FF352",
    x"BF4FEFA8",
    x"BF4FEBFD",
    x"BF4FE853",
    x"BF4FE4A8",
    x"BF4FE0FE",
    x"BF4FDD53",
    x"BF4FD9A8",
    x"BF4FD5FD",
    x"BF4FD252",
    x"BF4FCEA6",
    x"BF4FCAFB",
    x"BF4FC74F",
    x"BF4FC3A4",
    x"BF4FBFF8",
    x"BF4FBC4C",
    x"BF4FB8A0",
    x"BF4FB4F4",
    x"BF4FB147",
    x"BF4FAD9B",
    x"BF4FA9EE",
    x"BF4FA642",
    x"BF4FA295",
    x"BF4F9EE8",
    x"BF4F9B3B",
    x"BF4F978D",
    x"BF4F93E0",
    x"BF4F9033",
    x"BF4F8C85",
    x"BF4F88D7",
    x"BF4F852A",
    x"BF4F817C",
    x"BF4F7DCE",
    x"BF4F7A1F",
    x"BF4F7671",
    x"BF4F72C3",
    x"BF4F6F14",
    x"BF4F6B65",
    x"BF4F67B7",
    x"BF4F6408",
    x"BF4F6059",
    x"BF4F5CA9",
    x"BF4F58FA",
    x"BF4F554B",
    x"BF4F519B",
    x"BF4F4DEB",
    x"BF4F4A3C",
    x"BF4F468C",
    x"BF4F42DC",
    x"BF4F3F2B",
    x"BF4F3B7B",
    x"BF4F37CB",
    x"BF4F341A",
    x"BF4F3069",
    x"BF4F2CB9",
    x"BF4F2908",
    x"BF4F2557",
    x"BF4F21A5",
    x"BF4F1DF4",
    x"BF4F1A43",
    x"BF4F1691",
    x"BF4F12DF",
    x"BF4F0F2E",
    x"BF4F0B7C",
    x"BF4F07CA",
    x"BF4F0417",
    x"BF4F0065",
    x"BF4EFCB3",
    x"BF4EF900",
    x"BF4EF54D",
    x"BF4EF19B",
    x"BF4EEDE8",
    x"BF4EEA35",
    x"BF4EE681",
    x"BF4EE2CE",
    x"BF4EDF1B",
    x"BF4EDB67",
    x"BF4ED7B3",
    x"BF4ED400",
    x"BF4ED04C",
    x"BF4ECC98",
    x"BF4EC8E4",
    x"BF4EC52F",
    x"BF4EC17B",
    x"BF4EBDC6",
    x"BF4EBA12",
    x"BF4EB65D",
    x"BF4EB2A8",
    x"BF4EAEF3",
    x"BF4EAB3E",
    x"BF4EA788",
    x"BF4EA3D3",
    x"BF4EA01D",
    x"BF4E9C68",
    x"BF4E98B2",
    x"BF4E94FC",
    x"BF4E9146",
    x"BF4E8D90",
    x"BF4E89D9",
    x"BF4E8623",
    x"BF4E826C",
    x"BF4E7EB6",
    x"BF4E7AFF",
    x"BF4E7748",
    x"BF4E7391",
    x"BF4E6FDA",
    x"BF4E6C23",
    x"BF4E686B",
    x"BF4E64B4",
    x"BF4E60FC",
    x"BF4E5D44",
    x"BF4E598C",
    x"BF4E55D4",
    x"BF4E521C",
    x"BF4E4E64",
    x"BF4E4AAB",
    x"BF4E46F3",
    x"BF4E433A",
    x"BF4E3F81",
    x"BF4E3BC8",
    x"BF4E380F",
    x"BF4E3456",
    x"BF4E309D",
    x"BF4E2CE4",
    x"BF4E292A",
    x"BF4E2570",
    x"BF4E21B7",
    x"BF4E1DFD",
    x"BF4E1A43",
    x"BF4E1689",
    x"BF4E12CE",
    x"BF4E0F14",
    x"BF4E0B59",
    x"BF4E079F",
    x"BF4E03E4",
    x"BF4E0029",
    x"BF4DFC6E",
    x"BF4DF8B3",
    x"BF4DF4F8",
    x"BF4DF13C",
    x"BF4DED81",
    x"BF4DE9C5",
    x"BF4DE609",
    x"BF4DE24D",
    x"BF4DDE91",
    x"BF4DDAD5",
    x"BF4DD719",
    x"BF4DD35D",
    x"BF4DCFA0",
    x"BF4DCBE3",
    x"BF4DC827",
    x"BF4DC46A",
    x"BF4DC0AD",
    x"BF4DBCF0",
    x"BF4DB932",
    x"BF4DB575",
    x"BF4DB1B8",
    x"BF4DADFA",
    x"BF4DAA3C",
    x"BF4DA67E",
    x"BF4DA2C0",
    x"BF4D9F02",
    x"BF4D9B44",
    x"BF4D9786",
    x"BF4D93C7",
    x"BF4D9009",
    x"BF4D8C4A",
    x"BF4D888B",
    x"BF4D84CC",
    x"BF4D810D",
    x"BF4D7D4E",
    x"BF4D798E",
    x"BF4D75CF",
    x"BF4D720F",
    x"BF4D6E4F",
    x"BF4D6A90",
    x"BF4D66D0",
    x"BF4D6310",
    x"BF4D5F4F",
    x"BF4D5B8F",
    x"BF4D57CE",
    x"BF4D540E",
    x"BF4D504D",
    x"BF4D4C8C",
    x"BF4D48CB",
    x"BF4D450A",
    x"BF4D4149",
    x"BF4D3D88",
    x"BF4D39C6",
    x"BF4D3605",
    x"BF4D3243",
    x"BF4D2E81",
    x"BF4D2ABF",
    x"BF4D26FD",
    x"BF4D233B",
    x"BF4D1F79",
    x"BF4D1BB6",
    x"BF4D17F4",
    x"BF4D1431",
    x"BF4D106E",
    x"BF4D0CAB",
    x"BF4D08E8",
    x"BF4D0525",
    x"BF4D0162",
    x"BF4CFD9E",
    x"BF4CF9DB",
    x"BF4CF617",
    x"BF4CF253",
    x"BF4CEE8F",
    x"BF4CEACB",
    x"BF4CE707",
    x"BF4CE343",
    x"BF4CDF7E",
    x"BF4CDBBA",
    x"BF4CD7F5",
    x"BF4CD430",
    x"BF4CD06B",
    x"BF4CCCA6",
    x"BF4CC8E1",
    x"BF4CC51C",
    x"BF4CC156",
    x"BF4CBD91",
    x"BF4CB9CB",
    x"BF4CB605",
    x"BF4CB23F",
    x"BF4CAE79",
    x"BF4CAAB3",
    x"BF4CA6ED",
    x"BF4CA327",
    x"BF4C9F60",
    x"BF4C9B99",
    x"BF4C97D3",
    x"BF4C940C",
    x"BF4C9045",
    x"BF4C8C7E",
    x"BF4C88B6",
    x"BF4C84EF",
    x"BF4C8128",
    x"BF4C7D60",
    x"BF4C7998",
    x"BF4C75D0",
    x"BF4C7208",
    x"BF4C6E40",
    x"BF4C6A78",
    x"BF4C66B0",
    x"BF4C62E7",
    x"BF4C5F1E",
    x"BF4C5B56",
    x"BF4C578D",
    x"BF4C53C4",
    x"BF4C4FFB",
    x"BF4C4C32",
    x"BF4C4868",
    x"BF4C449F",
    x"BF4C40D5",
    x"BF4C3D0B",
    x"BF4C3942",
    x"BF4C3578",
    x"BF4C31AD",
    x"BF4C2DE3",
    x"BF4C2A19",
    x"BF4C264E",
    x"BF4C2284",
    x"BF4C1EB9",
    x"BF4C1AEE",
    x"BF4C1723",
    x"BF4C1358",
    x"BF4C0F8D",
    x"BF4C0BC2",
    x"BF4C07F6",
    x"BF4C042B",
    x"BF4C005F",
    x"BF4BFC93",
    x"BF4BF8C7",
    x"BF4BF4FB",
    x"BF4BF12F",
    x"BF4BED63",
    x"BF4BE996",
    x"BF4BE5CA",
    x"BF4BE1FD",
    x"BF4BDE30",
    x"BF4BDA63",
    x"BF4BD696",
    x"BF4BD2C9",
    x"BF4BCEFC",
    x"BF4BCB2F",
    x"BF4BC761",
    x"BF4BC393",
    x"BF4BBFC6",
    x"BF4BBBF8",
    x"BF4BB82A",
    x"BF4BB45B",
    x"BF4BB08D",
    x"BF4BACBF",
    x"BF4BA8F0",
    x"BF4BA522",
    x"BF4BA153",
    x"BF4B9D84",
    x"BF4B99B5",
    x"BF4B95E6",
    x"BF4B9217",
    x"BF4B8E47",
    x"BF4B8A78",
    x"BF4B86A8",
    x"BF4B82D8",
    x"BF4B7F09",
    x"BF4B7B39",
    x"BF4B7768",
    x"BF4B7398",
    x"BF4B6FC8",
    x"BF4B6BF7",
    x"BF4B6827",
    x"BF4B6456",
    x"BF4B6085",
    x"BF4B5CB4",
    x"BF4B58E3",
    x"BF4B5512",
    x"BF4B5141",
    x"BF4B4D6F",
    x"BF4B499E",
    x"BF4B45CC",
    x"BF4B41FA",
    x"BF4B3E28",
    x"BF4B3A56",
    x"BF4B3684",
    x"BF4B32B2",
    x"BF4B2EDF",
    x"BF4B2B0D",
    x"BF4B273A",
    x"BF4B2367",
    x"BF4B1F94",
    x"BF4B1BC1",
    x"BF4B17EE",
    x"BF4B141B",
    x"BF4B1047",
    x"BF4B0C74",
    x"BF4B08A0",
    x"BF4B04CC",
    x"BF4B00F8",
    x"BF4AFD24",
    x"BF4AF950",
    x"BF4AF57C",
    x"BF4AF1A8",
    x"BF4AEDD3",
    x"BF4AE9FE",
    x"BF4AE62A",
    x"BF4AE255",
    x"BF4ADE80",
    x"BF4ADAAB",
    x"BF4AD6D5",
    x"BF4AD300",
    x"BF4ACF2A",
    x"BF4ACB55",
    x"BF4AC77F",
    x"BF4AC3A9",
    x"BF4ABFD3",
    x"BF4ABBFD",
    x"BF4AB827",
    x"BF4AB451",
    x"BF4AB07A",
    x"BF4AACA4",
    x"BF4AA8CD",
    x"BF4AA4F6",
    x"BF4AA11F",
    x"BF4A9D48",
    x"BF4A9971",
    x"BF4A9599",
    x"BF4A91C2",
    x"BF4A8DEA",
    x"BF4A8A13",
    x"BF4A863B",
    x"BF4A8263",
    x"BF4A7E8B",
    x"BF4A7AB3",
    x"BF4A76DA",
    x"BF4A7302",
    x"BF4A6F29",
    x"BF4A6B51",
    x"BF4A6778",
    x"BF4A639F",
    x"BF4A5FC6",
    x"BF4A5BED",
    x"BF4A5814",
    x"BF4A543A",
    x"BF4A5061",
    x"BF4A4C87",
    x"BF4A48AD",
    x"BF4A44D3",
    x"BF4A40F9",
    x"BF4A3D1F",
    x"BF4A3945",
    x"BF4A356B",
    x"BF4A3190",
    x"BF4A2DB6",
    x"BF4A29DB",
    x"BF4A2600",
    x"BF4A2225",
    x"BF4A1E4A",
    x"BF4A1A6F",
    x"BF4A1693",
    x"BF4A12B8",
    x"BF4A0EDC",
    x"BF4A0B01",
    x"BF4A0725",
    x"BF4A0349",
    x"BF49FF6D",
    x"BF49FB91",
    x"BF49F7B4",
    x"BF49F3D8",
    x"BF49EFFB",
    x"BF49EC1F",
    x"BF49E842",
    x"BF49E465",
    x"BF49E088",
    x"BF49DCAB",
    x"BF49D8CD",
    x"BF49D4F0",
    x"BF49D112",
    x"BF49CD35",
    x"BF49C957",
    x"BF49C579",
    x"BF49C19B",
    x"BF49BDBD",
    x"BF49B9DF",
    x"BF49B600",
    x"BF49B222",
    x"BF49AE43",
    x"BF49AA64",
    x"BF49A685",
    x"BF49A2A6",
    x"BF499EC7",
    x"BF499AE8",
    x"BF499709",
    x"BF499329",
    x"BF498F4A",
    x"BF498B6A",
    x"BF49878A",
    x"BF4983AA",
    x"BF497FCA",
    x"BF497BEA",
    x"BF497809",
    x"BF497429",
    x"BF497048",
    x"BF496C68",
    x"BF496887",
    x"BF4964A6",
    x"BF4960C5",
    x"BF495CE4",
    x"BF495902",
    x"BF495521",
    x"BF49513F",
    x"BF494D5E",
    x"BF49497C",
    x"BF49459A",
    x"BF4941B8",
    x"BF493DD6",
    x"BF4939F4",
    x"BF493611",
    x"BF49322F",
    x"BF492E4C",
    x"BF492A69",
    x"BF492686",
    x"BF4922A3",
    x"BF491EC0",
    x"BF491ADD",
    x"BF4916FA",
    x"BF491316",
    x"BF490F33",
    x"BF490B4F",
    x"BF49076B",
    x"BF490387",
    x"BF48FFA3",
    x"BF48FBBF",
    x"BF48F7DA",
    x"BF48F3F6",
    x"BF48F011",
    x"BF48EC2D",
    x"BF48E848",
    x"BF48E463",
    x"BF48E07E",
    x"BF48DC99",
    x"BF48D8B3",
    x"BF48D4CE",
    x"BF48D0E9",
    x"BF48CD03",
    x"BF48C91D",
    x"BF48C537",
    x"BF48C151",
    x"BF48BD6B",
    x"BF48B985",
    x"BF48B59E",
    x"BF48B1B8",
    x"BF48ADD1",
    x"BF48A9EA",
    x"BF48A604",
    x"BF48A21D",
    x"BF489E36",
    x"BF489A4E",
    x"BF489667",
    x"BF48927F",
    x"BF488E98",
    x"BF488AB0",
    x"BF4886C8",
    x"BF4882E0",
    x"BF487EF8",
    x"BF487B10",
    x"BF487728",
    x"BF48733F",
    x"BF486F57",
    x"BF486B6E",
    x"BF486785",
    x"BF48639C",
    x"BF485FB3",
    x"BF485BCA",
    x"BF4857E1",
    x"BF4853F7",
    x"BF48500E",
    x"BF484C24",
    x"BF48483A",
    x"BF484451",
    x"BF484067",
    x"BF483C7C",
    x"BF483892",
    x"BF4834A8",
    x"BF4830BD",
    x"BF482CD3",
    x"BF4828E8",
    x"BF4824FD",
    x"BF482112",
    x"BF481D27",
    x"BF48193C",
    x"BF481550",
    x"BF481165",
    x"BF480D79",
    x"BF48098E",
    x"BF4805A2",
    x"BF4801B6",
    x"BF47FDCA",
    x"BF47F9DE",
    x"BF47F5F1",
    x"BF47F205",
    x"BF47EE18",
    x"BF47EA2C",
    x"BF47E63F",
    x"BF47E252",
    x"BF47DE65",
    x"BF47DA78",
    x"BF47D68B",
    x"BF47D29D",
    x"BF47CEB0",
    x"BF47CAC2",
    x"BF47C6D4",
    x"BF47C2E7",
    x"BF47BEF9",
    x"BF47BB0A",
    x"BF47B71C",
    x"BF47B32E",
    x"BF47AF3F",
    x"BF47AB51",
    x"BF47A762",
    x"BF47A373",
    x"BF479F84",
    x"BF479B95",
    x"BF4797A6",
    x"BF4793B7",
    x"BF478FC7",
    x"BF478BD8",
    x"BF4787E8",
    x"BF4783F8",
    x"BF478008",
    x"BF477C18",
    x"BF477828",
    x"BF477438",
    x"BF477048",
    x"BF476C57",
    x"BF476866",
    x"BF476476",
    x"BF476085",
    x"BF475C94",
    x"BF4758A3",
    x"BF4754B2",
    x"BF4750C0",
    x"BF474CCF",
    x"BF4748DD",
    x"BF4744EB",
    x"BF4740FA",
    x"BF473D08",
    x"BF473916",
    x"BF473523",
    x"BF473131",
    x"BF472D3F",
    x"BF47294C",
    x"BF472559",
    x"BF472167",
    x"BF471D74",
    x"BF471981",
    x"BF47158D",
    x"BF47119A",
    x"BF470DA7",
    x"BF4709B3",
    x"BF4705C0",
    x"BF4701CC",
    x"BF46FDD8",
    x"BF46F9E4",
    x"BF46F5F0",
    x"BF46F1FC",
    x"BF46EE07",
    x"BF46EA13",
    x"BF46E61E",
    x"BF46E22A",
    x"BF46DE35",
    x"BF46DA40",
    x"BF46D64B",
    x"BF46D256",
    x"BF46CE60",
    x"BF46CA6B",
    x"BF46C675",
    x"BF46C280",
    x"BF46BE8A",
    x"BF46BA94",
    x"BF46B69E",
    x"BF46B2A8",
    x"BF46AEB1",
    x"BF46AABB",
    x"BF46A6C5",
    x"BF46A2CE",
    x"BF469ED7",
    x"BF469AE0",
    x"BF4696E9",
    x"BF4692F2",
    x"BF468EFB",
    x"BF468B04",
    x"BF46870C",
    x"BF468315",
    x"BF467F1D",
    x"BF467B25",
    x"BF46772D",
    x"BF467335",
    x"BF466F3D",
    x"BF466B45",
    x"BF46674C",
    x"BF466354",
    x"BF465F5B",
    x"BF465B62",
    x"BF465769",
    x"BF465370",
    x"BF464F77",
    x"BF464B7E",
    x"BF464785",
    x"BF46438B",
    x"BF463F91",
    x"BF463B98",
    x"BF46379E",
    x"BF4633A4",
    x"BF462FAA",
    x"BF462BB0",
    x"BF4627B5",
    x"BF4623BB",
    x"BF461FC0",
    x"BF461BC6",
    x"BF4617CB",
    x"BF4613D0",
    x"BF460FD5",
    x"BF460BDA",
    x"BF4607DE",
    x"BF4603E3",
    x"BF45FFE7",
    x"BF45FBEC",
    x"BF45F7F0",
    x"BF45F3F4",
    x"BF45EFF8",
    x"BF45EBFC",
    x"BF45E800",
    x"BF45E403",
    x"BF45E007",
    x"BF45DC0A",
    x"BF45D80E",
    x"BF45D411",
    x"BF45D014",
    x"BF45CC17",
    x"BF45C819",
    x"BF45C41C",
    x"BF45C01F",
    x"BF45BC21",
    x"BF45B824",
    x"BF45B426",
    x"BF45B028",
    x"BF45AC2A",
    x"BF45A82C",
    x"BF45A42D",
    x"BF45A02F",
    x"BF459C31",
    x"BF459832",
    x"BF459433",
    x"BF459034",
    x"BF458C35",
    x"BF458836",
    x"BF458437",
    x"BF458038",
    x"BF457C38",
    x"BF457839",
    x"BF457439",
    x"BF457039",
    x"BF456C39",
    x"BF456839",
    x"BF456439",
    x"BF456039",
    x"BF455C38",
    x"BF455838",
    x"BF455437",
    x"BF455036",
    x"BF454C35",
    x"BF454834",
    x"BF454433",
    x"BF454032",
    x"BF453C31",
    x"BF45382F",
    x"BF45342E",
    x"BF45302C",
    x"BF452C2A",
    x"BF452828",
    x"BF452426",
    x"BF452024",
    x"BF451C22",
    x"BF45181F",
    x"BF45141D",
    x"BF45101A",
    x"BF450C17",
    x"BF450814",
    x"BF450411",
    x"BF45000E",
    x"BF44FC0B",
    x"BF44F807",
    x"BF44F404",
    x"BF44F000",
    x"BF44EBFD",
    x"BF44E7F9",
    x"BF44E3F5",
    x"BF44DFF1",
    x"BF44DBED",
    x"BF44D7E8",
    x"BF44D3E4",
    x"BF44CFDF",
    x"BF44CBDB",
    x"BF44C7D6",
    x"BF44C3D1",
    x"BF44BFCC",
    x"BF44BBC7",
    x"BF44B7C1",
    x"BF44B3BC",
    x"BF44AFB6",
    x"BF44ABB1",
    x"BF44A7AB",
    x"BF44A3A5",
    x"BF449F9F",
    x"BF449B99",
    x"BF449793",
    x"BF44938D",
    x"BF448F86",
    x"BF448B80",
    x"BF448779",
    x"BF448372",
    x"BF447F6B",
    x"BF447B64",
    x"BF44775D",
    x"BF447356",
    x"BF446F4E",
    x"BF446B47",
    x"BF44673F",
    x"BF446337",
    x"BF445F2F",
    x"BF445B27",
    x"BF44571F",
    x"BF445317",
    x"BF444F0F",
    x"BF444B06",
    x"BF4446FE",
    x"BF4442F5",
    x"BF443EEC",
    x"BF443AE3",
    x"BF4436DA",
    x"BF4432D1",
    x"BF442EC8",
    x"BF442ABE",
    x"BF4426B5",
    x"BF4422AB",
    x"BF441EA1",
    x"BF441A97",
    x"BF44168D",
    x"BF441283",
    x"BF440E79",
    x"BF440A6F",
    x"BF440664",
    x"BF44025A",
    x"BF43FE4F",
    x"BF43FA44",
    x"BF43F639",
    x"BF43F22E",
    x"BF43EE23",
    x"BF43EA17",
    x"BF43E60C",
    x"BF43E200",
    x"BF43DDF5",
    x"BF43D9E9",
    x"BF43D5DD",
    x"BF43D1D1",
    x"BF43CDC5",
    x"BF43C9B9",
    x"BF43C5AC",
    x"BF43C1A0",
    x"BF43BD93",
    x"BF43B987",
    x"BF43B57A",
    x"BF43B16D",
    x"BF43AD60",
    x"BF43A953",
    x"BF43A545",
    x"BF43A138",
    x"BF439D2A",
    x"BF43991D",
    x"BF43950F",
    x"BF439101",
    x"BF438CF3",
    x"BF4388E5",
    x"BF4384D6",
    x"BF4380C8",
    x"BF437CBA",
    x"BF4378AB",
    x"BF43749C",
    x"BF43708D",
    x"BF436C7F",
    x"BF43686F",
    x"BF436460",
    x"BF436051",
    x"BF435C41",
    x"BF435832",
    x"BF435422",
    x"BF435012",
    x"BF434C03",
    x"BF4347F3",
    x"BF4343E2",
    x"BF433FD2",
    x"BF433BC2",
    x"BF4337B1",
    x"BF4333A1",
    x"BF432F90",
    x"BF432B7F",
    x"BF43276E",
    x"BF43235D",
    x"BF431F4C",
    x"BF431B3B",
    x"BF431729",
    x"BF431318",
    x"BF430F06",
    x"BF430AF4",
    x"BF4306E2",
    x"BF4302D0",
    x"BF42FEBE",
    x"BF42FAAC",
    x"BF42F69A",
    x"BF42F287",
    x"BF42EE74",
    x"BF42EA62",
    x"BF42E64F",
    x"BF42E23C",
    x"BF42DE29",
    x"BF42DA16",
    x"BF42D602",
    x"BF42D1EF",
    x"BF42CDDB",
    x"BF42C9C8",
    x"BF42C5B4",
    x"BF42C1A0",
    x"BF42BD8C",
    x"BF42B978",
    x"BF42B564",
    x"BF42B14F",
    x"BF42AD3B",
    x"BF42A926",
    x"BF42A511",
    x"BF42A0FD",
    x"BF429CE8",
    x"BF4298D3",
    x"BF4294BD",
    x"BF4290A8",
    x"BF428C93",
    x"BF42887D",
    x"BF428468",
    x"BF428052",
    x"BF427C3C",
    x"BF427826",
    x"BF427410",
    x"BF426FFA",
    x"BF426BE3",
    x"BF4267CD",
    x"BF4263B6",
    x"BF425F9F",
    x"BF425B89",
    x"BF425772",
    x"BF42535B",
    x"BF424F43",
    x"BF424B2C",
    x"BF424715",
    x"BF4242FD",
    x"BF423EE5",
    x"BF423ACE",
    x"BF4236B6",
    x"BF42329E",
    x"BF422E86",
    x"BF422A6E",
    x"BF422655",
    x"BF42223D",
    x"BF421E24",
    x"BF421A0B",
    x"BF4215F3",
    x"BF4211DA",
    x"BF420DC1",
    x"BF4209A7",
    x"BF42058E",
    x"BF420175",
    x"BF41FD5B",
    x"BF41F942",
    x"BF41F528",
    x"BF41F10E",
    x"BF41ECF4",
    x"BF41E8DA",
    x"BF41E4C0",
    x"BF41E0A5",
    x"BF41DC8B",
    x"BF41D870",
    x"BF41D456",
    x"BF41D03B",
    x"BF41CC20",
    x"BF41C805",
    x"BF41C3EA",
    x"BF41BFCF",
    x"BF41BBB3",
    x"BF41B798",
    x"BF41B37C",
    x"BF41AF60",
    x"BF41AB44",
    x"BF41A728",
    x"BF41A30C",
    x"BF419EF0",
    x"BF419AD4",
    x"BF4196B7",
    x"BF41929B",
    x"BF418E7E",
    x"BF418A61",
    x"BF418645",
    x"BF418228",
    x"BF417E0A",
    x"BF4179ED",
    x"BF4175D0",
    x"BF4171B2",
    x"BF416D95",
    x"BF416977",
    x"BF416559",
    x"BF41613B",
    x"BF415D1D",
    x"BF4158FF",
    x"BF4154E1",
    x"BF4150C2",
    x"BF414CA4",
    x"BF414885",
    x"BF414466",
    x"BF414047",
    x"BF413C28",
    x"BF413809",
    x"BF4133EA",
    x"BF412FCB",
    x"BF412BAB",
    x"BF41278C",
    x"BF41236C",
    x"BF411F4C",
    x"BF411B2C",
    x"BF41170C",
    x"BF4112EC",
    x"BF410ECC",
    x"BF410AAB",
    x"BF41068B",
    x"BF41026A",
    x"BF40FE49",
    x"BF40FA29",
    x"BF40F608",
    x"BF40F1E7",
    x"BF40EDC5",
    x"BF40E9A4",
    x"BF40E583",
    x"BF40E161",
    x"BF40DD3F",
    x"BF40D91E",
    x"BF40D4FC",
    x"BF40D0DA",
    x"BF40CCB7",
    x"BF40C895",
    x"BF40C473",
    x"BF40C050",
    x"BF40BC2E",
    x"BF40B80B",
    x"BF40B3E8",
    x"BF40AFC5",
    x"BF40ABA2",
    x"BF40A77F",
    x"BF40A35C",
    x"BF409F38",
    x"BF409B15",
    x"BF4096F1",
    x"BF4092CD",
    x"BF408EA9",
    x"BF408A85",
    x"BF408661",
    x"BF40823D",
    x"BF407E19",
    x"BF4079F4",
    x"BF4075D0",
    x"BF4071AB",
    x"BF406D86",
    x"BF406961",
    x"BF40653C",
    x"BF406117",
    x"BF405CF2",
    x"BF4058CD",
    x"BF4054A7",
    x"BF405081",
    x"BF404C5C",
    x"BF404836",
    x"BF404410",
    x"BF403FEA",
    x"BF403BC4",
    x"BF40379D",
    x"BF403377",
    x"BF402F50",
    x"BF402B2A",
    x"BF402703",
    x"BF4022DC",
    x"BF401EB5",
    x"BF401A8E",
    x"BF401667",
    x"BF40123F",
    x"BF400E18",
    x"BF4009F0",
    x"BF4005C8",
    x"BF4001A1",
    x"BF3FFD79",
    x"BF3FF951",
    x"BF3FF529",
    x"BF3FF100",
    x"BF3FECD8",
    x"BF3FE8AF",
    x"BF3FE487",
    x"BF3FE05E",
    x"BF3FDC35",
    x"BF3FD80C",
    x"BF3FD3E3",
    x"BF3FCFBA",
    x"BF3FCB91",
    x"BF3FC767",
    x"BF3FC33E",
    x"BF3FBF14",
    x"BF3FBAEA",
    x"BF3FB6C0",
    x"BF3FB296",
    x"BF3FAE6C",
    x"BF3FAA42",
    x"BF3FA617",
    x"BF3FA1ED",
    x"BF3F9DC2",
    x"BF3F9998",
    x"BF3F956D",
    x"BF3F9142",
    x"BF3F8D17",
    x"BF3F88EC",
    x"BF3F84C0",
    x"BF3F8095",
    x"BF3F7C6A",
    x"BF3F783E",
    x"BF3F7412",
    x"BF3F6FE6",
    x"BF3F6BBA",
    x"BF3F678E",
    x"BF3F6362",
    x"BF3F5F36",
    x"BF3F5B09",
    x"BF3F56DD",
    x"BF3F52B0",
    x"BF3F4E83",
    x"BF3F4A56",
    x"BF3F4629",
    x"BF3F41FC",
    x"BF3F3DCF",
    x"BF3F39A2",
    x"BF3F3574",
    x"BF3F3147",
    x"BF3F2D19",
    x"BF3F28EB",
    x"BF3F24BD",
    x"BF3F208F",
    x"BF3F1C61",
    x"BF3F1833",
    x"BF3F1404",
    x"BF3F0FD6",
    x"BF3F0BA7",
    x"BF3F0778",
    x"BF3F034A",
    x"BF3EFF1B",
    x"BF3EFAEB",
    x"BF3EF6BC",
    x"BF3EF28D",
    x"BF3EEE5E",
    x"BF3EEA2E",
    x"BF3EE5FE",
    x"BF3EE1CF",
    x"BF3EDD9F",
    x"BF3ED96F",
    x"BF3ED53F",
    x"BF3ED10E",
    x"BF3ECCDE",
    x"BF3EC8AD",
    x"BF3EC47D",
    x"BF3EC04C",
    x"BF3EBC1B",
    x"BF3EB7EA",
    x"BF3EB3B9",
    x"BF3EAF88",
    x"BF3EAB57",
    x"BF3EA726",
    x"BF3EA2F4",
    x"BF3E9EC3",
    x"BF3E9A91",
    x"BF3E965F",
    x"BF3E922D",
    x"BF3E8DFB",
    x"BF3E89C9",
    x"BF3E8596",
    x"BF3E8164",
    x"BF3E7D31",
    x"BF3E78FF",
    x"BF3E74CC",
    x"BF3E7099",
    x"BF3E6C66",
    x"BF3E6833",
    x"BF3E6400",
    x"BF3E5FCD",
    x"BF3E5B99",
    x"BF3E5766",
    x"BF3E5332",
    x"BF3E4EFE",
    x"BF3E4ACA",
    x"BF3E4696",
    x"BF3E4262",
    x"BF3E3E2E",
    x"BF3E39F9",
    x"BF3E35C5",
    x"BF3E3190",
    x"BF3E2D5C",
    x"BF3E2927",
    x"BF3E24F2",
    x"BF3E20BD",
    x"BF3E1C88",
    x"BF3E1852",
    x"BF3E141D",
    x"BF3E0FE7",
    x"BF3E0BB2",
    x"BF3E077C",
    x"BF3E0346",
    x"BF3DFF10",
    x"BF3DFADA",
    x"BF3DF6A4",
    x"BF3DF26E",
    x"BF3DEE37",
    x"BF3DEA01",
    x"BF3DE5CA",
    x"BF3DE193",
    x"BF3DDD5C",
    x"BF3DD925",
    x"BF3DD4EE",
    x"BF3DD0B7",
    x"BF3DCC80",
    x"BF3DC848",
    x"BF3DC411",
    x"BF3DBFD9",
    x"BF3DBBA1",
    x"BF3DB769",
    x"BF3DB331",
    x"BF3DAEF9",
    x"BF3DAAC1",
    x"BF3DA688",
    x"BF3DA250",
    x"BF3D9E17",
    x"BF3D99DF",
    x"BF3D95A6",
    x"BF3D916D",
    x"BF3D8D34",
    x"BF3D88FB",
    x"BF3D84C1",
    x"BF3D8088",
    x"BF3D7C4E",
    x"BF3D7815",
    x"BF3D73DB",
    x"BF3D6FA1",
    x"BF3D6B67",
    x"BF3D672D",
    x"BF3D62F3",
    x"BF3D5EB9",
    x"BF3D5A7E",
    x"BF3D5644",
    x"BF3D5209",
    x"BF3D4DCE",
    x"BF3D4993",
    x"BF3D4558",
    x"BF3D411D",
    x"BF3D3CE2",
    x"BF3D38A7",
    x"BF3D346B",
    x"BF3D3030",
    x"BF3D2BF4",
    x"BF3D27B8",
    x"BF3D237C",
    x"BF3D1F40",
    x"BF3D1B04",
    x"BF3D16C8",
    x"BF3D128C",
    x"BF3D0E4F",
    x"BF3D0A12",
    x"BF3D05D6",
    x"BF3D0199",
    x"BF3CFD5C",
    x"BF3CF91F",
    x"BF3CF4E2",
    x"BF3CF0A5",
    x"BF3CEC67",
    x"BF3CE82A",
    x"BF3CE3EC",
    x"BF3CDFAE",
    x"BF3CDB70",
    x"BF3CD733",
    x"BF3CD2F4",
    x"BF3CCEB6",
    x"BF3CCA78",
    x"BF3CC63A",
    x"BF3CC1FB",
    x"BF3CBDBC",
    x"BF3CB97E",
    x"BF3CB53F",
    x"BF3CB100",
    x"BF3CACC1",
    x"BF3CA881",
    x"BF3CA442",
    x"BF3CA003",
    x"BF3C9BC3",
    x"BF3C9784",
    x"BF3C9344",
    x"BF3C8F04",
    x"BF3C8AC4",
    x"BF3C8684",
    x"BF3C8244",
    x"BF3C7E03",
    x"BF3C79C3",
    x"BF3C7582",
    x"BF3C7141",
    x"BF3C6D01",
    x"BF3C68C0",
    x"BF3C647F",
    x"BF3C603E",
    x"BF3C5BFC",
    x"BF3C57BB",
    x"BF3C5379",
    x"BF3C4F38",
    x"BF3C4AF6",
    x"BF3C46B4",
    x"BF3C4272",
    x"BF3C3E30",
    x"BF3C39EE",
    x"BF3C35AC",
    x"BF3C316A",
    x"BF3C2D27",
    x"BF3C28E4",
    x"BF3C24A2",
    x"BF3C205F",
    x"BF3C1C1C",
    x"BF3C17D9",
    x"BF3C1396",
    x"BF3C0F52",
    x"BF3C0B0F",
    x"BF3C06CB",
    x"BF3C0288",
    x"BF3BFE44",
    x"BF3BFA00",
    x"BF3BF5BC",
    x"BF3BF178",
    x"BF3BED34",
    x"BF3BE8F0",
    x"BF3BE4AB",
    x"BF3BE067",
    x"BF3BDC22",
    x"BF3BD7DD",
    x"BF3BD398",
    x"BF3BCF53",
    x"BF3BCB0E",
    x"BF3BC6C9",
    x"BF3BC284",
    x"BF3BBE3E",
    x"BF3BB9F9",
    x"BF3BB5B3",
    x"BF3BB16D",
    x"BF3BAD27",
    x"BF3BA8E1",
    x"BF3BA49B",
    x"BF3BA055",
    x"BF3B9C0F",
    x"BF3B97C8",
    x"BF3B9382",
    x"BF3B8F3B",
    x"BF3B8AF4",
    x"BF3B86AD",
    x"BF3B8266",
    x"BF3B7E1F",
    x"BF3B79D8",
    x"BF3B7590",
    x"BF3B7149",
    x"BF3B6D01",
    x"BF3B68BA",
    x"BF3B6472",
    x"BF3B602A",
    x"BF3B5BE2",
    x"BF3B579A",
    x"BF3B5351",
    x"BF3B4F09",
    x"BF3B4AC1",
    x"BF3B4678",
    x"BF3B422F",
    x"BF3B3DE6",
    x"BF3B399E",
    x"BF3B3554",
    x"BF3B310B",
    x"BF3B2CC2",
    x"BF3B2879",
    x"BF3B242F",
    x"BF3B1FE5",
    x"BF3B1B9C",
    x"BF3B1752",
    x"BF3B1308",
    x"BF3B0EBE",
    x"BF3B0A74",
    x"BF3B0629",
    x"BF3B01DF",
    x"BF3AFD94",
    x"BF3AF94A",
    x"BF3AF4FF",
    x"BF3AF0B4",
    x"BF3AEC69",
    x"BF3AE81E",
    x"BF3AE3D3",
    x"BF3ADF88",
    x"BF3ADB3C",
    x"BF3AD6F1",
    x"BF3AD2A5",
    x"BF3ACE59",
    x"BF3ACA0D",
    x"BF3AC5C1",
    x"BF3AC175",
    x"BF3ABD29",
    x"BF3AB8DD",
    x"BF3AB490",
    x"BF3AB044",
    x"BF3AABF7",
    x"BF3AA7AA",
    x"BF3AA35D",
    x"BF3A9F10",
    x"BF3A9AC3",
    x"BF3A9676",
    x"BF3A9229",
    x"BF3A8DDB",
    x"BF3A898E",
    x"BF3A8540",
    x"BF3A80F2",
    x"BF3A7CA4",
    x"BF3A7856",
    x"BF3A7408",
    x"BF3A6FBA",
    x"BF3A6B6C",
    x"BF3A671D",
    x"BF3A62CF",
    x"BF3A5E80",
    x"BF3A5A31",
    x"BF3A55E2",
    x"BF3A5193",
    x"BF3A4D44",
    x"BF3A48F5",
    x"BF3A44A6",
    x"BF3A4056",
    x"BF3A3C06",
    x"BF3A37B7",
    x"BF3A3367",
    x"BF3A2F17",
    x"BF3A2AC7",
    x"BF3A2677",
    x"BF3A2227",
    x"BF3A1DD6",
    x"BF3A1986",
    x"BF3A1535",
    x"BF3A10E4",
    x"BF3A0C94",
    x"BF3A0843",
    x"BF3A03F2",
    x"BF39FFA1",
    x"BF39FB4F",
    x"BF39F6FE",
    x"BF39F2AC",
    x"BF39EE5B",
    x"BF39EA09",
    x"BF39E5B7",
    x"BF39E165",
    x"BF39DD13",
    x"BF39D8C1",
    x"BF39D46F",
    x"BF39D01D",
    x"BF39CBCA",
    x"BF39C777",
    x"BF39C325",
    x"BF39BED2",
    x"BF39BA7F",
    x"BF39B62C",
    x"BF39B1D9",
    x"BF39AD85",
    x"BF39A932",
    x"BF39A4DF",
    x"BF39A08B",
    x"BF399C37",
    x"BF3997E3",
    x"BF39938F",
    x"BF398F3B",
    x"BF398AE7",
    x"BF398693",
    x"BF39823E",
    x"BF397DEA",
    x"BF397995",
    x"BF397541",
    x"BF3970EC",
    x"BF396C97",
    x"BF396842",
    x"BF3963ED",
    x"BF395F97",
    x"BF395B42",
    x"BF3956EC",
    x"BF395297",
    x"BF394E41",
    x"BF3949EB",
    x"BF394595",
    x"BF39413F",
    x"BF393CE9",
    x"BF393893",
    x"BF39343C",
    x"BF392FE6",
    x"BF392B8F",
    x"BF392738",
    x"BF3922E1",
    x"BF391E8B",
    x"BF391A33",
    x"BF3915DC",
    x"BF391185",
    x"BF390D2E",
    x"BF3908D6",
    x"BF39047E",
    x"BF390027",
    x"BF38FBCF",
    x"BF38F777",
    x"BF38F31F",
    x"BF38EEC7",
    x"BF38EA6E",
    x"BF38E616",
    x"BF38E1BD",
    x"BF38DD65",
    x"BF38D90C",
    x"BF38D4B3",
    x"BF38D05A",
    x"BF38CC01",
    x"BF38C7A8",
    x"BF38C34F",
    x"BF38BEF5",
    x"BF38BA9C",
    x"BF38B642",
    x"BF38B1E8",
    x"BF38AD8E",
    x"BF38A934",
    x"BF38A4DA",
    x"BF38A080",
    x"BF389C26",
    x"BF3897CB",
    x"BF389371",
    x"BF388F16",
    x"BF388ABB",
    x"BF388661",
    x"BF388206",
    x"BF387DAB",
    x"BF38794F",
    x"BF3874F4",
    x"BF387099",
    x"BF386C3D",
    x"BF3867E1",
    x"BF386386",
    x"BF385F2A",
    x"BF385ACE",
    x"BF385672",
    x"BF385216",
    x"BF384DB9",
    x"BF38495D",
    x"BF384500",
    x"BF3840A4",
    x"BF383C47",
    x"BF3837EA",
    x"BF38338D",
    x"BF382F30",
    x"BF382AD3",
    x"BF382676",
    x"BF382218",
    x"BF381DBB",
    x"BF38195D",
    x"BF3814FF",
    x"BF3810A1",
    x"BF380C43",
    x"BF3807E5",
    x"BF380387",
    x"BF37FF29",
    x"BF37FACA",
    x"BF37F66C",
    x"BF37F20D",
    x"BF37EDAF",
    x"BF37E950",
    x"BF37E4F1",
    x"BF37E092",
    x"BF37DC32",
    x"BF37D7D3",
    x"BF37D374",
    x"BF37CF14",
    x"BF37CAB5",
    x"BF37C655",
    x"BF37C1F5",
    x"BF37BD95",
    x"BF37B935",
    x"BF37B4D5",
    x"BF37B074",
    x"BF37AC14",
    x"BF37A7B4",
    x"BF37A353",
    x"BF379EF2",
    x"BF379A91",
    x"BF379630",
    x"BF3791CF",
    x"BF378D6E",
    x"BF37890D",
    x"BF3784AB",
    x"BF37804A",
    x"BF377BE8",
    x"BF377787",
    x"BF377325",
    x"BF376EC3",
    x"BF376A61",
    x"BF3765FE",
    x"BF37619C",
    x"BF375D3A",
    x"BF3758D7",
    x"BF375475",
    x"BF375012",
    x"BF374BAF",
    x"BF37474C",
    x"BF3742E9",
    x"BF373E86",
    x"BF373A23",
    x"BF3735BF",
    x"BF37315C",
    x"BF372CF8",
    x"BF372894",
    x"BF372431",
    x"BF371FCD",
    x"BF371B69",
    x"BF371704",
    x"BF3712A0",
    x"BF370E3C",
    x"BF3709D7",
    x"BF370573",
    x"BF37010E",
    x"BF36FCA9",
    x"BF36F844",
    x"BF36F3DF",
    x"BF36EF7A",
    x"BF36EB15",
    x"BF36E6AF",
    x"BF36E24A",
    x"BF36DDE4",
    x"BF36D97F",
    x"BF36D519",
    x"BF36D0B3",
    x"BF36CC4D",
    x"BF36C7E7",
    x"BF36C380",
    x"BF36BF1A",
    x"BF36BAB4",
    x"BF36B64D",
    x"BF36B1E6",
    x"BF36AD7F",
    x"BF36A919",
    x"BF36A4B2",
    x"BF36A04A",
    x"BF369BE3",
    x"BF36977C",
    x"BF369314",
    x"BF368EAD",
    x"BF368A45",
    x"BF3685DD",
    x"BF368175",
    x"BF367D0D",
    x"BF3678A5",
    x"BF36743D",
    x"BF366FD5",
    x"BF366B6C",
    x"BF366704",
    x"BF36629B",
    x"BF365E32",
    x"BF3659C9",
    x"BF365560",
    x"BF3650F7",
    x"BF364C8E",
    x"BF364825",
    x"BF3643BB",
    x"BF363F52",
    x"BF363AE8",
    x"BF36367E",
    x"BF363214",
    x"BF362DAA",
    x"BF362940",
    x"BF3624D6",
    x"BF36206C",
    x"BF361C01",
    x"BF361797",
    x"BF36132C",
    x"BF360EC1",
    x"BF360A56",
    x"BF3605EB",
    x"BF360180",
    x"BF35FD15",
    x"BF35F8AA",
    x"BF35F43E",
    x"BF35EFD3",
    x"BF35EB67",
    x"BF35E6FB",
    x"BF35E290",
    x"BF35DE24",
    x"BF35D9B8",
    x"BF35D54B",
    x"BF35D0DF",
    x"BF35CC73",
    x"BF35C806",
    x"BF35C39A",
    x"BF35BF2D",
    x"BF35BAC0",
    x"BF35B653",
    x"BF35B1E6",
    x"BF35AD79",
    x"BF35A90B",
    x"BF35A49E",
    x"BF35A031",
    x"BF359BC3",
    x"BF359755",
    x"BF3592E7",
    x"BF358E79",
    x"BF358A0B",
    x"BF35859D",
    x"BF35812F",
    x"BF357CC1",
    x"BF357852",
    x"BF3573E4",
    x"BF356F75",
    x"BF356B06",
    x"BF356697",
    x"BF356228",
    x"BF355DB9",
    x"BF35594A",
    x"BF3554DA",
    x"BF35506B",
    x"BF354BFB",
    x"BF35478C",
    x"BF35431C",
    x"BF353EAC",
    x"BF353A3C",
    x"BF3535CC",
    x"BF35315C",
    x"BF352CEB",
    x"BF35287B",
    x"BF35240A",
    x"BF351F9A",
    x"BF351B29",
    x"BF3516B8",
    x"BF351247",
    x"BF350DD6",
    x"BF350965",
    x"BF3504F3",
    x"BF350082",
    x"BF34FC10",
    x"BF34F79F",
    x"BF34F32D",
    x"BF34EEBB",
    x"BF34EA49",
    x"BF34E5D7",
    x"BF34E165",
    x"BF34DCF2",
    x"BF34D880",
    x"BF34D40D",
    x"BF34CF9B",
    x"BF34CB28",
    x"BF34C6B5",
    x"BF34C242",
    x"BF34BDCF",
    x"BF34B95C",
    x"BF34B4E9",
    x"BF34B075",
    x"BF34AC02",
    x"BF34A78E",
    x"BF34A31B",
    x"BF349EA7",
    x"BF349A33",
    x"BF3495BF",
    x"BF34914B",
    x"BF348CD6",
    x"BF348862",
    x"BF3483ED",
    x"BF347F79",
    x"BF347B04",
    x"BF34768F",
    x"BF34721A",
    x"BF346DA5",
    x"BF346930",
    x"BF3464BB",
    x"BF346046",
    x"BF345BD0",
    x"BF34575B",
    x"BF3452E5",
    x"BF344E6F",
    x"BF3449F9",
    x"BF344583",
    x"BF34410D",
    x"BF343C97",
    x"BF343821",
    x"BF3433AA",
    x"BF342F34",
    x"BF342ABD",
    x"BF342646",
    x"BF3421CF",
    x"BF341D58",
    x"BF3418E1",
    x"BF34146A",
    x"BF340FF3",
    x"BF340B7B",
    x"BF340704",
    x"BF34028C",
    x"BF33FE14",
    x"BF33F99D",
    x"BF33F525",
    x"BF33F0AD",
    x"BF33EC34",
    x"BF33E7BC",
    x"BF33E344",
    x"BF33DECB",
    x"BF33DA53",
    x"BF33D5DA",
    x"BF33D161",
    x"BF33CCE8",
    x"BF33C86F",
    x"BF33C3F6",
    x"BF33BF7D",
    x"BF33BB03",
    x"BF33B68A",
    x"BF33B210",
    x"BF33AD97",
    x"BF33A91D",
    x"BF33A4A3",
    x"BF33A029",
    x"BF339BAF",
    x"BF339735",
    x"BF3392BA",
    x"BF338E40",
    x"BF3389C5",
    x"BF33854B",
    x"BF3380D0",
    x"BF337C55",
    x"BF3377DA",
    x"BF33735F",
    x"BF336EE4",
    x"BF336A68",
    x"BF3365ED",
    x"BF336171",
    x"BF335CF6",
    x"BF33587A",
    x"BF3353FE",
    x"BF334F82",
    x"BF334B06",
    x"BF33468A",
    x"BF33420E",
    x"BF333D91",
    x"BF333915",
    x"BF333498",
    x"BF33301B",
    x"BF332B9F",
    x"BF332722",
    x"BF3322A5",
    x"BF331E27",
    x"BF3319AA",
    x"BF33152D",
    x"BF3310AF",
    x"BF330C32",
    x"BF3307B4",
    x"BF330336",
    x"BF32FEB8",
    x"BF32FA3A",
    x"BF32F5BC",
    x"BF32F13E",
    x"BF32ECC0",
    x"BF32E841",
    x"BF32E3C3",
    x"BF32DF44",
    x"BF32DAC5",
    x"BF32D646",
    x"BF32D1C7",
    x"BF32CD48",
    x"BF32C8C9",
    x"BF32C44A",
    x"BF32BFCA",
    x"BF32BB4B",
    x"BF32B6CB",
    x"BF32B24C",
    x"BF32ADCC",
    x"BF32A94C",
    x"BF32A4CC",
    x"BF32A04C",
    x"BF329BCB",
    x"BF32974B",
    x"BF3292CA",
    x"BF328E4A",
    x"BF3289C9",
    x"BF328548",
    x"BF3280C7",
    x"BF327C46",
    x"BF3277C5",
    x"BF327344",
    x"BF326EC3",
    x"BF326A41",
    x"BF3265C0",
    x"BF32613E",
    x"BF325CBC",
    x"BF32583A",
    x"BF3253B8",
    x"BF324F36",
    x"BF324AB4",
    x"BF324632",
    x"BF3241AF",
    x"BF323D2D",
    x"BF3238AA",
    x"BF323427",
    x"BF322FA5",
    x"BF322B22",
    x"BF32269E",
    x"BF32221B",
    x"BF321D98",
    x"BF321915",
    x"BF321491",
    x"BF32100E",
    x"BF320B8A",
    x"BF320706",
    x"BF320282",
    x"BF31FDFE",
    x"BF31F97A",
    x"BF31F4F6",
    x"BF31F071",
    x"BF31EBED",
    x"BF31E768",
    x"BF31E2E4",
    x"BF31DE5F",
    x"BF31D9DA",
    x"BF31D555",
    x"BF31D0D0",
    x"BF31CC4B",
    x"BF31C7C5",
    x"BF31C340",
    x"BF31BEBA",
    x"BF31BA35",
    x"BF31B5AF",
    x"BF31B129",
    x"BF31ACA3",
    x"BF31A81D",
    x"BF31A397",
    x"BF319F11",
    x"BF319A8A",
    x"BF319604",
    x"BF31917D",
    x"BF318CF6",
    x"BF318870",
    x"BF3183E9",
    x"BF317F62",
    x"BF317ADB",
    x"BF317653",
    x"BF3171CC",
    x"BF316D44",
    x"BF3168BD",
    x"BF316435",
    x"BF315FAD",
    x"BF315B26",
    x"BF31569E",
    x"BF315215",
    x"BF314D8D",
    x"BF314905",
    x"BF31447D",
    x"BF313FF4",
    x"BF313B6B",
    x"BF3136E3",
    x"BF31325A",
    x"BF312DD1",
    x"BF312948",
    x"BF3124BF",
    x"BF312035",
    x"BF311BAC",
    x"BF311722",
    x"BF311299",
    x"BF310E0F",
    x"BF310985",
    x"BF3104FB",
    x"BF310071",
    x"BF30FBE7",
    x"BF30F75D",
    x"BF30F2D3",
    x"BF30EE48",
    x"BF30E9BE",
    x"BF30E533",
    x"BF30E0A8",
    x"BF30DC1D",
    x"BF30D792",
    x"BF30D307",
    x"BF30CE7C",
    x"BF30C9F1",
    x"BF30C566",
    x"BF30C0DA",
    x"BF30BC4E",
    x"BF30B7C3",
    x"BF30B337",
    x"BF30AEAB",
    x"BF30AA1F",
    x"BF30A593",
    x"BF30A106",
    x"BF309C7A",
    x"BF3097EE",
    x"BF309361",
    x"BF308ED4",
    x"BF308A48",
    x"BF3085BB",
    x"BF30812E",
    x"BF307CA1",
    x"BF307813",
    x"BF307386",
    x"BF306EF9",
    x"BF306A6B",
    x"BF3065DD",
    x"BF306150",
    x"BF305CC2",
    x"BF305834",
    x"BF3053A6",
    x"BF304F18",
    x"BF304A89",
    x"BF3045FB",
    x"BF30416C",
    x"BF303CDE",
    x"BF30384F",
    x"BF3033C0",
    x"BF302F31",
    x"BF302AA2",
    x"BF302613",
    x"BF302184",
    x"BF301CF5",
    x"BF301865",
    x"BF3013D6",
    x"BF300F46",
    x"BF300AB6",
    x"BF300626",
    x"BF300196",
    x"BF2FFD06",
    x"BF2FF876",
    x"BF2FF3E6",
    x"BF2FEF56",
    x"BF2FEAC5",
    x"BF2FE634",
    x"BF2FE1A4",
    x"BF2FDD13",
    x"BF2FD882",
    x"BF2FD3F1",
    x"BF2FCF60",
    x"BF2FCACF",
    x"BF2FC63D",
    x"BF2FC1AC",
    x"BF2FBD1A",
    x"BF2FB888",
    x"BF2FB3F7",
    x"BF2FAF65",
    x"BF2FAAD3",
    x"BF2FA641",
    x"BF2FA1AF",
    x"BF2F9D1C",
    x"BF2F988A",
    x"BF2F93F7",
    x"BF2F8F65",
    x"BF2F8AD2",
    x"BF2F863F",
    x"BF2F81AC",
    x"BF2F7D19",
    x"BF2F7886",
    x"BF2F73F3",
    x"BF2F6F5F",
    x"BF2F6ACC",
    x"BF2F6638",
    x"BF2F61A5",
    x"BF2F5D11",
    x"BF2F587D",
    x"BF2F53E9",
    x"BF2F4F55",
    x"BF2F4AC1",
    x"BF2F462C",
    x"BF2F4198",
    x"BF2F3D03",
    x"BF2F386F",
    x"BF2F33DA",
    x"BF2F2F45",
    x"BF2F2AB0",
    x"BF2F261B",
    x"BF2F2186",
    x"BF2F1CF1",
    x"BF2F185B",
    x"BF2F13C6",
    x"BF2F0F30",
    x"BF2F0A9B",
    x"BF2F0605",
    x"BF2F016F",
    x"BF2EFCD9",
    x"BF2EF843",
    x"BF2EF3AD",
    x"BF2EEF16",
    x"BF2EEA80",
    x"BF2EE5E9",
    x"BF2EE153",
    x"BF2EDCBC",
    x"BF2ED825",
    x"BF2ED38E",
    x"BF2ECEF7",
    x"BF2ECA60",
    x"BF2EC5C9",
    x"BF2EC131",
    x"BF2EBC9A",
    x"BF2EB802",
    x"BF2EB36B",
    x"BF2EAED3",
    x"BF2EAA3B",
    x"BF2EA5A3",
    x"BF2EA10B",
    x"BF2E9C73",
    x"BF2E97DA",
    x"BF2E9342",
    x"BF2E8EA9",
    x"BF2E8A11",
    x"BF2E8578",
    x"BF2E80DF",
    x"BF2E7C46",
    x"BF2E77AD",
    x"BF2E7314",
    x"BF2E6E7B",
    x"BF2E69E1",
    x"BF2E6548",
    x"BF2E60AE",
    x"BF2E5C15",
    x"BF2E577B",
    x"BF2E52E1",
    x"BF2E4E47",
    x"BF2E49AD",
    x"BF2E4513",
    x"BF2E4078",
    x"BF2E3BDE",
    x"BF2E3743",
    x"BF2E32A9",
    x"BF2E2E0E",
    x"BF2E2973",
    x"BF2E24D8",
    x"BF2E203D",
    x"BF2E1BA2",
    x"BF2E1707",
    x"BF2E126B",
    x"BF2E0DD0",
    x"BF2E0934",
    x"BF2E0499",
    x"BF2DFFFD",
    x"BF2DFB61",
    x"BF2DF6C5",
    x"BF2DF229",
    x"BF2DED8D",
    x"BF2DE8F0",
    x"BF2DE454",
    x"BF2DDFB8",
    x"BF2DDB1B",
    x"BF2DD67E",
    x"BF2DD1E1",
    x"BF2DCD44",
    x"BF2DC8A7",
    x"BF2DC40A",
    x"BF2DBF6D",
    x"BF2DBAD0",
    x"BF2DB632",
    x"BF2DB195",
    x"BF2DACF7",
    x"BF2DA859",
    x"BF2DA3BB",
    x"BF2D9F1D",
    x"BF2D9A7F",
    x"BF2D95E1",
    x"BF2D9143",
    x"BF2D8CA4",
    x"BF2D8806",
    x"BF2D8367",
    x"BF2D7EC9",
    x"BF2D7A2A",
    x"BF2D758B",
    x"BF2D70EC",
    x"BF2D6C4D",
    x"BF2D67AD",
    x"BF2D630E",
    x"BF2D5E6F",
    x"BF2D59CF",
    x"BF2D552F",
    x"BF2D5090",
    x"BF2D4BF0",
    x"BF2D4750",
    x"BF2D42B0",
    x"BF2D3E10",
    x"BF2D396F",
    x"BF2D34CF",
    x"BF2D302E",
    x"BF2D2B8E",
    x"BF2D26ED",
    x"BF2D224C",
    x"BF2D1DAB",
    x"BF2D190A",
    x"BF2D1469",
    x"BF2D0FC8",
    x"BF2D0B27",
    x"BF2D0685",
    x"BF2D01E4",
    x"BF2CFD42",
    x"BF2CF8A0",
    x"BF2CF3FF",
    x"BF2CEF5D",
    x"BF2CEABB",
    x"BF2CE618",
    x"BF2CE176",
    x"BF2CDCD4",
    x"BF2CD831",
    x"BF2CD38F",
    x"BF2CCEEC",
    x"BF2CCA49",
    x"BF2CC5A6",
    x"BF2CC103",
    x"BF2CBC60",
    x"BF2CB7BD",
    x"BF2CB31A",
    x"BF2CAE76",
    x"BF2CA9D3",
    x"BF2CA52F",
    x"BF2CA08C",
    x"BF2C9BE8",
    x"BF2C9744",
    x"BF2C92A0",
    x"BF2C8DFC",
    x"BF2C8957",
    x"BF2C84B3",
    x"BF2C800F",
    x"BF2C7B6A",
    x"BF2C76C5",
    x"BF2C7221",
    x"BF2C6D7C",
    x"BF2C68D7",
    x"BF2C6432",
    x"BF2C5F8D",
    x"BF2C5AE7",
    x"BF2C5642",
    x"BF2C519D",
    x"BF2C4CF7",
    x"BF2C4851",
    x"BF2C43AB",
    x"BF2C3F06",
    x"BF2C3A60",
    x"BF2C35B9",
    x"BF2C3113",
    x"BF2C2C6D",
    x"BF2C27C7",
    x"BF2C2320",
    x"BF2C1E79",
    x"BF2C19D3",
    x"BF2C152C",
    x"BF2C1085",
    x"BF2C0BDE",
    x"BF2C0737",
    x"BF2C028F",
    x"BF2BFDE8",
    x"BF2BF941",
    x"BF2BF499",
    x"BF2BEFF1",
    x"BF2BEB4A",
    x"BF2BE6A2",
    x"BF2BE1FA",
    x"BF2BDD52",
    x"BF2BD8AA",
    x"BF2BD401",
    x"BF2BCF59",
    x"BF2BCAB0",
    x"BF2BC608",
    x"BF2BC15F",
    x"BF2BBCB6",
    x"BF2BB80D",
    x"BF2BB364",
    x"BF2BAEBB",
    x"BF2BAA12",
    x"BF2BA569",
    x"BF2BA0BF",
    x"BF2B9C16",
    x"BF2B976C",
    x"BF2B92C2",
    x"BF2B8E19",
    x"BF2B896F",
    x"BF2B84C5",
    x"BF2B801A",
    x"BF2B7B70",
    x"BF2B76C6",
    x"BF2B721B",
    x"BF2B6D71",
    x"BF2B68C6",
    x"BF2B641B",
    x"BF2B5F71",
    x"BF2B5AC6",
    x"BF2B561B",
    x"BF2B516F",
    x"BF2B4CC4",
    x"BF2B4819",
    x"BF2B436D",
    x"BF2B3EC2",
    x"BF2B3A16",
    x"BF2B356A",
    x"BF2B30BE",
    x"BF2B2C12",
    x"BF2B2766",
    x"BF2B22BA",
    x"BF2B1E0E",
    x"BF2B1961",
    x"BF2B14B5",
    x"BF2B1008",
    x"BF2B0B5B",
    x"BF2B06AF",
    x"BF2B0202",
    x"BF2AFD55",
    x"BF2AF8A7",
    x"BF2AF3FA",
    x"BF2AEF4D",
    x"BF2AEA9F",
    x"BF2AE5F2",
    x"BF2AE144",
    x"BF2ADC96",
    x"BF2AD7E9",
    x"BF2AD33B",
    x"BF2ACE8D",
    x"BF2AC9DE",
    x"BF2AC530",
    x"BF2AC082",
    x"BF2ABBD3",
    x"BF2AB725",
    x"BF2AB276",
    x"BF2AADC7",
    x"BF2AA918",
    x"BF2AA469",
    x"BF2A9FBA",
    x"BF2A9B0B",
    x"BF2A965C",
    x"BF2A91AC",
    x"BF2A8CFD",
    x"BF2A884D",
    x"BF2A839E",
    x"BF2A7EEE",
    x"BF2A7A3E",
    x"BF2A758E",
    x"BF2A70DE",
    x"BF2A6C2E",
    x"BF2A677D",
    x"BF2A62CD",
    x"BF2A5E1C",
    x"BF2A596C",
    x"BF2A54BB",
    x"BF2A500A",
    x"BF2A4B59",
    x"BF2A46A8",
    x"BF2A41F7",
    x"BF2A3D46",
    x"BF2A3894",
    x"BF2A33E3",
    x"BF2A2F31",
    x"BF2A2A80",
    x"BF2A25CE",
    x"BF2A211C",
    x"BF2A1C6A",
    x"BF2A17B8",
    x"BF2A1306",
    x"BF2A0E54",
    x"BF2A09A1",
    x"BF2A04EF",
    x"BF2A003C",
    x"BF29FB89",
    x"BF29F6D7",
    x"BF29F224",
    x"BF29ED71",
    x"BF29E8BE",
    x"BF29E40B",
    x"BF29DF57",
    x"BF29DAA4",
    x"BF29D5F0",
    x"BF29D13D",
    x"BF29CC89",
    x"BF29C7D5",
    x"BF29C321",
    x"BF29BE6D",
    x"BF29B9B9",
    x"BF29B505",
    x"BF29B051",
    x"BF29AB9C",
    x"BF29A6E8",
    x"BF29A233",
    x"BF299D7E",
    x"BF2998CA",
    x"BF299415",
    x"BF298F60",
    x"BF298AAA",
    x"BF2985F5",
    x"BF298140",
    x"BF297C8A",
    x"BF2977D5",
    x"BF29731F",
    x"BF296E69",
    x"BF2969B4",
    x"BF2964FE",
    x"BF296048",
    x"BF295B91",
    x"BF2956DB",
    x"BF295225",
    x"BF294D6E",
    x"BF2948B8",
    x"BF294401",
    x"BF293F4A",
    x"BF293A93",
    x"BF2935DD",
    x"BF293125",
    x"BF292C6E",
    x"BF2927B7",
    x"BF292300",
    x"BF291E48",
    x"BF291991",
    x"BF2914D9",
    x"BF291021",
    x"BF290B69",
    x"BF2906B1",
    x"BF2901F9",
    x"BF28FD41",
    x"BF28F889",
    x"BF28F3D0",
    x"BF28EF18",
    x"BF28EA5F",
    x"BF28E5A6",
    x"BF28E0EE",
    x"BF28DC35",
    x"BF28D77C",
    x"BF28D2C3",
    x"BF28CE09",
    x"BF28C950",
    x"BF28C497",
    x"BF28BFDD",
    x"BF28BB23",
    x"BF28B66A",
    x"BF28B1B0",
    x"BF28ACF6",
    x"BF28A83C",
    x"BF28A382",
    x"BF289EC8",
    x"BF289A0D",
    x"BF289553",
    x"BF289098",
    x"BF288BDE",
    x"BF288723",
    x"BF288268",
    x"BF287DAD",
    x"BF2878F2",
    x"BF287437",
    x"BF286F7C",
    x"BF286AC0",
    x"BF286605",
    x"BF286149",
    x"BF285C8E",
    x"BF2857D2",
    x"BF285316",
    x"BF284E5A",
    x"BF28499E",
    x"BF2844E2",
    x"BF284026",
    x"BF283B69",
    x"BF2836AD",
    x"BF2831F0",
    x"BF282D34",
    x"BF282877",
    x"BF2823BA",
    x"BF281EFD",
    x"BF281A40",
    x"BF281583",
    x"BF2810C6",
    x"BF280C08",
    x"BF28074B",
    x"BF28028D",
    x"BF27FDD0",
    x"BF27F912",
    x"BF27F454",
    x"BF27EF96",
    x"BF27EAD8",
    x"BF27E61A",
    x"BF27E15B",
    x"BF27DC9D",
    x"BF27D7DE",
    x"BF27D320",
    x"BF27CE61",
    x"BF27C9A2",
    x"BF27C4E4",
    x"BF27C025",
    x"BF27BB65",
    x"BF27B6A6",
    x"BF27B1E7",
    x"BF27AD28",
    x"BF27A868",
    x"BF27A3A8",
    x"BF279EE9",
    x"BF279A29",
    x"BF279569",
    x"BF2790A9",
    x"BF278BE9",
    x"BF278729",
    x"BF278268",
    x"BF277DA8",
    x"BF2778E8",
    x"BF277427",
    x"BF276F66",
    x"BF276AA5",
    x"BF2765E5",
    x"BF276123",
    x"BF275C62",
    x"BF2757A1",
    x"BF2752E0",
    x"BF274E1E",
    x"BF27495D",
    x"BF27449B",
    x"BF273FDA",
    x"BF273B18",
    x"BF273656",
    x"BF273194",
    x"BF272CD2",
    x"BF272810",
    x"BF27234D",
    x"BF271E8B",
    x"BF2719C8",
    x"BF271506",
    x"BF271043",
    x"BF270B80",
    x"BF2706BD",
    x"BF2701FA",
    x"BF26FD37",
    x"BF26F874",
    x"BF26F3B0",
    x"BF26EEED",
    x"BF26EA2A",
    x"BF26E566",
    x"BF26E0A2",
    x"BF26DBDE",
    x"BF26D71A",
    x"BF26D256",
    x"BF26CD92",
    x"BF26C8CE",
    x"BF26C40A",
    x"BF26BF45",
    x"BF26BA81",
    x"BF26B5BC",
    x"BF26B0F7",
    x"BF26AC33",
    x"BF26A76E",
    x"BF26A2A9",
    x"BF269DE3",
    x"BF26991E",
    x"BF269459",
    x"BF268F93",
    x"BF268ACE",
    x"BF268608",
    x"BF268143",
    x"BF267C7D",
    x"BF2677B7",
    x"BF2672F1",
    x"BF266E2B",
    x"BF266964",
    x"BF26649E",
    x"BF265FD8",
    x"BF265B11",
    x"BF26564A",
    x"BF265184",
    x"BF264CBD",
    x"BF2647F6",
    x"BF26432F",
    x"BF263E68",
    x"BF2639A0",
    x"BF2634D9",
    x"BF263012",
    x"BF262B4A",
    x"BF262682",
    x"BF2621BB",
    x"BF261CF3",
    x"BF26182B",
    x"BF261363",
    x"BF260E9B",
    x"BF2609D3",
    x"BF26050A",
    x"BF260042",
    x"BF25FB79",
    x"BF25F6B1",
    x"BF25F1E8",
    x"BF25ED1F",
    x"BF25E856",
    x"BF25E38D",
    x"BF25DEC4",
    x"BF25D9FB",
    x"BF25D531",
    x"BF25D068",
    x"BF25CB9E",
    x"BF25C6D5",
    x"BF25C20B",
    x"BF25BD41",
    x"BF25B877",
    x"BF25B3AD",
    x"BF25AEE3",
    x"BF25AA19",
    x"BF25A54E",
    x"BF25A084",
    x"BF259BB9",
    x"BF2596EF",
    x"BF259224",
    x"BF258D59",
    x"BF25888E",
    x"BF2583C3",
    x"BF257EF8",
    x"BF257A2D",
    x"BF257562",
    x"BF257096",
    x"BF256BCB",
    x"BF2566FF",
    x"BF256233",
    x"BF255D67",
    x"BF25589B",
    x"BF2553CF",
    x"BF254F03",
    x"BF254A37",
    x"BF25456B",
    x"BF25409E",
    x"BF253BD2",
    x"BF253705",
    x"BF253238",
    x"BF252D6C",
    x"BF25289F",
    x"BF2523D2",
    x"BF251F04",
    x"BF251A37",
    x"BF25156A",
    x"BF25109C",
    x"BF250BCF",
    x"BF250701",
    x"BF250234",
    x"BF24FD66",
    x"BF24F898",
    x"BF24F3CA",
    x"BF24EEFC",
    x"BF24EA2D",
    x"BF24E55F",
    x"BF24E091",
    x"BF24DBC2",
    x"BF24D6F4",
    x"BF24D225",
    x"BF24CD56",
    x"BF24C887",
    x"BF24C3B8",
    x"BF24BEE9",
    x"BF24BA1A",
    x"BF24B54A",
    x"BF24B07B",
    x"BF24ABAC",
    x"BF24A6DC",
    x"BF24A20C",
    x"BF249D3C",
    x"BF24986D",
    x"BF24939C",
    x"BF248ECC",
    x"BF2489FC",
    x"BF24852C",
    x"BF24805B",
    x"BF247B8B",
    x"BF2476BA",
    x"BF2471EA",
    x"BF246D19",
    x"BF246848",
    x"BF246377",
    x"BF245EA6",
    x"BF2459D5",
    x"BF245503",
    x"BF245032",
    x"BF244B60",
    x"BF24468F",
    x"BF2441BD",
    x"BF243CEB",
    x"BF24381A",
    x"BF243348",
    x"BF242E75",
    x"BF2429A3",
    x"BF2424D1",
    x"BF241FFF",
    x"BF241B2C",
    x"BF24165A",
    x"BF241187",
    x"BF240CB4",
    x"BF2407E1",
    x"BF24030E",
    x"BF23FE3B",
    x"BF23F968",
    x"BF23F495",
    x"BF23EFC1",
    x"BF23EAEE",
    x"BF23E61A",
    x"BF23E147",
    x"BF23DC73",
    x"BF23D79F",
    x"BF23D2CB",
    x"BF23CDF7",
    x"BF23C923",
    x"BF23C44F",
    x"BF23BF7A",
    x"BF23BAA6",
    x"BF23B5D1",
    x"BF23B0FC",
    x"BF23AC28",
    x"BF23A753",
    x"BF23A27E",
    x"BF239DA9",
    x"BF2398D4",
    x"BF2393FE",
    x"BF238F29",
    x"BF238A54",
    x"BF23857E",
    x"BF2380A8",
    x"BF237BD3",
    x"BF2376FD",
    x"BF237227",
    x"BF236D51",
    x"BF23687B",
    x"BF2363A5",
    x"BF235ECE",
    x"BF2359F8",
    x"BF235521",
    x"BF23504B",
    x"BF234B74",
    x"BF23469D",
    x"BF2341C6",
    x"BF233CEF",
    x"BF233818",
    x"BF233341",
    x"BF232E6A",
    x"BF232992",
    x"BF2324BB",
    x"BF231FE3",
    x"BF231B0B",
    x"BF231633",
    x"BF23115C",
    x"BF230C84",
    x"BF2307AB",
    x"BF2302D3",
    x"BF22FDFB",
    x"BF22F923",
    x"BF22F44A",
    x"BF22EF72",
    x"BF22EA99",
    x"BF22E5C0",
    x"BF22E0E7",
    x"BF22DC0E",
    x"BF22D735",
    x"BF22D25C",
    x"BF22CD83",
    x"BF22C8A9",
    x"BF22C3D0",
    x"BF22BEF6",
    x"BF22BA1D",
    x"BF22B543",
    x"BF22B069",
    x"BF22AB8F",
    x"BF22A6B5",
    x"BF22A1DB",
    x"BF229D00",
    x"BF229826",
    x"BF22934C",
    x"BF228E71",
    x"BF228996",
    x"BF2284BC",
    x"BF227FE1",
    x"BF227B06",
    x"BF22762B",
    x"BF227150",
    x"BF226C74",
    x"BF226799",
    x"BF2262BE",
    x"BF225DE2",
    x"BF225907",
    x"BF22542B",
    x"BF224F4F",
    x"BF224A73",
    x"BF224597",
    x"BF2240BB",
    x"BF223BDF",
    x"BF223702",
    x"BF223226",
    x"BF222D4A",
    x"BF22286D",
    x"BF222390",
    x"BF221EB3",
    x"BF2219D7",
    x"BF2214FA",
    x"BF22101C",
    x"BF220B3F",
    x"BF220662",
    x"BF220185",
    x"BF21FCA7",
    x"BF21F7C9",
    x"BF21F2EC",
    x"BF21EE0E",
    x"BF21E930",
    x"BF21E452",
    x"BF21DF74",
    x"BF21DA96",
    x"BF21D5B8",
    x"BF21D0D9",
    x"BF21CBFB",
    x"BF21C71C",
    x"BF21C23E",
    x"BF21BD5F",
    x"BF21B880",
    x"BF21B3A1",
    x"BF21AEC2",
    x"BF21A9E3",
    x"BF21A504",
    x"BF21A024",
    x"BF219B45",
    x"BF219665",
    x"BF219186",
    x"BF218CA6",
    x"BF2187C6",
    x"BF2182E6",
    x"BF217E06",
    x"BF217926",
    x"BF217446",
    x"BF216F66",
    x"BF216A85",
    x"BF2165A5",
    x"BF2160C4",
    x"BF215BE3",
    x"BF215703",
    x"BF215222",
    x"BF214D41",
    x"BF214860",
    x"BF21437E",
    x"BF213E9D",
    x"BF2139BC",
    x"BF2134DA",
    x"BF212FF9",
    x"BF212B17",
    x"BF212635",
    x"BF212153",
    x"BF211C71",
    x"BF21178F",
    x"BF2112AD",
    x"BF210DCB",
    x"BF2108E9",
    x"BF210406",
    x"BF20FF24",
    x"BF20FA41",
    x"BF20F55E",
    x"BF20F07B",
    x"BF20EB99",
    x"BF20E6B5",
    x"BF20E1D2",
    x"BF20DCEF",
    x"BF20D80C",
    x"BF20D328",
    x"BF20CE45",
    x"BF20C961",
    x"BF20C47E",
    x"BF20BF9A",
    x"BF20BAB6",
    x"BF20B5D2",
    x"BF20B0EE",
    x"BF20AC0A",
    x"BF20A725",
    x"BF20A241",
    x"BF209D5C",
    x"BF209878",
    x"BF209393",
    x"BF208EAE",
    x"BF2089CA",
    x"BF2084E5",
    x"BF208000",
    x"BF207B1A",
    x"BF207635",
    x"BF207150",
    x"BF206C6A",
    x"BF206785",
    x"BF20629F",
    x"BF205DB9",
    x"BF2058D4",
    x"BF2053EE",
    x"BF204F08",
    x"BF204A21",
    x"BF20453B",
    x"BF204055",
    x"BF203B6F",
    x"BF203688",
    x"BF2031A1",
    x"BF202CBB",
    x"BF2027D4",
    x"BF2022ED",
    x"BF201E06",
    x"BF20191F",
    x"BF201438",
    x"BF200F50",
    x"BF200A69",
    x"BF200582",
    x"BF20009A",
    x"BF1FFBB2",
    x"BF1FF6CB",
    x"BF1FF1E3",
    x"BF1FECFB",
    x"BF1FE813",
    x"BF1FE32B",
    x"BF1FDE42",
    x"BF1FD95A",
    x"BF1FD472",
    x"BF1FCF89",
    x"BF1FCAA0",
    x"BF1FC5B8",
    x"BF1FC0CF",
    x"BF1FBBE6",
    x"BF1FB6FD",
    x"BF1FB214",
    x"BF1FAD2B",
    x"BF1FA841",
    x"BF1FA358",
    x"BF1F9E6E",
    x"BF1F9985",
    x"BF1F949B",
    x"BF1F8FB1",
    x"BF1F8AC7",
    x"BF1F85DD",
    x"BF1F80F3",
    x"BF1F7C09",
    x"BF1F771F",
    x"BF1F7235",
    x"BF1F6D4A",
    x"BF1F6860",
    x"BF1F6375",
    x"BF1F5E8A",
    x"BF1F599F",
    x"BF1F54B4",
    x"BF1F4FC9",
    x"BF1F4ADE",
    x"BF1F45F3",
    x"BF1F4108",
    x"BF1F3C1C",
    x"BF1F3731",
    x"BF1F3245",
    x"BF1F2D59",
    x"BF1F286E",
    x"BF1F2382",
    x"BF1F1E96",
    x"BF1F19AA",
    x"BF1F14BD",
    x"BF1F0FD1",
    x"BF1F0AE5",
    x"BF1F05F8",
    x"BF1F010C",
    x"BF1EFC1F",
    x"BF1EF732",
    x"BF1EF245",
    x"BF1EED59",
    x"BF1EE86C",
    x"BF1EE37E",
    x"BF1EDE91",
    x"BF1ED9A4",
    x"BF1ED4B6",
    x"BF1ECFC9",
    x"BF1ECADB",
    x"BF1EC5ED",
    x"BF1EC100",
    x"BF1EBC12",
    x"BF1EB724",
    x"BF1EB236",
    x"BF1EAD47",
    x"BF1EA859",
    x"BF1EA36B",
    x"BF1E9E7C",
    x"BF1E998E",
    x"BF1E949F",
    x"BF1E8FB0",
    x"BF1E8AC1",
    x"BF1E85D2",
    x"BF1E80E3",
    x"BF1E7BF4",
    x"BF1E7705",
    x"BF1E7216",
    x"BF1E6D26",
    x"BF1E6837",
    x"BF1E6347",
    x"BF1E5E57",
    x"BF1E5968",
    x"BF1E5478",
    x"BF1E4F88",
    x"BF1E4A98",
    x"BF1E45A7",
    x"BF1E40B7",
    x"BF1E3BC7",
    x"BF1E36D6",
    x"BF1E31E6",
    x"BF1E2CF5",
    x"BF1E2804",
    x"BF1E2313",
    x"BF1E1E22",
    x"BF1E1931",
    x"BF1E1440",
    x"BF1E0F4F",
    x"BF1E0A5D",
    x"BF1E056C",
    x"BF1E007B",
    x"BF1DFB89",
    x"BF1DF697",
    x"BF1DF1A5",
    x"BF1DECB3",
    x"BF1DE7C1",
    x"BF1DE2CF",
    x"BF1DDDDD",
    x"BF1DD8EB",
    x"BF1DD3F8",
    x"BF1DCF06",
    x"BF1DCA13",
    x"BF1DC521",
    x"BF1DC02E",
    x"BF1DBB3B",
    x"BF1DB648",
    x"BF1DB155",
    x"BF1DAC62",
    x"BF1DA76F",
    x"BF1DA27B",
    x"BF1D9D88",
    x"BF1D9894",
    x"BF1D93A1",
    x"BF1D8EAD",
    x"BF1D89B9",
    x"BF1D84C5",
    x"BF1D7FD1",
    x"BF1D7ADD",
    x"BF1D75E9",
    x"BF1D70F5",
    x"BF1D6C00",
    x"BF1D670C",
    x"BF1D6217",
    x"BF1D5D23",
    x"BF1D582E",
    x"BF1D5339",
    x"BF1D4E44",
    x"BF1D494F",
    x"BF1D445A",
    x"BF1D3F65",
    x"BF1D3A6F",
    x"BF1D357A",
    x"BF1D3084",
    x"BF1D2B8F",
    x"BF1D2699",
    x"BF1D21A3",
    x"BF1D1CAD",
    x"BF1D17B7",
    x"BF1D12C1",
    x"BF1D0DCB",
    x"BF1D08D5",
    x"BF1D03DE",
    x"BF1CFEE8",
    x"BF1CF9F1",
    x"BF1CF4FB",
    x"BF1CF004",
    x"BF1CEB0D",
    x"BF1CE616",
    x"BF1CE11F",
    x"BF1CDC28",
    x"BF1CD731",
    x"BF1CD239",
    x"BF1CCD42",
    x"BF1CC84B",
    x"BF1CC353",
    x"BF1CBE5B",
    x"BF1CB963",
    x"BF1CB46C",
    x"BF1CAF74",
    x"BF1CAA7C",
    x"BF1CA583",
    x"BF1CA08B",
    x"BF1C9B93",
    x"BF1C969A",
    x"BF1C91A2",
    x"BF1C8CA9",
    x"BF1C87B0",
    x"BF1C82B8",
    x"BF1C7DBF",
    x"BF1C78C6",
    x"BF1C73CC",
    x"BF1C6ED3",
    x"BF1C69DA",
    x"BF1C64E1",
    x"BF1C5FE7",
    x"BF1C5AEE",
    x"BF1C55F4",
    x"BF1C50FA",
    x"BF1C4C00",
    x"BF1C4706",
    x"BF1C420C",
    x"BF1C3D12",
    x"BF1C3818",
    x"BF1C331D",
    x"BF1C2E23",
    x"BF1C2929",
    x"BF1C242E",
    x"BF1C1F33",
    x"BF1C1A38",
    x"BF1C153D",
    x"BF1C1042",
    x"BF1C0B47",
    x"BF1C064C",
    x"BF1C0151",
    x"BF1BFC56",
    x"BF1BF75A",
    x"BF1BF25F",
    x"BF1BED63",
    x"BF1BE867",
    x"BF1BE36B",
    x"BF1BDE6F",
    x"BF1BD973",
    x"BF1BD477",
    x"BF1BCF7B",
    x"BF1BCA7F",
    x"BF1BC582",
    x"BF1BC086",
    x"BF1BBB89",
    x"BF1BB68D",
    x"BF1BB190",
    x"BF1BAC93",
    x"BF1BA796",
    x"BF1BA299",
    x"BF1B9D9C",
    x"BF1B989E",
    x"BF1B93A1",
    x"BF1B8EA4",
    x"BF1B89A6",
    x"BF1B84A9",
    x"BF1B7FAB",
    x"BF1B7AAD",
    x"BF1B75AF",
    x"BF1B70B1",
    x"BF1B6BB3",
    x"BF1B66B5",
    x"BF1B61B7",
    x"BF1B5CB8",
    x"BF1B57BA",
    x"BF1B52BB",
    x"BF1B4DBD",
    x"BF1B48BE",
    x"BF1B43BF",
    x"BF1B3EC0",
    x"BF1B39C1",
    x"BF1B34C2",
    x"BF1B2FC3",
    x"BF1B2AC3",
    x"BF1B25C4",
    x"BF1B20C4",
    x"BF1B1BC5",
    x"BF1B16C5",
    x"BF1B11C5",
    x"BF1B0CC6",
    x"BF1B07C6",
    x"BF1B02C6",
    x"BF1AFDC5",
    x"BF1AF8C5",
    x"BF1AF3C5",
    x"BF1AEEC4",
    x"BF1AE9C4",
    x"BF1AE4C3",
    x"BF1ADFC3",
    x"BF1ADAC2",
    x"BF1AD5C1",
    x"BF1AD0C0",
    x"BF1ACBBF",
    x"BF1AC6BE",
    x"BF1AC1BC",
    x"BF1ABCBB",
    x"BF1AB7BA",
    x"BF1AB2B8",
    x"BF1AADB6",
    x"BF1AA8B5",
    x"BF1AA3B3",
    x"BF1A9EB1",
    x"BF1A99AF",
    x"BF1A94AD",
    x"BF1A8FAB",
    x"BF1A8AA8",
    x"BF1A85A6",
    x"BF1A80A3",
    x"BF1A7BA1",
    x"BF1A769E",
    x"BF1A719B",
    x"BF1A6C99",
    x"BF1A6796",
    x"BF1A6293",
    x"BF1A5D8F",
    x"BF1A588C",
    x"BF1A5389",
    x"BF1A4E86",
    x"BF1A4982",
    x"BF1A447E",
    x"BF1A3F7B",
    x"BF1A3A77",
    x"BF1A3573",
    x"BF1A306F",
    x"BF1A2B6B",
    x"BF1A2667",
    x"BF1A2163",
    x"BF1A1C5E",
    x"BF1A175A",
    x"BF1A1255",
    x"BF1A0D51",
    x"BF1A084C",
    x"BF1A0347",
    x"BF19FE42",
    x"BF19F93D",
    x"BF19F438",
    x"BF19EF33",
    x"BF19EA2E",
    x"BF19E529",
    x"BF19E023",
    x"BF19DB1E",
    x"BF19D618",
    x"BF19D112",
    x"BF19CC0C",
    x"BF19C706",
    x"BF19C200",
    x"BF19BCFA",
    x"BF19B7F4",
    x"BF19B2EE",
    x"BF19ADE7",
    x"BF19A8E1",
    x"BF19A3DA",
    x"BF199ED4",
    x"BF1999CD",
    x"BF1994C6",
    x"BF198FBF",
    x"BF198AB8",
    x"BF1985B1",
    x"BF1980AA",
    x"BF197BA3",
    x"BF19769B",
    x"BF197194",
    x"BF196C8C",
    x"BF196784",
    x"BF19627D",
    x"BF195D75",
    x"BF19586D",
    x"BF195365",
    x"BF194E5D",
    x"BF194955",
    x"BF19444C",
    x"BF193F44",
    x"BF193A3B",
    x"BF193533",
    x"BF19302A",
    x"BF192B21",
    x"BF192618",
    x"BF19210F",
    x"BF191C06",
    x"BF1916FD",
    x"BF1911F4",
    x"BF190CEB",
    x"BF1907E1",
    x"BF1902D8",
    x"BF18FDCE",
    x"BF18F8C4",
    x"BF18F3BB",
    x"BF18EEB1",
    x"BF18E9A7",
    x"BF18E49D",
    x"BF18DF92",
    x"BF18DA88",
    x"BF18D57E",
    x"BF18D073",
    x"BF18CB69",
    x"BF18C65E",
    x"BF18C154",
    x"BF18BC49",
    x"BF18B73E",
    x"BF18B233",
    x"BF18AD28",
    x"BF18A81D",
    x"BF18A311",
    x"BF189E06",
    x"BF1898FB",
    x"BF1893EF",
    x"BF188EE3",
    x"BF1889D8",
    x"BF1884CC",
    x"BF187FC0",
    x"BF187AB4",
    x"BF1875A8",
    x"BF18709C",
    x"BF186B8F",
    x"BF186683",
    x"BF186177",
    x"BF185C6A",
    x"BF18575D",
    x"BF185251",
    x"BF184D44",
    x"BF184837",
    x"BF18432A",
    x"BF183E1D",
    x"BF183910",
    x"BF183402",
    x"BF182EF5",
    x"BF1829E7",
    x"BF1824DA",
    x"BF181FCC",
    x"BF181ABE",
    x"BF1815B1",
    x"BF1810A3",
    x"BF180B95",
    x"BF180687",
    x"BF180178",
    x"BF17FC6A",
    x"BF17F75C",
    x"BF17F24D",
    x"BF17ED3F",
    x"BF17E830",
    x"BF17E321",
    x"BF17DE12",
    x"BF17D903",
    x"BF17D3F4",
    x"BF17CEE5",
    x"BF17C9D6",
    x"BF17C4C7",
    x"BF17BFB7",
    x"BF17BAA8",
    x"BF17B598",
    x"BF17B089",
    x"BF17AB79",
    x"BF17A669",
    x"BF17A159",
    x"BF179C49",
    x"BF179739",
    x"BF179229",
    x"BF178D18",
    x"BF178808",
    x"BF1782F8",
    x"BF177DE7",
    x"BF1778D6",
    x"BF1773C6",
    x"BF176EB5",
    x"BF1769A4",
    x"BF176493",
    x"BF175F82",
    x"BF175A70",
    x"BF17555F",
    x"BF17504E",
    x"BF174B3C",
    x"BF17462B",
    x"BF174119",
    x"BF173C07",
    x"BF1736F5",
    x"BF1731E3",
    x"BF172CD1",
    x"BF1727BF",
    x"BF1722AD",
    x"BF171D9B",
    x"BF171888",
    x"BF171376",
    x"BF170E63",
    x"BF170950",
    x"BF17043E",
    x"BF16FF2B",
    x"BF16FA18",
    x"BF16F505",
    x"BF16EFF2",
    x"BF16EADE",
    x"BF16E5CB",
    x"BF16E0B8",
    x"BF16DBA4",
    x"BF16D691",
    x"BF16D17D",
    x"BF16CC69",
    x"BF16C755",
    x"BF16C241",
    x"BF16BD2D",
    x"BF16B819",
    x"BF16B305",
    x"BF16ADF1",
    x"BF16A8DC",
    x"BF16A3C8",
    x"BF169EB3",
    x"BF16999F",
    x"BF16948A",
    x"BF168F75",
    x"BF168A60",
    x"BF16854B",
    x"BF168036",
    x"BF167B21",
    x"BF16760B",
    x"BF1670F6",
    x"BF166BE0",
    x"BF1666CB",
    x"BF1661B5",
    x"BF165C9F",
    x"BF16578A",
    x"BF165274",
    x"BF164D5E",
    x"BF164847",
    x"BF164331",
    x"BF163E1B",
    x"BF163905",
    x"BF1633EE",
    x"BF162ED8",
    x"BF1629C1",
    x"BF1624AA",
    x"BF161F93",
    x"BF161A7C",
    x"BF161565",
    x"BF16104E",
    x"BF160B37",
    x"BF160620",
    x"BF160108",
    x"BF15FBF1",
    x"BF15F6D9",
    x"BF15F1C2",
    x"BF15ECAA",
    x"BF15E792",
    x"BF15E27A",
    x"BF15DD62",
    x"BF15D84A",
    x"BF15D332",
    x"BF15CE19",
    x"BF15C901",
    x"BF15C3E9",
    x"BF15BED0",
    x"BF15B9B7",
    x"BF15B49F",
    x"BF15AF86",
    x"BF15AA6D",
    x"BF15A554",
    x"BF15A03B",
    x"BF159B21",
    x"BF159608",
    x"BF1590EF",
    x"BF158BD5",
    x"BF1586BC",
    x"BF1581A2",
    x"BF157C88",
    x"BF15776F",
    x"BF157255",
    x"BF156D3B",
    x"BF156821",
    x"BF156306",
    x"BF155DEC",
    x"BF1558D2",
    x"BF1553B7",
    x"BF154E9D",
    x"BF154982",
    x"BF154467",
    x"BF153F4D",
    x"BF153A32",
    x"BF153517",
    x"BF152FFC",
    x"BF152AE0",
    x"BF1525C5",
    x"BF1520AA",
    x"BF151B8E",
    x"BF151673",
    x"BF151157",
    x"BF150C3B",
    x"BF150720",
    x"BF150204",
    x"BF14FCE8",
    x"BF14F7CC",
    x"BF14F2B0",
    x"BF14ED93",
    x"BF14E877",
    x"BF14E35A",
    x"BF14DE3E",
    x"BF14D921",
    x"BF14D405",
    x"BF14CEE8",
    x"BF14C9CB",
    x"BF14C4AE",
    x"BF14BF91",
    x"BF14BA74",
    x"BF14B557",
    x"BF14B039",
    x"BF14AB1C",
    x"BF14A5FE",
    x"BF14A0E1",
    x"BF149BC3",
    x"BF1496A5",
    x"BF149187",
    x"BF148C69",
    x"BF14874B",
    x"BF14822D",
    x"BF147D0F",
    x"BF1477F1",
    x"BF1472D2",
    x"BF146DB4",
    x"BF146895",
    x"BF146377",
    x"BF145E58",
    x"BF145939",
    x"BF14541A",
    x"BF144EFB",
    x"BF1449DC",
    x"BF1444BD",
    x"BF143F9D",
    x"BF143A7E",
    x"BF14355E",
    x"BF14303F",
    x"BF142B1F",
    x"BF142600",
    x"BF1420E0",
    x"BF141BC0",
    x"BF1416A0",
    x"BF141180",
    x"BF140C5F",
    x"BF14073F",
    x"BF14021F",
    x"BF13FCFE",
    x"BF13F7DE",
    x"BF13F2BD",
    x"BF13ED9C",
    x"BF13E87C",
    x"BF13E35B",
    x"BF13DE3A",
    x"BF13D919",
    x"BF13D3F8",
    x"BF13CED6",
    x"BF13C9B5",
    x"BF13C493",
    x"BF13BF72",
    x"BF13BA50",
    x"BF13B52F",
    x"BF13B00D",
    x"BF13AAEB",
    x"BF13A5C9",
    x"BF13A0A7",
    x"BF139B85",
    x"BF139663",
    x"BF139140",
    x"BF138C1E",
    x"BF1386FB",
    x"BF1381D9",
    x"BF137CB6",
    x"BF137793",
    x"BF137270",
    x"BF136D4D",
    x"BF13682A",
    x"BF136307",
    x"BF135DE4",
    x"BF1358C1",
    x"BF13539D",
    x"BF134E7A",
    x"BF134956",
    x"BF134433",
    x"BF133F0F",
    x"BF1339EB",
    x"BF1334C7",
    x"BF132FA3",
    x"BF132A7F",
    x"BF13255B",
    x"BF132037",
    x"BF131B12",
    x"BF1315EE",
    x"BF1310C9",
    x"BF130BA5",
    x"BF130680",
    x"BF13015B",
    x"BF12FC36",
    x"BF12F711",
    x"BF12F1EC",
    x"BF12ECC7",
    x"BF12E7A2",
    x"BF12E27C",
    x"BF12DD57",
    x"BF12D831",
    x"BF12D30C",
    x"BF12CDE6",
    x"BF12C8C0",
    x"BF12C39A",
    x"BF12BE74",
    x"BF12B94E",
    x"BF12B428",
    x"BF12AF02",
    x"BF12A9DC",
    x"BF12A4B5",
    x"BF129F8F",
    x"BF129A68",
    x"BF129542",
    x"BF12901B",
    x"BF128AF4",
    x"BF1285CD",
    x"BF1280A6",
    x"BF127B7F",
    x"BF127658",
    x"BF127130",
    x"BF126C09",
    x"BF1266E2",
    x"BF1261BA",
    x"BF125C92",
    x"BF12576B",
    x"BF125243",
    x"BF124D1B",
    x"BF1247F3",
    x"BF1242CB",
    x"BF123DA3",
    x"BF12387A",
    x"BF123352",
    x"BF122E2A",
    x"BF122901",
    x"BF1223D9",
    x"BF121EB0",
    x"BF121987",
    x"BF12145E",
    x"BF120F35",
    x"BF120A0C",
    x"BF1204E3",
    x"BF11FFBA",
    x"BF11FA91",
    x"BF11F567",
    x"BF11F03E",
    x"BF11EB14",
    x"BF11E5EA",
    x"BF11E0C1",
    x"BF11DB97",
    x"BF11D66D",
    x"BF11D143",
    x"BF11CC19",
    x"BF11C6EF",
    x"BF11C1C4",
    x"BF11BC9A",
    x"BF11B76F",
    x"BF11B245",
    x"BF11AD1A",
    x"BF11A7F0",
    x"BF11A2C5",
    x"BF119D9A",
    x"BF11986F",
    x"BF119344",
    x"BF118E19",
    x"BF1188ED",
    x"BF1183C2",
    x"BF117E97",
    x"BF11796B",
    x"BF117440",
    x"BF116F14",
    x"BF1169E8",
    x"BF1164BC",
    x"BF115F90",
    x"BF115A64",
    x"BF115538",
    x"BF11500C",
    x"BF114AE0",
    x"BF1145B3",
    x"BF114087",
    x"BF113B5A",
    x"BF11362E",
    x"BF113101",
    x"BF112BD4",
    x"BF1126A7",
    x"BF11217A",
    x"BF111C4D",
    x"BF111720",
    x"BF1111F3",
    x"BF110CC5",
    x"BF110798",
    x"BF11026A",
    x"BF10FD3D",
    x"BF10F80F",
    x"BF10F2E1",
    x"BF10EDB3",
    x"BF10E885",
    x"BF10E357",
    x"BF10DE29",
    x"BF10D8FB",
    x"BF10D3CD",
    x"BF10CE9E",
    x"BF10C970",
    x"BF10C441",
    x"BF10BF13",
    x"BF10B9E4",
    x"BF10B4B5",
    x"BF10AF86",
    x"BF10AA57",
    x"BF10A528",
    x"BF109FF9",
    x"BF109ACA",
    x"BF10959A",
    x"BF10906B",
    x"BF108B3B",
    x"BF10860C",
    x"BF1080DC",
    x"BF107BAC",
    x"BF10767C",
    x"BF10714C",
    x"BF106C1C",
    x"BF1066EC",
    x"BF1061BC",
    x"BF105C8C",
    x"BF10575B",
    x"BF10522B",
    x"BF104CFA",
    x"BF1047CA",
    x"BF104299",
    x"BF103D68",
    x"BF103837",
    x"BF103306",
    x"BF102DD5",
    x"BF1028A4",
    x"BF102373",
    x"BF101E41",
    x"BF101910",
    x"BF1013DE",
    x"BF100EAD",
    x"BF10097B",
    x"BF100449",
    x"BF0FFF17",
    x"BF0FF9E5",
    x"BF0FF4B3",
    x"BF0FEF81",
    x"BF0FEA4F",
    x"BF0FE51D",
    x"BF0FDFEA",
    x"BF0FDAB8",
    x"BF0FD585",
    x"BF0FD053",
    x"BF0FCB20",
    x"BF0FC5ED",
    x"BF0FC0BA",
    x"BF0FBB87",
    x"BF0FB654",
    x"BF0FB121",
    x"BF0FABEE",
    x"BF0FA6BA",
    x"BF0FA187",
    x"BF0F9C53",
    x"BF0F9720",
    x"BF0F91EC",
    x"BF0F8CB8",
    x"BF0F8784",
    x"BF0F8250",
    x"BF0F7D1C",
    x"BF0F77E8",
    x"BF0F72B4",
    x"BF0F6D80",
    x"BF0F684B",
    x"BF0F6317",
    x"BF0F5DE2",
    x"BF0F58AE",
    x"BF0F5379",
    x"BF0F4E44",
    x"BF0F490F",
    x"BF0F43DA",
    x"BF0F3EA5",
    x"BF0F3970",
    x"BF0F343B",
    x"BF0F2F05",
    x"BF0F29D0",
    x"BF0F249B",
    x"BF0F1F65",
    x"BF0F1A2F",
    x"BF0F14FA",
    x"BF0F0FC4",
    x"BF0F0A8E",
    x"BF0F0558",
    x"BF0F0022",
    x"BF0EFAEB",
    x"BF0EF5B5",
    x"BF0EF07F",
    x"BF0EEB48",
    x"BF0EE612",
    x"BF0EE0DB",
    x"BF0EDBA4",
    x"BF0ED66E",
    x"BF0ED137",
    x"BF0ECC00",
    x"BF0EC6C9",
    x"BF0EC192",
    x"BF0EBC5A",
    x"BF0EB723",
    x"BF0EB1EC",
    x"BF0EACB4",
    x"BF0EA77D",
    x"BF0EA245",
    x"BF0E9D0D",
    x"BF0E97D5",
    x"BF0E929D",
    x"BF0E8D65",
    x"BF0E882D",
    x"BF0E82F5",
    x"BF0E7DBD",
    x"BF0E7885",
    x"BF0E734C",
    x"BF0E6E14",
    x"BF0E68DB",
    x"BF0E63A2",
    x"BF0E5E6A",
    x"BF0E5931",
    x"BF0E53F8",
    x"BF0E4EBF",
    x"BF0E4986",
    x"BF0E444C",
    x"BF0E3F13",
    x"BF0E39DA",
    x"BF0E34A0",
    x"BF0E2F67",
    x"BF0E2A2D",
    x"BF0E24F3",
    x"BF0E1FBA",
    x"BF0E1A80",
    x"BF0E1546",
    x"BF0E100C",
    x"BF0E0AD2",
    x"BF0E0597",
    x"BF0E005D",
    x"BF0DFB23",
    x"BF0DF5E8",
    x"BF0DF0AE",
    x"BF0DEB73",
    x"BF0DE638",
    x"BF0DE0FD",
    x"BF0DDBC2",
    x"BF0DD687",
    x"BF0DD14C",
    x"BF0DCC11",
    x"BF0DC6D6",
    x"BF0DC19B",
    x"BF0DBC5F",
    x"BF0DB724",
    x"BF0DB1E8",
    x"BF0DACAC",
    x"BF0DA771",
    x"BF0DA235",
    x"BF0D9CF9",
    x"BF0D97BD",
    x"BF0D9281",
    x"BF0D8D45",
    x"BF0D8808",
    x"BF0D82CC",
    x"BF0D7D8F",
    x"BF0D7853",
    x"BF0D7316",
    x"BF0D6DDA",
    x"BF0D689D",
    x"BF0D6360",
    x"BF0D5E23",
    x"BF0D58E6",
    x"BF0D53A9",
    x"BF0D4E6C",
    x"BF0D492E",
    x"BF0D43F1",
    x"BF0D3EB3",
    x"BF0D3976",
    x"BF0D3438",
    x"BF0D2EFA",
    x"BF0D29BD",
    x"BF0D247F",
    x"BF0D1F41",
    x"BF0D1A03",
    x"BF0D14C5",
    x"BF0D0F86",
    x"BF0D0A48",
    x"BF0D050A",
    x"BF0CFFCB",
    x"BF0CFA8D",
    x"BF0CF54E",
    x"BF0CF00F",
    x"BF0CEAD0",
    x"BF0CE591",
    x"BF0CE052",
    x"BF0CDB13",
    x"BF0CD5D4",
    x"BF0CD095",
    x"BF0CCB56",
    x"BF0CC616",
    x"BF0CC0D7",
    x"BF0CBB97",
    x"BF0CB657",
    x"BF0CB118",
    x"BF0CABD8",
    x"BF0CA698",
    x"BF0CA158",
    x"BF0C9C18",
    x"BF0C96D7",
    x"BF0C9197",
    x"BF0C8C57",
    x"BF0C8716",
    x"BF0C81D6",
    x"BF0C7C95",
    x"BF0C7755",
    x"BF0C7214",
    x"BF0C6CD3",
    x"BF0C6792",
    x"BF0C6251",
    x"BF0C5D10",
    x"BF0C57CF",
    x"BF0C528D",
    x"BF0C4D4C",
    x"BF0C480B",
    x"BF0C42C9",
    x"BF0C3D87",
    x"BF0C3846",
    x"BF0C3304",
    x"BF0C2DC2",
    x"BF0C2880",
    x"BF0C233E",
    x"BF0C1DFC",
    x"BF0C18BA",
    x"BF0C1377",
    x"BF0C0E35",
    x"BF0C08F2",
    x"BF0C03B0",
    x"BF0BFE6D",
    x"BF0BF92B",
    x"BF0BF3E8",
    x"BF0BEEA5",
    x"BF0BE962",
    x"BF0BE41F",
    x"BF0BDEDC",
    x"BF0BD998",
    x"BF0BD455",
    x"BF0BCF12",
    x"BF0BC9CE",
    x"BF0BC48B",
    x"BF0BBF47",
    x"BF0BBA03",
    x"BF0BB4BF",
    x"BF0BAF7C",
    x"BF0BAA38",
    x"BF0BA4F4",
    x"BF0B9FAF",
    x"BF0B9A6B",
    x"BF0B9527",
    x"BF0B8FE2",
    x"BF0B8A9E",
    x"BF0B8559",
    x"BF0B8015",
    x"BF0B7AD0",
    x"BF0B758B",
    x"BF0B7046",
    x"BF0B6B01",
    x"BF0B65BC",
    x"BF0B6077",
    x"BF0B5B32",
    x"BF0B55EC",
    x"BF0B50A7",
    x"BF0B4B61",
    x"BF0B461C",
    x"BF0B40D6",
    x"BF0B3B90",
    x"BF0B364B",
    x"BF0B3105",
    x"BF0B2BBF",
    x"BF0B2679",
    x"BF0B2132",
    x"BF0B1BEC",
    x"BF0B16A6",
    x"BF0B115F",
    x"BF0B0C19",
    x"BF0B06D2",
    x"BF0B018C",
    x"BF0AFC45",
    x"BF0AF6FE",
    x"BF0AF1B7",
    x"BF0AEC70",
    x"BF0AE729",
    x"BF0AE1E2",
    x"BF0ADC9B",
    x"BF0AD753",
    x"BF0AD20C",
    x"BF0ACCC4",
    x"BF0AC77D",
    x"BF0AC235",
    x"BF0ABCED",
    x"BF0AB7A5",
    x"BF0AB25E",
    x"BF0AAD16",
    x"BF0AA7CD",
    x"BF0AA285",
    x"BF0A9D3D",
    x"BF0A97F5",
    x"BF0A92AC",
    x"BF0A8D64",
    x"BF0A881B",
    x"BF0A82D2",
    x"BF0A7D8A",
    x"BF0A7841",
    x"BF0A72F8",
    x"BF0A6DAF",
    x"BF0A6866",
    x"BF0A631D",
    x"BF0A5DD3",
    x"BF0A588A",
    x"BF0A5341",
    x"BF0A4DF7",
    x"BF0A48AD",
    x"BF0A4364",
    x"BF0A3E1A",
    x"BF0A38D0",
    x"BF0A3386",
    x"BF0A2E3C",
    x"BF0A28F2",
    x"BF0A23A8",
    x"BF0A1E5E",
    x"BF0A1913",
    x"BF0A13C9",
    x"BF0A0E7E",
    x"BF0A0934",
    x"BF0A03E9",
    x"BF09FE9E",
    x"BF09F954",
    x"BF09F409",
    x"BF09EEBE",
    x"BF09E973",
    x"BF09E427",
    x"BF09DEDC",
    x"BF09D991",
    x"BF09D445",
    x"BF09CEFA",
    x"BF09C9AE",
    x"BF09C463",
    x"BF09BF17",
    x"BF09B9CB",
    x"BF09B47F",
    x"BF09AF33",
    x"BF09A9E7",
    x"BF09A49B",
    x"BF099F4E",
    x"BF099A02",
    x"BF0994B6",
    x"BF098F69",
    x"BF098A1D",
    x"BF0984D0",
    x"BF097F83",
    x"BF097A36",
    x"BF0974E9",
    x"BF096F9C",
    x"BF096A4F",
    x"BF096502",
    x"BF095FB5",
    x"BF095A68",
    x"BF09551A",
    x"BF094FCD",
    x"BF094A7F",
    x"BF094531",
    x"BF093FE4",
    x"BF093A96",
    x"BF093548",
    x"BF092FFA",
    x"BF092AAC",
    x"BF09255E",
    x"BF092010",
    x"BF091AC1",
    x"BF091573",
    x"BF091024",
    x"BF090AD6",
    x"BF090587",
    x"BF090038",
    x"BF08FAEA",
    x"BF08F59B",
    x"BF08F04C",
    x"BF08EAFD",
    x"BF08E5AD",
    x"BF08E05E",
    x"BF08DB0F",
    x"BF08D5BF",
    x"BF08D070",
    x"BF08CB20",
    x"BF08C5D1",
    x"BF08C081",
    x"BF08BB31",
    x"BF08B5E1",
    x"BF08B091",
    x"BF08AB41",
    x"BF08A5F1",
    x"BF08A0A1",
    x"BF089B51",
    x"BF089600",
    x"BF0890B0",
    x"BF088B5F",
    x"BF08860F",
    x"BF0880BE",
    x"BF087B6D",
    x"BF08761C",
    x"BF0870CB",
    x"BF086B7A",
    x"BF086629",
    x"BF0860D8",
    x"BF085B87",
    x"BF085635",
    x"BF0850E4",
    x"BF084B92",
    x"BF084641",
    x"BF0840EF",
    x"BF083B9D",
    x"BF08364B",
    x"BF0830F9",
    x"BF082BA7",
    x"BF082655",
    x"BF082103",
    x"BF081BB1",
    x"BF08165E",
    x"BF08110C",
    x"BF080BB9",
    x"BF080667",
    x"BF080114",
    x"BF07FBC1",
    x"BF07F66F",
    x"BF07F11C",
    x"BF07EBC9",
    x"BF07E676",
    x"BF07E122",
    x"BF07DBCF",
    x"BF07D67C",
    x"BF07D128",
    x"BF07CBD5",
    x"BF07C681",
    x"BF07C12E",
    x"BF07BBDA",
    x"BF07B686",
    x"BF07B132",
    x"BF07ABDE",
    x"BF07A68A",
    x"BF07A136",
    x"BF079BE2",
    x"BF07968D",
    x"BF079139",
    x"BF078BE4",
    x"BF078690",
    x"BF07813B",
    x"BF077BE6",
    x"BF077692",
    x"BF07713D",
    x"BF076BE8",
    x"BF076693",
    x"BF07613E",
    x"BF075BE8",
    x"BF075693",
    x"BF07513E",
    x"BF074BE8",
    x"BF074693",
    x"BF07413D",
    x"BF073BE7",
    x"BF073692",
    x"BF07313C",
    x"BF072BE6",
    x"BF072690",
    x"BF07213A",
    x"BF071BE3",
    x"BF07168D",
    x"BF071137",
    x"BF070BE0",
    x"BF07068A",
    x"BF070133",
    x"BF06FBDD",
    x"BF06F686",
    x"BF06F12F",
    x"BF06EBD8",
    x"BF06E681",
    x"BF06E12A",
    x"BF06DBD3",
    x"BF06D67B",
    x"BF06D124",
    x"BF06CBCD",
    x"BF06C675",
    x"BF06C11E",
    x"BF06BBC6",
    x"BF06B66E",
    x"BF06B116",
    x"BF06ABBF",
    x"BF06A667",
    x"BF06A10E",
    x"BF069BB6",
    x"BF06965E",
    x"BF069106",
    x"BF068BAD",
    x"BF068655",
    x"BF0680FC",
    x"BF067BA4",
    x"BF06764B",
    x"BF0670F2",
    x"BF066B99",
    x"BF066640",
    x"BF0660E7",
    x"BF065B8E",
    x"BF065635",
    x"BF0650DC",
    x"BF064B82",
    x"BF064629",
    x"BF0640CF",
    x"BF063B76",
    x"BF06361C",
    x"BF0630C2",
    x"BF062B69",
    x"BF06260F",
    x"BF0620B5",
    x"BF061B5B",
    x"BF061600",
    x"BF0610A6",
    x"BF060B4C",
    x"BF0605F1",
    x"BF060097",
    x"BF05FB3C",
    x"BF05F5E2",
    x"BF05F087",
    x"BF05EB2C",
    x"BF05E5D1",
    x"BF05E076",
    x"BF05DB1B",
    x"BF05D5C0",
    x"BF05D065",
    x"BF05CB0A",
    x"BF05C5AE",
    x"BF05C053",
    x"BF05BAF7",
    x"BF05B59C",
    x"BF05B040",
    x"BF05AAE4",
    x"BF05A588",
    x"BF05A02C",
    x"BF059AD0",
    x"BF059574",
    x"BF059018",
    x"BF058ABC",
    x"BF05855F",
    x"BF058003",
    x"BF057AA6",
    x"BF05754A",
    x"BF056FED",
    x"BF056A90",
    x"BF056534",
    x"BF055FD7",
    x"BF055A7A",
    x"BF05551D",
    x"BF054FBF",
    x"BF054A62",
    x"BF054505",
    x"BF053FA8",
    x"BF053A4A",
    x"BF0534EC",
    x"BF052F8F",
    x"BF052A31",
    x"BF0524D3",
    x"BF051F75",
    x"BF051A18",
    x"BF0514BA",
    x"BF050F5B",
    x"BF0509FD",
    x"BF05049F",
    x"BF04FF41",
    x"BF04F9E2",
    x"BF04F484",
    x"BF04EF25",
    x"BF04E9C6",
    x"BF04E468",
    x"BF04DF09",
    x"BF04D9AA",
    x"BF04D44B",
    x"BF04CEEC",
    x"BF04C98D",
    x"BF04C42D",
    x"BF04BECE",
    x"BF04B96F",
    x"BF04B40F",
    x"BF04AEB0",
    x"BF04A950",
    x"BF04A3F0",
    x"BF049E91",
    x"BF049931",
    x"BF0493D1",
    x"BF048E71",
    x"BF048911",
    x"BF0483B0",
    x"BF047E50",
    x"BF0478F0",
    x"BF04738F",
    x"BF046E2F",
    x"BF0468CE",
    x"BF04636E",
    x"BF045E0D",
    x"BF0458AC",
    x"BF04534B",
    x"BF044DEA",
    x"BF044889",
    x"BF044328",
    x"BF043DC7",
    x"BF043865",
    x"BF043304",
    x"BF042DA2",
    x"BF042841",
    x"BF0422DF",
    x"BF041D7E",
    x"BF04181C",
    x"BF0412BA",
    x"BF040D58",
    x"BF0407F6",
    x"BF040294",
    x"BF03FD32",
    x"BF03F7CF",
    x"BF03F26D",
    x"BF03ED0B",
    x"BF03E7A8",
    x"BF03E246",
    x"BF03DCE3",
    x"BF03D780",
    x"BF03D21D",
    x"BF03CCBA",
    x"BF03C757",
    x"BF03C1F4",
    x"BF03BC91",
    x"BF03B72E",
    x"BF03B1CB",
    x"BF03AC67",
    x"BF03A704",
    x"BF03A1A0",
    x"BF039C3D",
    x"BF0396D9",
    x"BF039175",
    x"BF038C11",
    x"BF0386AE",
    x"BF03814A",
    x"BF037BE5",
    x"BF037681",
    x"BF03711D",
    x"BF036BB9",
    x"BF036654",
    x"BF0360F0",
    x"BF035B8B",
    x"BF035627",
    x"BF0350C2",
    x"BF034B5D",
    x"BF0345F8",
    x"BF034093",
    x"BF033B2E",
    x"BF0335C9",
    x"BF033064",
    x"BF032AFF",
    x"BF032599",
    x"BF032034",
    x"BF031ACE",
    x"BF031569",
    x"BF031003",
    x"BF030A9D",
    x"BF030537",
    x"BF02FFD2",
    x"BF02FA6C",
    x"BF02F506",
    x"BF02EF9F",
    x"BF02EA39",
    x"BF02E4D3",
    x"BF02DF6C",
    x"BF02DA06",
    x"BF02D49F",
    x"BF02CF39",
    x"BF02C9D2",
    x"BF02C46B",
    x"BF02BF05",
    x"BF02B99E",
    x"BF02B437",
    x"BF02AED0",
    x"BF02A968",
    x"BF02A401",
    x"BF029E9A",
    x"BF029932",
    x"BF0293CB",
    x"BF028E63",
    x"BF0288FC",
    x"BF028394",
    x"BF027E2C",
    x"BF0278C4",
    x"BF02735C",
    x"BF026DF4",
    x"BF02688C",
    x"BF026324",
    x"BF025DBC",
    x"BF025853",
    x"BF0252EB",
    x"BF024D82",
    x"BF02481A",
    x"BF0242B1",
    x"BF023D48",
    x"BF0237E0",
    x"BF023277",
    x"BF022D0E",
    x"BF0227A5",
    x"BF02223C",
    x"BF021CD2",
    x"BF021769",
    x"BF021200",
    x"BF020C96",
    x"BF02072D",
    x"BF0201C3",
    x"BF01FC59",
    x"BF01F6F0",
    x"BF01F186",
    x"BF01EC1C",
    x"BF01E6B2",
    x"BF01E148",
    x"BF01DBDE",
    x"BF01D674",
    x"BF01D109",
    x"BF01CB9F",
    x"BF01C634",
    x"BF01C0CA",
    x"BF01BB5F",
    x"BF01B5F5",
    x"BF01B08A",
    x"BF01AB1F",
    x"BF01A5B4",
    x"BF01A049",
    x"BF019ADE",
    x"BF019573",
    x"BF019007",
    x"BF018A9C",
    x"BF018531",
    x"BF017FC5",
    x"BF017A5A",
    x"BF0174EE",
    x"BF016F82",
    x"BF016A17",
    x"BF0164AB",
    x"BF015F3F",
    x"BF0159D3",
    x"BF015467",
    x"BF014EFA",
    x"BF01498E",
    x"BF014422",
    x"BF013EB5",
    x"BF013949",
    x"BF0133DC",
    x"BF012E70",
    x"BF012903",
    x"BF012396",
    x"BF011E29",
    x"BF0118BC",
    x"BF01134F",
    x"BF010DE2",
    x"BF010875",
    x"BF010308",
    x"BF00FD9A",
    x"BF00F82D",
    x"BF00F2BF",
    x"BF00ED52",
    x"BF00E7E4",
    x"BF00E276",
    x"BF00DD09",
    x"BF00D79B",
    x"BF00D22D",
    x"BF00CCBF",
    x"BF00C751",
    x"BF00C1E2",
    x"BF00BC74",
    x"BF00B706",
    x"BF00B197",
    x"BF00AC29",
    x"BF00A6BA",
    x"BF00A14C",
    x"BF009BDD",
    x"BF00966E",
    x"BF0090FF",
    x"BF008B90",
    x"BF008621",
    x"BF0080B2",
    x"BF007B43",
    x"BF0075D4",
    x"BF007064",
    x"BF006AF5",
    x"BF006585",
    x"BF006016",
    x"BF005AA6",
    x"BF005536",
    x"BF004FC6",
    x"BF004A56",
    x"BF0044E6",
    x"BF003F76",
    x"BF003A06",
    x"BF003496",
    x"BF002F26",
    x"BF0029B5",
    x"BF002445",
    x"BF001ED4",
    x"BF001964",
    x"BF0013F3",
    x"BF000E82",
    x"BF000912",
    x"BF0003A1",
    x"BEFFFC5F",
    x"BEFFF17D",
    x"BEFFE69B",
    x"BEFFDBB8",
    x"BEFFD0D6",
    x"BEFFC5F3",
    x"BEFFBB10",
    x"BEFFB02D",
    x"BEFFA54A",
    x"BEFF9A67",
    x"BEFF8F83",
    x"BEFF849F",
    x"BEFF79BC",
    x"BEFF6ED8",
    x"BEFF63F4",
    x"BEFF590F",
    x"BEFF4E2B",
    x"BEFF4346",
    x"BEFF3862",
    x"BEFF2D7D",
    x"BEFF2298",
    x"BEFF17B2",
    x"BEFF0CCD",
    x"BEFF01E8",
    x"BEFEF702",
    x"BEFEEC1C",
    x"BEFEE136",
    x"BEFED650",
    x"BEFECB6A",
    x"BEFEC083",
    x"BEFEB59D",
    x"BEFEAAB6",
    x"BEFE9FCF",
    x"BEFE94E8",
    x"BEFE8A01",
    x"BEFE7F19",
    x"BEFE7432",
    x"BEFE694A",
    x"BEFE5E62",
    x"BEFE537A",
    x"BEFE4892",
    x"BEFE3DAA",
    x"BEFE32C2",
    x"BEFE27D9",
    x"BEFE1CF0",
    x"BEFE1207",
    x"BEFE071E",
    x"BEFDFC35",
    x"BEFDF14C",
    x"BEFDE662",
    x"BEFDDB79",
    x"BEFDD08F",
    x"BEFDC5A5",
    x"BEFDBABB",
    x"BEFDAFD1",
    x"BEFDA4E6",
    x"BEFD99FC",
    x"BEFD8F11",
    x"BEFD8426",
    x"BEFD793B",
    x"BEFD6E50",
    x"BEFD6365",
    x"BEFD5879",
    x"BEFD4D8D",
    x"BEFD42A2",
    x"BEFD37B6",
    x"BEFD2CCA",
    x"BEFD21DD",
    x"BEFD16F1",
    x"BEFD0C04",
    x"BEFD0118",
    x"BEFCF62B",
    x"BEFCEB3E",
    x"BEFCE051",
    x"BEFCD563",
    x"BEFCCA76",
    x"BEFCBF88",
    x"BEFCB49B",
    x"BEFCA9AD",
    x"BEFC9EBF",
    x"BEFC93D0",
    x"BEFC88E2",
    x"BEFC7DF3",
    x"BEFC7305",
    x"BEFC6816",
    x"BEFC5D27",
    x"BEFC5238",
    x"BEFC4748",
    x"BEFC3C59",
    x"BEFC3169",
    x"BEFC267A",
    x"BEFC1B8A",
    x"BEFC109A",
    x"BEFC05AA",
    x"BEFBFAB9",
    x"BEFBEFC9",
    x"BEFBE4D8",
    x"BEFBD9E7",
    x"BEFBCEF6",
    x"BEFBC405",
    x"BEFBB914",
    x"BEFBAE22",
    x"BEFBA331",
    x"BEFB983F",
    x"BEFB8D4D",
    x"BEFB825B",
    x"BEFB7769",
    x"BEFB6C77",
    x"BEFB6184",
    x"BEFB5692",
    x"BEFB4B9F",
    x"BEFB40AC",
    x"BEFB35B9",
    x"BEFB2AC6",
    x"BEFB1FD2",
    x"BEFB14DF",
    x"BEFB09EB",
    x"BEFAFEF7",
    x"BEFAF403",
    x"BEFAE90F",
    x"BEFADE1B",
    x"BEFAD326",
    x"BEFAC832",
    x"BEFABD3D",
    x"BEFAB248",
    x"BEFAA753",
    x"BEFA9C5E",
    x"BEFA9169",
    x"BEFA8673",
    x"BEFA7B7D",
    x"BEFA7088",
    x"BEFA6592",
    x"BEFA5A9C",
    x"BEFA4FA5",
    x"BEFA44AF",
    x"BEFA39B8",
    x"BEFA2EC2",
    x"BEFA23CB",
    x"BEFA18D4",
    x"BEFA0DDD",
    x"BEFA02E5",
    x"BEF9F7EE",
    x"BEF9ECF6",
    x"BEF9E1FE",
    x"BEF9D707",
    x"BEF9CC0E",
    x"BEF9C116",
    x"BEF9B61E",
    x"BEF9AB25",
    x"BEF9A02D",
    x"BEF99534",
    x"BEF98A3B",
    x"BEF97F42",
    x"BEF97449",
    x"BEF9694F",
    x"BEF95E56",
    x"BEF9535C",
    x"BEF94862",
    x"BEF93D68",
    x"BEF9326E",
    x"BEF92773",
    x"BEF91C79",
    x"BEF9117E",
    x"BEF90684",
    x"BEF8FB89",
    x"BEF8F08E",
    x"BEF8E592",
    x"BEF8DA97",
    x"BEF8CF9C",
    x"BEF8C4A0",
    x"BEF8B9A4",
    x"BEF8AEA8",
    x"BEF8A3AC",
    x"BEF898B0",
    x"BEF88DB3",
    x"BEF882B7",
    x"BEF877BA",
    x"BEF86CBD",
    x"BEF861C0",
    x"BEF856C3",
    x"BEF84BC6",
    x"BEF840C8",
    x"BEF835CB",
    x"BEF82ACD",
    x"BEF81FCF",
    x"BEF814D1",
    x"BEF809D3",
    x"BEF7FED4",
    x"BEF7F3D6",
    x"BEF7E8D7",
    x"BEF7DDD8",
    x"BEF7D2D9",
    x"BEF7C7DA",
    x"BEF7BCDB",
    x"BEF7B1DC",
    x"BEF7A6DC",
    x"BEF79BDC",
    x"BEF790DC",
    x"BEF785DC",
    x"BEF77ADC",
    x"BEF76FDC",
    x"BEF764DC",
    x"BEF759DB",
    x"BEF74EDA",
    x"BEF743D9",
    x"BEF738D8",
    x"BEF72DD7",
    x"BEF722D6",
    x"BEF717D4",
    x"BEF70CD3",
    x"BEF701D1",
    x"BEF6F6CF",
    x"BEF6EBCD",
    x"BEF6E0CB",
    x"BEF6D5C8",
    x"BEF6CAC6",
    x"BEF6BFC3",
    x"BEF6B4C0",
    x"BEF6A9BD",
    x"BEF69EBA",
    x"BEF693B7",
    x"BEF688B3",
    x"BEF67DB0",
    x"BEF672AC",
    x"BEF667A8",
    x"BEF65CA4",
    x"BEF651A0",
    x"BEF6469C",
    x"BEF63B97",
    x"BEF63093",
    x"BEF6258E",
    x"BEF61A89",
    x"BEF60F84",
    x"BEF6047F",
    x"BEF5F979",
    x"BEF5EE74",
    x"BEF5E36E",
    x"BEF5D868",
    x"BEF5CD62",
    x"BEF5C25C",
    x"BEF5B756",
    x"BEF5AC50",
    x"BEF5A149",
    x"BEF59643",
    x"BEF58B3C",
    x"BEF58035",
    x"BEF5752E",
    x"BEF56A26",
    x"BEF55F1F",
    x"BEF55417",
    x"BEF54910",
    x"BEF53E08",
    x"BEF53300",
    x"BEF527F8",
    x"BEF51CEF",
    x"BEF511E7",
    x"BEF506DE",
    x"BEF4FBD5",
    x"BEF4F0CC",
    x"BEF4E5C3",
    x"BEF4DABA",
    x"BEF4CFB1",
    x"BEF4C4A7",
    x"BEF4B99E",
    x"BEF4AE94",
    x"BEF4A38A",
    x"BEF49880",
    x"BEF48D76",
    x"BEF4826B",
    x"BEF47761",
    x"BEF46C56",
    x"BEF4614B",
    x"BEF45640",
    x"BEF44B35",
    x"BEF4402A",
    x"BEF4351F",
    x"BEF42A13",
    x"BEF41F07",
    x"BEF413FB",
    x"BEF408F0",
    x"BEF3FDE3",
    x"BEF3F2D7",
    x"BEF3E7CB",
    x"BEF3DCBE",
    x"BEF3D1B1",
    x"BEF3C6A4",
    x"BEF3BB97",
    x"BEF3B08A",
    x"BEF3A57D",
    x"BEF39A6F",
    x"BEF38F62",
    x"BEF38454",
    x"BEF37946",
    x"BEF36E38",
    x"BEF3632A",
    x"BEF3581C",
    x"BEF34D0D",
    x"BEF341FE",
    x"BEF336F0",
    x"BEF32BE1",
    x"BEF320D2",
    x"BEF315C2",
    x"BEF30AB3",
    x"BEF2FFA4",
    x"BEF2F494",
    x"BEF2E984",
    x"BEF2DE74",
    x"BEF2D364",
    x"BEF2C854",
    x"BEF2BD43",
    x"BEF2B233",
    x"BEF2A722",
    x"BEF29C11",
    x"BEF29100",
    x"BEF285EF",
    x"BEF27ADE",
    x"BEF26FCD",
    x"BEF264BB",
    x"BEF259A9",
    x"BEF24E97",
    x"BEF24385",
    x"BEF23873",
    x"BEF22D61",
    x"BEF2224F",
    x"BEF2173C",
    x"BEF20C29",
    x"BEF20116",
    x"BEF1F603",
    x"BEF1EAF0",
    x"BEF1DFDD",
    x"BEF1D4C9",
    x"BEF1C9B6",
    x"BEF1BEA2",
    x"BEF1B38E",
    x"BEF1A87A",
    x"BEF19D66",
    x"BEF19252",
    x"BEF1873D",
    x"BEF17C28",
    x"BEF17114",
    x"BEF165FF",
    x"BEF15AEA",
    x"BEF14FD5",
    x"BEF144BF",
    x"BEF139AA",
    x"BEF12E94",
    x"BEF1237E",
    x"BEF11868",
    x"BEF10D52",
    x"BEF1023C",
    x"BEF0F726",
    x"BEF0EC0F",
    x"BEF0E0F9",
    x"BEF0D5E2",
    x"BEF0CACB",
    x"BEF0BFB4",
    x"BEF0B49C",
    x"BEF0A985",
    x"BEF09E6E",
    x"BEF09356",
    x"BEF0883E",
    x"BEF07D26",
    x"BEF0720E",
    x"BEF066F6",
    x"BEF05BDD",
    x"BEF050C5",
    x"BEF045AC",
    x"BEF03A93",
    x"BEF02F7A",
    x"BEF02461",
    x"BEF01948",
    x"BEF00E2E",
    x"BEF00315",
    x"BEEFF7FB",
    x"BEEFECE1",
    x"BEEFE1C7",
    x"BEEFD6AD",
    x"BEEFCB93",
    x"BEEFC079",
    x"BEEFB55E",
    x"BEEFAA43",
    x"BEEF9F28",
    x"BEEF940D",
    x"BEEF88F2",
    x"BEEF7DD7",
    x"BEEF72BC",
    x"BEEF67A0",
    x"BEEF5C84",
    x"BEEF5168",
    x"BEEF464C",
    x"BEEF3B30",
    x"BEEF3014",
    x"BEEF24F7",
    x"BEEF19DB",
    x"BEEF0EBE",
    x"BEEF03A1",
    x"BEEEF884",
    x"BEEEED67",
    x"BEEEE24A",
    x"BEEED72C",
    x"BEEECC0F",
    x"BEEEC0F1",
    x"BEEEB5D3",
    x"BEEEAAB5",
    x"BEEE9F97",
    x"BEEE9479",
    x"BEEE895A",
    x"BEEE7E3C",
    x"BEEE731D",
    x"BEEE67FE",
    x"BEEE5CDF",
    x"BEEE51C0",
    x"BEEE46A0",
    x"BEEE3B81",
    x"BEEE3061",
    x"BEEE2542",
    x"BEEE1A22",
    x"BEEE0F02",
    x"BEEE03E2",
    x"BEEDF8C1",
    x"BEEDEDA1",
    x"BEEDE280",
    x"BEEDD75F",
    x"BEEDCC3E",
    x"BEEDC11D",
    x"BEEDB5FC",
    x"BEEDAADB",
    x"BEED9FB9",
    x"BEED9498",
    x"BEED8976",
    x"BEED7E54",
    x"BEED7332",
    x"BEED6810",
    x"BEED5CEE",
    x"BEED51CB",
    x"BEED46A9",
    x"BEED3B86",
    x"BEED3063",
    x"BEED2540",
    x"BEED1A1D",
    x"BEED0EF9",
    x"BEED03D6",
    x"BEECF8B2",
    x"BEECED8F",
    x"BEECE26B",
    x"BEECD747",
    x"BEECCC22",
    x"BEECC0FE",
    x"BEECB5DA",
    x"BEECAAB5",
    x"BEEC9F90",
    x"BEEC946B",
    x"BEEC8946",
    x"BEEC7E21",
    x"BEEC72FC",
    x"BEEC67D6",
    x"BEEC5CB1",
    x"BEEC518B",
    x"BEEC4665",
    x"BEEC3B3F",
    x"BEEC3019",
    x"BEEC24F3",
    x"BEEC19CC",
    x"BEEC0EA5",
    x"BEEC037F",
    x"BEEBF858",
    x"BEEBED31",
    x"BEEBE20A",
    x"BEEBD6E2",
    x"BEEBCBBB",
    x"BEEBC093",
    x"BEEBB56C",
    x"BEEBAA44",
    x"BEEB9F1C",
    x"BEEB93F3",
    x"BEEB88CB",
    x"BEEB7DA3",
    x"BEEB727A",
    x"BEEB6751",
    x"BEEB5C28",
    x"BEEB50FF",
    x"BEEB45D6",
    x"BEEB3AAD",
    x"BEEB2F84",
    x"BEEB245A",
    x"BEEB1930",
    x"BEEB0E06",
    x"BEEB02DC",
    x"BEEAF7B2",
    x"BEEAEC88",
    x"BEEAE15D",
    x"BEEAD633",
    x"BEEACB08",
    x"BEEABFDD",
    x"BEEAB4B2",
    x"BEEAA987",
    x"BEEA9E5C",
    x"BEEA9330",
    x"BEEA8805",
    x"BEEA7CD9",
    x"BEEA71AD",
    x"BEEA6681",
    x"BEEA5B55",
    x"BEEA5029",
    x"BEEA44FD",
    x"BEEA39D0",
    x"BEEA2EA3",
    x"BEEA2376",
    x"BEEA1849",
    x"BEEA0D1C",
    x"BEEA01EF",
    x"BEE9F6C2",
    x"BEE9EB94",
    x"BEE9E066",
    x"BEE9D539",
    x"BEE9CA0B",
    x"BEE9BEDD",
    x"BEE9B3AE",
    x"BEE9A880",
    x"BEE99D51",
    x"BEE99223",
    x"BEE986F4",
    x"BEE97BC5",
    x"BEE97096",
    x"BEE96567",
    x"BEE95A37",
    x"BEE94F08",
    x"BEE943D8",
    x"BEE938A8",
    x"BEE92D78",
    x"BEE92248",
    x"BEE91718",
    x"BEE90BE8",
    x"BEE900B7",
    x"BEE8F587",
    x"BEE8EA56",
    x"BEE8DF25",
    x"BEE8D3F4",
    x"BEE8C8C3",
    x"BEE8BD91",
    x"BEE8B260",
    x"BEE8A72E",
    x"BEE89BFD",
    x"BEE890CB",
    x"BEE88599",
    x"BEE87A66",
    x"BEE86F34",
    x"BEE86402",
    x"BEE858CF",
    x"BEE84D9C",
    x"BEE84269",
    x"BEE83736",
    x"BEE82C03",
    x"BEE820D0",
    x"BEE8159C",
    x"BEE80A69",
    x"BEE7FF35",
    x"BEE7F401",
    x"BEE7E8CD",
    x"BEE7DD99",
    x"BEE7D265",
    x"BEE7C731",
    x"BEE7BBFC",
    x"BEE7B0C7",
    x"BEE7A592",
    x"BEE79A5D",
    x"BEE78F28",
    x"BEE783F3",
    x"BEE778BE",
    x"BEE76D88",
    x"BEE76253",
    x"BEE7571D",
    x"BEE74BE7",
    x"BEE740B1",
    x"BEE7357A",
    x"BEE72A44",
    x"BEE71F0E",
    x"BEE713D7",
    x"BEE708A0",
    x"BEE6FD69",
    x"BEE6F232",
    x"BEE6E6FB",
    x"BEE6DBC4",
    x"BEE6D08C",
    x"BEE6C554",
    x"BEE6BA1D",
    x"BEE6AEE5",
    x"BEE6A3AD",
    x"BEE69875",
    x"BEE68D3C",
    x"BEE68204",
    x"BEE676CB",
    x"BEE66B93",
    x"BEE6605A",
    x"BEE65521",
    x"BEE649E7",
    x"BEE63EAE",
    x"BEE63375",
    x"BEE6283B",
    x"BEE61D02",
    x"BEE611C8",
    x"BEE6068E",
    x"BEE5FB54",
    x"BEE5F019",
    x"BEE5E4DF",
    x"BEE5D9A4",
    x"BEE5CE6A",
    x"BEE5C32F",
    x"BEE5B7F4",
    x"BEE5ACB9",
    x"BEE5A17E",
    x"BEE59642",
    x"BEE58B07",
    x"BEE57FCB",
    x"BEE5748F",
    x"BEE56953",
    x"BEE55E17",
    x"BEE552DB",
    x"BEE5479F",
    x"BEE53C62",
    x"BEE53126",
    x"BEE525E9",
    x"BEE51AAC",
    x"BEE50F6F",
    x"BEE50432",
    x"BEE4F8F5",
    x"BEE4EDB7",
    x"BEE4E27A",
    x"BEE4D73C",
    x"BEE4CBFE",
    x"BEE4C0C0",
    x"BEE4B582",
    x"BEE4AA44",
    x"BEE49F05",
    x"BEE493C7",
    x"BEE48888",
    x"BEE47D49",
    x"BEE4720A",
    x"BEE466CB",
    x"BEE45B8C",
    x"BEE4504D",
    x"BEE4450D",
    x"BEE439CE",
    x"BEE42E8E",
    x"BEE4234E",
    x"BEE4180E",
    x"BEE40CCE",
    x"BEE4018D",
    x"BEE3F64D",
    x"BEE3EB0C",
    x"BEE3DFCB",
    x"BEE3D48B",
    x"BEE3C94A",
    x"BEE3BE08",
    x"BEE3B2C7",
    x"BEE3A786",
    x"BEE39C44",
    x"BEE39102",
    x"BEE385C1",
    x"BEE37A7F",
    x"BEE36F3D",
    x"BEE363FA",
    x"BEE358B8",
    x"BEE34D75",
    x"BEE34233",
    x"BEE336F0",
    x"BEE32BAD",
    x"BEE3206A",
    x"BEE31527",
    x"BEE309E3",
    x"BEE2FEA0",
    x"BEE2F35C",
    x"BEE2E819",
    x"BEE2DCD5",
    x"BEE2D191",
    x"BEE2C64C",
    x"BEE2BB08",
    x"BEE2AFC4",
    x"BEE2A47F",
    x"BEE2993A",
    x"BEE28DF6",
    x"BEE282B1",
    x"BEE2776C",
    x"BEE26C26",
    x"BEE260E1",
    x"BEE2559B",
    x"BEE24A56",
    x"BEE23F10",
    x"BEE233CA",
    x"BEE22884",
    x"BEE21D3E",
    x"BEE211F7",
    x"BEE206B1",
    x"BEE1FB6A",
    x"BEE1F023",
    x"BEE1E4DD",
    x"BEE1D996",
    x"BEE1CE4E",
    x"BEE1C307",
    x"BEE1B7C0",
    x"BEE1AC78",
    x"BEE1A130",
    x"BEE195E9",
    x"BEE18AA1",
    x"BEE17F58",
    x"BEE17410",
    x"BEE168C8",
    x"BEE15D7F",
    x"BEE15237",
    x"BEE146EE",
    x"BEE13BA5",
    x"BEE1305C",
    x"BEE12513",
    x"BEE119C9",
    x"BEE10E80",
    x"BEE10336",
    x"BEE0F7ED",
    x"BEE0ECA3",
    x"BEE0E159",
    x"BEE0D60E",
    x"BEE0CAC4",
    x"BEE0BF7A",
    x"BEE0B42F",
    x"BEE0A8E5",
    x"BEE09D9A",
    x"BEE0924F",
    x"BEE08704",
    x"BEE07BB8",
    x"BEE0706D",
    x"BEE06522",
    x"BEE059D6",
    x"BEE04E8A",
    x"BEE0433E",
    x"BEE037F2",
    x"BEE02CA6",
    x"BEE0215A",
    x"BEE0160D",
    x"BEE00AC1",
    x"BEDFFF74",
    x"BEDFF427",
    x"BEDFE8DA",
    x"BEDFDD8D",
    x"BEDFD240",
    x"BEDFC6F2",
    x"BEDFBBA5",
    x"BEDFB057",
    x"BEDFA509",
    x"BEDF99BB",
    x"BEDF8E6D",
    x"BEDF831F",
    x"BEDF77D1",
    x"BEDF6C82",
    x"BEDF6134",
    x"BEDF55E5",
    x"BEDF4A96",
    x"BEDF3F47",
    x"BEDF33F8",
    x"BEDF28A9",
    x"BEDF1D59",
    x"BEDF120A",
    x"BEDF06BA",
    x"BEDEFB6A",
    x"BEDEF01A",
    x"BEDEE4CA",
    x"BEDED97A",
    x"BEDECE2A",
    x"BEDEC2D9",
    x"BEDEB789",
    x"BEDEAC38",
    x"BEDEA0E7",
    x"BEDE9596",
    x"BEDE8A45",
    x"BEDE7EF3",
    x"BEDE73A2",
    x"BEDE6851",
    x"BEDE5CFF",
    x"BEDE51AD",
    x"BEDE465B",
    x"BEDE3B09",
    x"BEDE2FB7",
    x"BEDE2464",
    x"BEDE1912",
    x"BEDE0DBF",
    x"BEDE026C",
    x"BEDDF71A",
    x"BEDDEBC7",
    x"BEDDE073",
    x"BEDDD520",
    x"BEDDC9CD",
    x"BEDDBE79",
    x"BEDDB325",
    x"BEDDA7D2",
    x"BEDD9C7E",
    x"BEDD912A",
    x"BEDD85D5",
    x"BEDD7A81",
    x"BEDD6F2C",
    x"BEDD63D8",
    x"BEDD5883",
    x"BEDD4D2E",
    x"BEDD41D9",
    x"BEDD3684",
    x"BEDD2B2F",
    x"BEDD1FD9",
    x"BEDD1484",
    x"BEDD092E",
    x"BEDCFDD8",
    x"BEDCF282",
    x"BEDCE72C",
    x"BEDCDBD6",
    x"BEDCD07F",
    x"BEDCC529",
    x"BEDCB9D2",
    x"BEDCAE7C",
    x"BEDCA325",
    x"BEDC97CE",
    x"BEDC8C76",
    x"BEDC811F",
    x"BEDC75C8",
    x"BEDC6A70",
    x"BEDC5F18",
    x"BEDC53C1",
    x"BEDC4869",
    x"BEDC3D11",
    x"BEDC31B8",
    x"BEDC2660",
    x"BEDC1B08",
    x"BEDC0FAF",
    x"BEDC0456",
    x"BEDBF8FD",
    x"BEDBEDA4",
    x"BEDBE24B",
    x"BEDBD6F2",
    x"BEDBCB98",
    x"BEDBC03F",
    x"BEDBB4E5",
    x"BEDBA98B",
    x"BEDB9E31",
    x"BEDB92D7",
    x"BEDB877D",
    x"BEDB7C23",
    x"BEDB70C8",
    x"BEDB656E",
    x"BEDB5A13",
    x"BEDB4EB8",
    x"BEDB435D",
    x"BEDB3802",
    x"BEDB2CA7",
    x"BEDB214B",
    x"BEDB15F0",
    x"BEDB0A94",
    x"BEDAFF38",
    x"BEDAF3DC",
    x"BEDAE880",
    x"BEDADD24",
    x"BEDAD1C8",
    x"BEDAC66B",
    x"BEDABB0F",
    x"BEDAAFB2",
    x"BEDAA455",
    x"BEDA98F8",
    x"BEDA8D9B",
    x"BEDA823E",
    x"BEDA76E0",
    x"BEDA6B83",
    x"BEDA6025",
    x"BEDA54C8",
    x"BEDA496A",
    x"BEDA3E0C",
    x"BEDA32AD",
    x"BEDA274F",
    x"BEDA1BF1",
    x"BEDA1092",
    x"BEDA0533",
    x"BED9F9D5",
    x"BED9EE76",
    x"BED9E317",
    x"BED9D7B7",
    x"BED9CC58",
    x"BED9C0F9",
    x"BED9B599",
    x"BED9AA39",
    x"BED99ED9",
    x"BED99379",
    x"BED98819",
    x"BED97CB9",
    x"BED97159",
    x"BED965F8",
    x"BED95A97",
    x"BED94F37",
    x"BED943D6",
    x"BED93875",
    x"BED92D13",
    x"BED921B2",
    x"BED91651",
    x"BED90AEF",
    x"BED8FF8D",
    x"BED8F42C",
    x"BED8E8CA",
    x"BED8DD67",
    x"BED8D205",
    x"BED8C6A3",
    x"BED8BB40",
    x"BED8AFDE",
    x"BED8A47B",
    x"BED89918",
    x"BED88DB5",
    x"BED88252",
    x"BED876EF",
    x"BED86B8B",
    x"BED86028",
    x"BED854C4",
    x"BED84960",
    x"BED83DFC",
    x"BED83298",
    x"BED82734",
    x"BED81BD0",
    x"BED8106B",
    x"BED80507",
    x"BED7F9A2",
    x"BED7EE3D",
    x"BED7E2D8",
    x"BED7D773",
    x"BED7CC0E",
    x"BED7C0A9",
    x"BED7B543",
    x"BED7A9DE",
    x"BED79E78",
    x"BED79312",
    x"BED787AC",
    x"BED77C46",
    x"BED770E0",
    x"BED76579",
    x"BED75A13",
    x"BED74EAC",
    x"BED74345",
    x"BED737DE",
    x"BED72C77",
    x"BED72110",
    x"BED715A9",
    x"BED70A41",
    x"BED6FEDA",
    x"BED6F372",
    x"BED6E80A",
    x"BED6DCA2",
    x"BED6D13A",
    x"BED6C5D2",
    x"BED6BA6A",
    x"BED6AF01",
    x"BED6A399",
    x"BED69830",
    x"BED68CC7",
    x"BED6815E",
    x"BED675F5",
    x"BED66A8C",
    x"BED65F22",
    x"BED653B9",
    x"BED6484F",
    x"BED63CE5",
    x"BED6317B",
    x"BED62611",
    x"BED61AA7",
    x"BED60F3D",
    x"BED603D3",
    x"BED5F868",
    x"BED5ECFD",
    x"BED5E193",
    x"BED5D628",
    x"BED5CABD",
    x"BED5BF52",
    x"BED5B3E6",
    x"BED5A87B",
    x"BED59D0F",
    x"BED591A4",
    x"BED58638",
    x"BED57ACC",
    x"BED56F60",
    x"BED563F3",
    x"BED55887",
    x"BED54D1B",
    x"BED541AE",
    x"BED53641",
    x"BED52AD5",
    x"BED51F68",
    x"BED513FA",
    x"BED5088D",
    x"BED4FD20",
    x"BED4F1B2",
    x"BED4E645",
    x"BED4DAD7",
    x"BED4CF69",
    x"BED4C3FB",
    x"BED4B88D",
    x"BED4AD1F",
    x"BED4A1B0",
    x"BED49642",
    x"BED48AD3",
    x"BED47F64",
    x"BED473F5",
    x"BED46886",
    x"BED45D17",
    x"BED451A8",
    x"BED44639",
    x"BED43AC9",
    x"BED42F59",
    x"BED423EA",
    x"BED4187A",
    x"BED40D0A",
    x"BED40199",
    x"BED3F629",
    x"BED3EAB9",
    x"BED3DF48",
    x"BED3D3D7",
    x"BED3C867",
    x"BED3BCF6",
    x"BED3B185",
    x"BED3A613",
    x"BED39AA2",
    x"BED38F31",
    x"BED383BF",
    x"BED3784D",
    x"BED36CDB",
    x"BED3616A",
    x"BED355F7",
    x"BED34A85",
    x"BED33F13",
    x"BED333A0",
    x"BED3282E",
    x"BED31CBB",
    x"BED31148",
    x"BED305D5",
    x"BED2FA62",
    x"BED2EEEF",
    x"BED2E37C",
    x"BED2D808",
    x"BED2CC94",
    x"BED2C121",
    x"BED2B5AD",
    x"BED2AA39",
    x"BED29EC5",
    x"BED29350",
    x"BED287DC",
    x"BED27C68",
    x"BED270F3",
    x"BED2657E",
    x"BED25A09",
    x"BED24E94",
    x"BED2431F",
    x"BED237AA",
    x"BED22C34",
    x"BED220BF",
    x"BED21549",
    x"BED209D3",
    x"BED1FE5E",
    x"BED1F2E8",
    x"BED1E771",
    x"BED1DBFB",
    x"BED1D085",
    x"BED1C50E",
    x"BED1B998",
    x"BED1AE21",
    x"BED1A2AA",
    x"BED19733",
    x"BED18BBC",
    x"BED18044",
    x"BED174CD",
    x"BED16955",
    x"BED15DDE",
    x"BED15266",
    x"BED146EE",
    x"BED13B76",
    x"BED12FFE",
    x"BED12485",
    x"BED1190D",
    x"BED10D95",
    x"BED1021C",
    x"BED0F6A3",
    x"BED0EB2A",
    x"BED0DFB1",
    x"BED0D438",
    x"BED0C8BF",
    x"BED0BD45",
    x"BED0B1CC",
    x"BED0A652",
    x"BED09AD8",
    x"BED08F5E",
    x"BED083E4",
    x"BED0786A",
    x"BED06CF0",
    x"BED06175",
    x"BED055FB",
    x"BED04A80",
    x"BED03F05",
    x"BED0338A",
    x"BED0280F",
    x"BED01C94",
    x"BED01119",
    x"BED0059D",
    x"BECFFA22",
    x"BECFEEA6",
    x"BECFE32A",
    x"BECFD7AE",
    x"BECFCC32",
    x"BECFC0B6",
    x"BECFB53A",
    x"BECFA9BD",
    x"BECF9E41",
    x"BECF92C4",
    x"BECF8747",
    x"BECF7BCA",
    x"BECF704D",
    x"BECF64D0",
    x"BECF5953",
    x"BECF4DD5",
    x"BECF4258",
    x"BECF36DA",
    x"BECF2B5C",
    x"BECF1FDE",
    x"BECF1460",
    x"BECF08E2",
    x"BECEFD64",
    x"BECEF1E5",
    x"BECEE667",
    x"BECEDAE8",
    x"BECECF69",
    x"BECEC3EA",
    x"BECEB86B",
    x"BECEACEC",
    x"BECEA16D",
    x"BECE95ED",
    x"BECE8A6E",
    x"BECE7EEE",
    x"BECE736E",
    x"BECE67EE",
    x"BECE5C6E",
    x"BECE50EE",
    x"BECE456E",
    x"BECE39ED",
    x"BECE2E6D",
    x"BECE22EC",
    x"BECE176B",
    x"BECE0BEA",
    x"BECE0069",
    x"BECDF4E8",
    x"BECDE967",
    x"BECDDDE5",
    x"BECDD264",
    x"BECDC6E2",
    x"BECDBB60",
    x"BECDAFDE",
    x"BECDA45C",
    x"BECD98DA",
    x"BECD8D58",
    x"BECD81D5",
    x"BECD7653",
    x"BECD6AD0",
    x"BECD5F4D",
    x"BECD53CA",
    x"BECD4847",
    x"BECD3CC4",
    x"BECD3141",
    x"BECD25BE",
    x"BECD1A3A",
    x"BECD0EB6",
    x"BECD0333",
    x"BECCF7AF",
    x"BECCEC2B",
    x"BECCE0A7",
    x"BECCD522",
    x"BECCC99E",
    x"BECCBE19",
    x"BECCB295",
    x"BECCA710",
    x"BECC9B8B",
    x"BECC9006",
    x"BECC8481",
    x"BECC78FC",
    x"BECC6D76",
    x"BECC61F1",
    x"BECC566B",
    x"BECC4AE5",
    x"BECC3F60",
    x"BECC33DA",
    x"BECC2853",
    x"BECC1CCD",
    x"BECC1147",
    x"BECC05C0",
    x"BECBFA3A",
    x"BECBEEB3",
    x"BECBE32C",
    x"BECBD7A5",
    x"BECBCC1E",
    x"BECBC097",
    x"BECBB50F",
    x"BECBA988",
    x"BECB9E00",
    x"BECB9279",
    x"BECB86F1",
    x"BECB7B69",
    x"BECB6FE1",
    x"BECB6459",
    x"BECB58D0",
    x"BECB4D48",
    x"BECB41BF",
    x"BECB3637",
    x"BECB2AAE",
    x"BECB1F25",
    x"BECB139C",
    x"BECB0813",
    x"BECAFC89",
    x"BECAF100",
    x"BECAE576",
    x"BECAD9ED",
    x"BECACE63",
    x"BECAC2D9",
    x"BECAB74F",
    x"BECAABC5",
    x"BECAA03A",
    x"BECA94B0",
    x"BECA8925",
    x"BECA7D9B",
    x"BECA7210",
    x"BECA6685",
    x"BECA5AFA",
    x"BECA4F6F",
    x"BECA43E4",
    x"BECA3858",
    x"BECA2CCD",
    x"BECA2141",
    x"BECA15B5",
    x"BECA0A2A",
    x"BEC9FE9E",
    x"BEC9F312",
    x"BEC9E785",
    x"BEC9DBF9",
    x"BEC9D06C",
    x"BEC9C4E0",
    x"BEC9B953",
    x"BEC9ADC6",
    x"BEC9A239",
    x"BEC996AC",
    x"BEC98B1F",
    x"BEC97F92",
    x"BEC97404",
    x"BEC96877",
    x"BEC95CE9",
    x"BEC9515B",
    x"BEC945CD",
    x"BEC93A3F",
    x"BEC92EB1",
    x"BEC92323",
    x"BEC91794",
    x"BEC90C06",
    x"BEC90077",
    x"BEC8F4E8",
    x"BEC8E959",
    x"BEC8DDCA",
    x"BEC8D23B",
    x"BEC8C6AC",
    x"BEC8BB1D",
    x"BEC8AF8D",
    x"BEC8A3FD",
    x"BEC8986E",
    x"BEC88CDE",
    x"BEC8814E",
    x"BEC875BE",
    x"BEC86A2D",
    x"BEC85E9D",
    x"BEC8530D",
    x"BEC8477C",
    x"BEC83BEB",
    x"BEC8305B",
    x"BEC824CA",
    x"BEC81938",
    x"BEC80DA7",
    x"BEC80216",
    x"BEC7F685",
    x"BEC7EAF3",
    x"BEC7DF61",
    x"BEC7D3CF",
    x"BEC7C83E",
    x"BEC7BCAC",
    x"BEC7B119",
    x"BEC7A587",
    x"BEC799F5",
    x"BEC78E62",
    x"BEC782D0",
    x"BEC7773D",
    x"BEC76BAA",
    x"BEC76017",
    x"BEC75484",
    x"BEC748F0",
    x"BEC73D5D",
    x"BEC731CA",
    x"BEC72636",
    x"BEC71AA2",
    x"BEC70F0E",
    x"BEC7037B",
    x"BEC6F7E6",
    x"BEC6EC52",
    x"BEC6E0BE",
    x"BEC6D529",
    x"BEC6C995",
    x"BEC6BE00",
    x"BEC6B26B",
    x"BEC6A6D6",
    x"BEC69B41",
    x"BEC68FAC",
    x"BEC68417",
    x"BEC67882",
    x"BEC66CEC",
    x"BEC66156",
    x"BEC655C1",
    x"BEC64A2B",
    x"BEC63E95",
    x"BEC632FF",
    x"BEC62768",
    x"BEC61BD2",
    x"BEC6103C",
    x"BEC604A5",
    x"BEC5F90E",
    x"BEC5ED77",
    x"BEC5E1E1",
    x"BEC5D649",
    x"BEC5CAB2",
    x"BEC5BF1B",
    x"BEC5B384",
    x"BEC5A7EC",
    x"BEC59C54",
    x"BEC590BD",
    x"BEC58525",
    x"BEC5798D",
    x"BEC56DF4",
    x"BEC5625C",
    x"BEC556C4",
    x"BEC54B2B",
    x"BEC53F93",
    x"BEC533FA",
    x"BEC52861",
    x"BEC51CC8",
    x"BEC5112F",
    x"BEC50596",
    x"BEC4F9FD",
    x"BEC4EE63",
    x"BEC4E2C9",
    x"BEC4D730",
    x"BEC4CB96",
    x"BEC4BFFC",
    x"BEC4B462",
    x"BEC4A8C8",
    x"BEC49D2E",
    x"BEC49193",
    x"BEC485F9",
    x"BEC47A5E",
    x"BEC46EC3",
    x"BEC46328",
    x"BEC4578D",
    x"BEC44BF2",
    x"BEC44057",
    x"BEC434BC",
    x"BEC42920",
    x"BEC41D85",
    x"BEC411E9",
    x"BEC4064D",
    x"BEC3FAB1",
    x"BEC3EF15",
    x"BEC3E379",
    x"BEC3D7DD",
    x"BEC3CC40",
    x"BEC3C0A4",
    x"BEC3B507",
    x"BEC3A96A",
    x"BEC39DCE",
    x"BEC39231",
    x"BEC38693",
    x"BEC37AF6",
    x"BEC36F59",
    x"BEC363BB",
    x"BEC3581E",
    x"BEC34C80",
    x"BEC340E2",
    x"BEC33544",
    x"BEC329A6",
    x"BEC31E08",
    x"BEC3126A",
    x"BEC306CB",
    x"BEC2FB2D",
    x"BEC2EF8E",
    x"BEC2E3EF",
    x"BEC2D851",
    x"BEC2CCB2",
    x"BEC2C112",
    x"BEC2B573",
    x"BEC2A9D4",
    x"BEC29E34",
    x"BEC29295",
    x"BEC286F5",
    x"BEC27B55",
    x"BEC26FB5",
    x"BEC26415",
    x"BEC25875",
    x"BEC24CD5",
    x"BEC24135",
    x"BEC23594",
    x"BEC229F3",
    x"BEC21E53",
    x"BEC212B2",
    x"BEC20711",
    x"BEC1FB70",
    x"BEC1EFCE",
    x"BEC1E42D",
    x"BEC1D88C",
    x"BEC1CCEA",
    x"BEC1C148",
    x"BEC1B5A7",
    x"BEC1AA05",
    x"BEC19E63",
    x"BEC192C0",
    x"BEC1871E",
    x"BEC17B7C",
    x"BEC16FD9",
    x"BEC16437",
    x"BEC15894",
    x"BEC14CF1",
    x"BEC1414E",
    x"BEC135AB",
    x"BEC12A08",
    x"BEC11E64",
    x"BEC112C1",
    x"BEC1071E",
    x"BEC0FB7A",
    x"BEC0EFD6",
    x"BEC0E432",
    x"BEC0D88E",
    x"BEC0CCEA",
    x"BEC0C146",
    x"BEC0B5A1",
    x"BEC0A9FD",
    x"BEC09E58",
    x"BEC092B4",
    x"BEC0870F",
    x"BEC07B6A",
    x"BEC06FC5",
    x"BEC06420",
    x"BEC0587A",
    x"BEC04CD5",
    x"BEC0412F",
    x"BEC0358A",
    x"BEC029E4",
    x"BEC01E3E",
    x"BEC01298",
    x"BEC006F2",
    x"BEBFFB4C",
    x"BEBFEFA5",
    x"BEBFE3FF",
    x"BEBFD858",
    x"BEBFCCB2",
    x"BEBFC10B",
    x"BEBFB564",
    x"BEBFA9BD",
    x"BEBF9E16",
    x"BEBF926F",
    x"BEBF86C7",
    x"BEBF7B20",
    x"BEBF6F78",
    x"BEBF63D0",
    x"BEBF5829",
    x"BEBF4C81",
    x"BEBF40D9",
    x"BEBF3530",
    x"BEBF2988",
    x"BEBF1DE0",
    x"BEBF1237",
    x"BEBF068F",
    x"BEBEFAE6",
    x"BEBEEF3D",
    x"BEBEE394",
    x"BEBED7EB",
    x"BEBECC42",
    x"BEBEC098",
    x"BEBEB4EF",
    x"BEBEA945",
    x"BEBE9D9C",
    x"BEBE91F2",
    x"BEBE8648",
    x"BEBE7A9E",
    x"BEBE6EF4",
    x"BEBE6349",
    x"BEBE579F",
    x"BEBE4BF5",
    x"BEBE404A",
    x"BEBE349F",
    x"BEBE28F4",
    x"BEBE1D4A",
    x"BEBE119E",
    x"BEBE05F3",
    x"BEBDFA48",
    x"BEBDEE9D",
    x"BEBDE2F1",
    x"BEBDD746",
    x"BEBDCB9A",
    x"BEBDBFEE",
    x"BEBDB442",
    x"BEBDA896",
    x"BEBD9CEA",
    x"BEBD913D",
    x"BEBD8591",
    x"BEBD79E4",
    x"BEBD6E38",
    x"BEBD628B",
    x"BEBD56DE",
    x"BEBD4B31",
    x"BEBD3F84",
    x"BEBD33D7",
    x"BEBD2829",
    x"BEBD1C7C",
    x"BEBD10CE",
    x"BEBD0521",
    x"BEBCF973",
    x"BEBCEDC5",
    x"BEBCE217",
    x"BEBCD669",
    x"BEBCCABB",
    x"BEBCBF0C",
    x"BEBCB35E",
    x"BEBCA7AF",
    x"BEBC9C00",
    x"BEBC9052",
    x"BEBC84A3",
    x"BEBC78F4",
    x"BEBC6D45",
    x"BEBC6195",
    x"BEBC55E6",
    x"BEBC4A36",
    x"BEBC3E87",
    x"BEBC32D7",
    x"BEBC2727",
    x"BEBC1B77",
    x"BEBC0FC7",
    x"BEBC0417",
    x"BEBBF867",
    x"BEBBECB6",
    x"BEBBE106",
    x"BEBBD555",
    x"BEBBC9A4",
    x"BEBBBDF4",
    x"BEBBB243",
    x"BEBBA692",
    x"BEBB9AE0",
    x"BEBB8F2F",
    x"BEBB837E",
    x"BEBB77CC",
    x"BEBB6C1A",
    x"BEBB6069",
    x"BEBB54B7",
    x"BEBB4905",
    x"BEBB3D53",
    x"BEBB31A0",
    x"BEBB25EE",
    x"BEBB1A3C",
    x"BEBB0E89",
    x"BEBB02D6",
    x"BEBAF724",
    x"BEBAEB71",
    x"BEBADFBE",
    x"BEBAD40B",
    x"BEBAC857",
    x"BEBABCA4",
    x"BEBAB0F1",
    x"BEBAA53D",
    x"BEBA9989",
    x"BEBA8DD6",
    x"BEBA8222",
    x"BEBA766E",
    x"BEBA6ABA",
    x"BEBA5F05",
    x"BEBA5351",
    x"BEBA479D",
    x"BEBA3BE8",
    x"BEBA3033",
    x"BEBA247F",
    x"BEBA18CA",
    x"BEBA0D15",
    x"BEBA015F",
    x"BEB9F5AA",
    x"BEB9E9F5",
    x"BEB9DE3F",
    x"BEB9D28A",
    x"BEB9C6D4",
    x"BEB9BB1E",
    x"BEB9AF68",
    x"BEB9A3B2",
    x"BEB997FC",
    x"BEB98C46",
    x"BEB98090",
    x"BEB974D9",
    x"BEB96923",
    x"BEB95D6C",
    x"BEB951B5",
    x"BEB945FE",
    x"BEB93A47",
    x"BEB92E90",
    x"BEB922D9",
    x"BEB91721",
    x"BEB90B6A",
    x"BEB8FFB2",
    x"BEB8F3FA",
    x"BEB8E843",
    x"BEB8DC8B",
    x"BEB8D0D3",
    x"BEB8C51B",
    x"BEB8B962",
    x"BEB8ADAA",
    x"BEB8A1F1",
    x"BEB89639",
    x"BEB88A80",
    x"BEB87EC7",
    x"BEB8730E",
    x"BEB86755",
    x"BEB85B9C",
    x"BEB84FE3",
    x"BEB8442A",
    x"BEB83870",
    x"BEB82CB6",
    x"BEB820FD",
    x"BEB81543",
    x"BEB80989",
    x"BEB7FDCF",
    x"BEB7F215",
    x"BEB7E65B",
    x"BEB7DAA0",
    x"BEB7CEE6",
    x"BEB7C32B",
    x"BEB7B770",
    x"BEB7ABB6",
    x"BEB79FFB",
    x"BEB79440",
    x"BEB78884",
    x"BEB77CC9",
    x"BEB7710E",
    x"BEB76552",
    x"BEB75997",
    x"BEB74DDB",
    x"BEB7421F",
    x"BEB73663",
    x"BEB72AA7",
    x"BEB71EEB",
    x"BEB7132F",
    x"BEB70773",
    x"BEB6FBB6",
    x"BEB6EFFA",
    x"BEB6E43D",
    x"BEB6D880",
    x"BEB6CCC3",
    x"BEB6C106",
    x"BEB6B549",
    x"BEB6A98C",
    x"BEB69DCE",
    x"BEB69211",
    x"BEB68653",
    x"BEB67A96",
    x"BEB66ED8",
    x"BEB6631A",
    x"BEB6575C",
    x"BEB64B9E",
    x"BEB63FE0",
    x"BEB63421",
    x"BEB62863",
    x"BEB61CA4",
    x"BEB610E6",
    x"BEB60527",
    x"BEB5F968",
    x"BEB5EDA9",
    x"BEB5E1EA",
    x"BEB5D62B",
    x"BEB5CA6B",
    x"BEB5BEAC",
    x"BEB5B2EC",
    x"BEB5A72D",
    x"BEB59B6D",
    x"BEB58FAD",
    x"BEB583ED",
    x"BEB5782D",
    x"BEB56C6D",
    x"BEB560AC",
    x"BEB554EC",
    x"BEB5492B",
    x"BEB53D6B",
    x"BEB531AA",
    x"BEB525E9",
    x"BEB51A28",
    x"BEB50E67",
    x"BEB502A6",
    x"BEB4F6E5",
    x"BEB4EB23",
    x"BEB4DF62",
    x"BEB4D3A0",
    x"BEB4C7DE",
    x"BEB4BC1D",
    x"BEB4B05B",
    x"BEB4A499",
    x"BEB498D6",
    x"BEB48D14",
    x"BEB48152",
    x"BEB4758F",
    x"BEB469CD",
    x"BEB45E0A",
    x"BEB45247",
    x"BEB44684",
    x"BEB43AC1",
    x"BEB42EFE",
    x"BEB4233B",
    x"BEB41777",
    x"BEB40BB4",
    x"BEB3FFF0",
    x"BEB3F42D",
    x"BEB3E869",
    x"BEB3DCA5",
    x"BEB3D0E1",
    x"BEB3C51D",
    x"BEB3B959",
    x"BEB3AD94",
    x"BEB3A1D0",
    x"BEB3960B",
    x"BEB38A47",
    x"BEB37E82",
    x"BEB372BD",
    x"BEB366F8",
    x"BEB35B33",
    x"BEB34F6E",
    x"BEB343A8",
    x"BEB337E3",
    x"BEB32C1D",
    x"BEB32058",
    x"BEB31492",
    x"BEB308CC",
    x"BEB2FD06",
    x"BEB2F140",
    x"BEB2E57A",
    x"BEB2D9B4",
    x"BEB2CDED",
    x"BEB2C227",
    x"BEB2B660",
    x"BEB2AA99",
    x"BEB29ED3",
    x"BEB2930C",
    x"BEB28745",
    x"BEB27B7E",
    x"BEB26FB6",
    x"BEB263EF",
    x"BEB25827",
    x"BEB24C60",
    x"BEB24098",
    x"BEB234D0",
    x"BEB22909",
    x"BEB21D41",
    x"BEB21178",
    x"BEB205B0",
    x"BEB1F9E8",
    x"BEB1EE1F",
    x"BEB1E257",
    x"BEB1D68E",
    x"BEB1CAC5",
    x"BEB1BEFD",
    x"BEB1B334",
    x"BEB1A76B",
    x"BEB19BA1",
    x"BEB18FD8",
    x"BEB1840F",
    x"BEB17845",
    x"BEB16C7C",
    x"BEB160B2",
    x"BEB154E8",
    x"BEB1491E",
    x"BEB13D54",
    x"BEB1318A",
    x"BEB125C0",
    x"BEB119F5",
    x"BEB10E2B",
    x"BEB10260",
    x"BEB0F696",
    x"BEB0EACB",
    x"BEB0DF00",
    x"BEB0D335",
    x"BEB0C76A",
    x"BEB0BB9F",
    x"BEB0AFD3",
    x"BEB0A408",
    x"BEB0983C",
    x"BEB08C71",
    x"BEB080A5",
    x"BEB074D9",
    x"BEB0690D",
    x"BEB05D41",
    x"BEB05175",
    x"BEB045A9",
    x"BEB039DC",
    x"BEB02E10",
    x"BEB02243",
    x"BEB01677",
    x"BEB00AAA",
    x"BEAFFEDD",
    x"BEAFF310",
    x"BEAFE743",
    x"BEAFDB76",
    x"BEAFCFA8",
    x"BEAFC3DB",
    x"BEAFB80D",
    x"BEAFAC40",
    x"BEAFA072",
    x"BEAF94A4",
    x"BEAF88D6",
    x"BEAF7D08",
    x"BEAF713A",
    x"BEAF656B",
    x"BEAF599D",
    x"BEAF4DCF",
    x"BEAF4200",
    x"BEAF3631",
    x"BEAF2A62",
    x"BEAF1E94",
    x"BEAF12C5",
    x"BEAF06F5",
    x"BEAEFB26",
    x"BEAEEF57",
    x"BEAEE387",
    x"BEAED7B8",
    x"BEAECBE8",
    x"BEAEC018",
    x"BEAEB449",
    x"BEAEA879",
    x"BEAE9CA8",
    x"BEAE90D8",
    x"BEAE8508",
    x"BEAE7938",
    x"BEAE6D67",
    x"BEAE6197",
    x"BEAE55C6",
    x"BEAE49F5",
    x"BEAE3E24",
    x"BEAE3253",
    x"BEAE2682",
    x"BEAE1AB1",
    x"BEAE0EDF",
    x"BEAE030E",
    x"BEADF73C",
    x"BEADEB6B",
    x"BEADDF99",
    x"BEADD3C7",
    x"BEADC7F5",
    x"BEADBC23",
    x"BEADB051",
    x"BEADA47F",
    x"BEAD98AC",
    x"BEAD8CDA",
    x"BEAD8107",
    x"BEAD7534",
    x"BEAD6962",
    x"BEAD5D8F",
    x"BEAD51BC",
    x"BEAD45E9",
    x"BEAD3A15",
    x"BEAD2E42",
    x"BEAD226F",
    x"BEAD169B",
    x"BEAD0AC7",
    x"BEACFEF4",
    x"BEACF320",
    x"BEACE74C",
    x"BEACDB78",
    x"BEACCFA4",
    x"BEACC3CF",
    x"BEACB7FB",
    x"BEACAC27",
    x"BEACA052",
    x"BEAC947D",
    x"BEAC88A9",
    x"BEAC7CD4",
    x"BEAC70FF",
    x"BEAC652A",
    x"BEAC5954",
    x"BEAC4D7F",
    x"BEAC41AA",
    x"BEAC35D4",
    x"BEAC29FF",
    x"BEAC1E29",
    x"BEAC1253",
    x"BEAC067D",
    x"BEABFAA7",
    x"BEABEED1",
    x"BEABE2FB",
    x"BEABD724",
    x"BEABCB4E",
    x"BEABBF77",
    x"BEABB3A1",
    x"BEABA7CA",
    x"BEAB9BF3",
    x"BEAB901C",
    x"BEAB8445",
    x"BEAB786E",
    x"BEAB6C97",
    x"BEAB60BF",
    x"BEAB54E8",
    x"BEAB4910",
    x"BEAB3D39",
    x"BEAB3161",
    x"BEAB2589",
    x"BEAB19B1",
    x"BEAB0DD9",
    x"BEAB0201",
    x"BEAAF628",
    x"BEAAEA50",
    x"BEAADE77",
    x"BEAAD29F",
    x"BEAAC6C6",
    x"BEAABAED",
    x"BEAAAF14",
    x"BEAAA33B",
    x"BEAA9762",
    x"BEAA8B89",
    x"BEAA7FB0",
    x"BEAA73D6",
    x"BEAA67FD",
    x"BEAA5C23",
    x"BEAA5049",
    x"BEAA446F",
    x"BEAA3895",
    x"BEAA2CBB",
    x"BEAA20E1",
    x"BEAA1507",
    x"BEAA092D",
    x"BEA9FD52",
    x"BEA9F178",
    x"BEA9E59D",
    x"BEA9D9C2",
    x"BEA9CDE7",
    x"BEA9C20C",
    x"BEA9B631",
    x"BEA9AA56",
    x"BEA99E7B",
    x"BEA992A0",
    x"BEA986C4",
    x"BEA97AE8",
    x"BEA96F0D",
    x"BEA96331",
    x"BEA95755",
    x"BEA94B79",
    x"BEA93F9D",
    x"BEA933C1",
    x"BEA927E5",
    x"BEA91C08",
    x"BEA9102C",
    x"BEA9044F",
    x"BEA8F872",
    x"BEA8EC95",
    x"BEA8E0B9",
    x"BEA8D4DC",
    x"BEA8C8FE",
    x"BEA8BD21",
    x"BEA8B144",
    x"BEA8A567",
    x"BEA89989",
    x"BEA88DAB",
    x"BEA881CE",
    x"BEA875F0",
    x"BEA86A12",
    x"BEA85E34",
    x"BEA85256",
    x"BEA84678",
    x"BEA83A99",
    x"BEA82EBB",
    x"BEA822DC",
    x"BEA816FE",
    x"BEA80B1F",
    x"BEA7FF40",
    x"BEA7F361",
    x"BEA7E782",
    x"BEA7DBA3",
    x"BEA7CFC4",
    x"BEA7C3E4",
    x"BEA7B805",
    x"BEA7AC25",
    x"BEA7A046",
    x"BEA79466",
    x"BEA78886",
    x"BEA77CA6",
    x"BEA770C6",
    x"BEA764E6",
    x"BEA75906",
    x"BEA74D25",
    x"BEA74145",
    x"BEA73564",
    x"BEA72984",
    x"BEA71DA3",
    x"BEA711C2",
    x"BEA705E1",
    x"BEA6FA00",
    x"BEA6EE1F",
    x"BEA6E23E",
    x"BEA6D65C",
    x"BEA6CA7B",
    x"BEA6BE99",
    x"BEA6B2B8",
    x"BEA6A6D6",
    x"BEA69AF4",
    x"BEA68F12",
    x"BEA68330",
    x"BEA6774E",
    x"BEA66B6C",
    x"BEA65F89",
    x"BEA653A7",
    x"BEA647C4",
    x"BEA63BE2",
    x"BEA62FFF",
    x"BEA6241C",
    x"BEA61839",
    x"BEA60C56",
    x"BEA60073",
    x"BEA5F48F",
    x"BEA5E8AC",
    x"BEA5DCC9",
    x"BEA5D0E5",
    x"BEA5C501",
    x"BEA5B91E",
    x"BEA5AD3A",
    x"BEA5A156",
    x"BEA59572",
    x"BEA5898E",
    x"BEA57DA9",
    x"BEA571C5",
    x"BEA565E1",
    x"BEA559FC",
    x"BEA54E17",
    x"BEA54233",
    x"BEA5364E",
    x"BEA52A69",
    x"BEA51E84",
    x"BEA5129F",
    x"BEA506B9",
    x"BEA4FAD4",
    x"BEA4EEEE",
    x"BEA4E309",
    x"BEA4D723",
    x"BEA4CB3E",
    x"BEA4BF58",
    x"BEA4B372",
    x"BEA4A78C",
    x"BEA49BA6",
    x"BEA48FBF",
    x"BEA483D9",
    x"BEA477F2",
    x"BEA46C0C",
    x"BEA46025",
    x"BEA4543F",
    x"BEA44858",
    x"BEA43C71",
    x"BEA4308A",
    x"BEA424A3",
    x"BEA418BB",
    x"BEA40CD4",
    x"BEA400ED",
    x"BEA3F505",
    x"BEA3E91D",
    x"BEA3DD36",
    x"BEA3D14E",
    x"BEA3C566",
    x"BEA3B97E",
    x"BEA3AD96",
    x"BEA3A1AD",
    x"BEA395C5",
    x"BEA389DD",
    x"BEA37DF4",
    x"BEA3720C",
    x"BEA36623",
    x"BEA35A3A",
    x"BEA34E51",
    x"BEA34268",
    x"BEA3367F",
    x"BEA32A96",
    x"BEA31EAD",
    x"BEA312C3",
    x"BEA306DA",
    x"BEA2FAF0",
    x"BEA2EF06",
    x"BEA2E31C",
    x"BEA2D733",
    x"BEA2CB49",
    x"BEA2BF5E",
    x"BEA2B374",
    x"BEA2A78A",
    x"BEA29BA0",
    x"BEA28FB5",
    x"BEA283CB",
    x"BEA277E0",
    x"BEA26BF5",
    x"BEA2600A",
    x"BEA2541F",
    x"BEA24834",
    x"BEA23C49",
    x"BEA2305E",
    x"BEA22472",
    x"BEA21887",
    x"BEA20C9B",
    x"BEA200B0",
    x"BEA1F4C4",
    x"BEA1E8D8",
    x"BEA1DCEC",
    x"BEA1D100",
    x"BEA1C514",
    x"BEA1B928",
    x"BEA1AD3B",
    x"BEA1A14F",
    x"BEA19562",
    x"BEA18976",
    x"BEA17D89",
    x"BEA1719C",
    x"BEA165AF",
    x"BEA159C2",
    x"BEA14DD5",
    x"BEA141E8",
    x"BEA135FB",
    x"BEA12A0D",
    x"BEA11E20",
    x"BEA11232",
    x"BEA10644",
    x"BEA0FA57",
    x"BEA0EE69",
    x"BEA0E27B",
    x"BEA0D68D",
    x"BEA0CA9E",
    x"BEA0BEB0",
    x"BEA0B2C2",
    x"BEA0A6D3",
    x"BEA09AE5",
    x"BEA08EF6",
    x"BEA08307",
    x"BEA07718",
    x"BEA06B29",
    x"BEA05F3A",
    x"BEA0534B",
    x"BEA0475C",
    x"BEA03B6D",
    x"BEA02F7D",
    x"BEA0238E",
    x"BEA0179E",
    x"BEA00BAE",
    x"BE9FFFBE",
    x"BE9FF3CE",
    x"BE9FE7DE",
    x"BE9FDBEE",
    x"BE9FCFFE",
    x"BE9FC40E",
    x"BE9FB81D",
    x"BE9FAC2D",
    x"BE9FA03C",
    x"BE9F944C",
    x"BE9F885B",
    x"BE9F7C6A",
    x"BE9F7079",
    x"BE9F6488",
    x"BE9F5897",
    x"BE9F4CA5",
    x"BE9F40B4",
    x"BE9F34C3",
    x"BE9F28D1",
    x"BE9F1CDF",
    x"BE9F10EE",
    x"BE9F04FC",
    x"BE9EF90A",
    x"BE9EED18",
    x"BE9EE126",
    x"BE9ED533",
    x"BE9EC941",
    x"BE9EBD4F",
    x"BE9EB15C",
    x"BE9EA569",
    x"BE9E9977",
    x"BE9E8D84",
    x"BE9E8191",
    x"BE9E759E",
    x"BE9E69AB",
    x"BE9E5DB8",
    x"BE9E51C4",
    x"BE9E45D1",
    x"BE9E39DE",
    x"BE9E2DEA",
    x"BE9E21F6",
    x"BE9E1603",
    x"BE9E0A0F",
    x"BE9DFE1B",
    x"BE9DF227",
    x"BE9DE633",
    x"BE9DDA3E",
    x"BE9DCE4A",
    x"BE9DC256",
    x"BE9DB661",
    x"BE9DAA6D",
    x"BE9D9E78",
    x"BE9D9283",
    x"BE9D868E",
    x"BE9D7A99",
    x"BE9D6EA4",
    x"BE9D62AF",
    x"BE9D56BA",
    x"BE9D4AC4",
    x"BE9D3ECF",
    x"BE9D32D9",
    x"BE9D26E3",
    x"BE9D1AEE",
    x"BE9D0EF8",
    x"BE9D0302",
    x"BE9CF70C",
    x"BE9CEB16",
    x"BE9CDF20",
    x"BE9CD329",
    x"BE9CC733",
    x"BE9CBB3C",
    x"BE9CAF46",
    x"BE9CA34F",
    x"BE9C9758",
    x"BE9C8B61",
    x"BE9C7F6A",
    x"BE9C7373",
    x"BE9C677C",
    x"BE9C5B85",
    x"BE9C4F8D",
    x"BE9C4396",
    x"BE9C379E",
    x"BE9C2BA7",
    x"BE9C1FAF",
    x"BE9C13B7",
    x"BE9C07BF",
    x"BE9BFBC7",
    x"BE9BEFCF",
    x"BE9BE3D7",
    x"BE9BD7DF",
    x"BE9BCBE6",
    x"BE9BBFEE",
    x"BE9BB3F5",
    x"BE9BA7FD",
    x"BE9B9C04",
    x"BE9B900B",
    x"BE9B8412",
    x"BE9B7819",
    x"BE9B6C20",
    x"BE9B6027",
    x"BE9B542D",
    x"BE9B4834",
    x"BE9B3C3A",
    x"BE9B3041",
    x"BE9B2447",
    x"BE9B184D",
    x"BE9B0C53",
    x"BE9B0059",
    x"BE9AF45F",
    x"BE9AE865",
    x"BE9ADC6B",
    x"BE9AD070",
    x"BE9AC476",
    x"BE9AB87B",
    x"BE9AAC81",
    x"BE9AA086",
    x"BE9A948B",
    x"BE9A8890",
    x"BE9A7C95",
    x"BE9A709A",
    x"BE9A649F",
    x"BE9A58A4",
    x"BE9A4CA8",
    x"BE9A40AD",
    x"BE9A34B1",
    x"BE9A28B6",
    x"BE9A1CBA",
    x"BE9A10BE",
    x"BE9A04C2",
    x"BE99F8C6",
    x"BE99ECCA",
    x"BE99E0CE",
    x"BE99D4D1",
    x"BE99C8D5",
    x"BE99BCD9",
    x"BE99B0DC",
    x"BE99A4DF",
    x"BE9998E3",
    x"BE998CE6",
    x"BE9980E9",
    x"BE9974EC",
    x"BE9968EE",
    x"BE995CF1",
    x"BE9950F4",
    x"BE9944F7",
    x"BE9938F9",
    x"BE992CFB",
    x"BE9920FE",
    x"BE991500",
    x"BE990902",
    x"BE98FD04",
    x"BE98F106",
    x"BE98E508",
    x"BE98D90A",
    x"BE98CD0B",
    x"BE98C10D",
    x"BE98B50E",
    x"BE98A910",
    x"BE989D11",
    x"BE989112",
    x"BE988513",
    x"BE987914",
    x"BE986D15",
    x"BE986116",
    x"BE985517",
    x"BE984917",
    x"BE983D18",
    x"BE983118",
    x"BE982519",
    x"BE981919",
    x"BE980D19",
    x"BE980119",
    x"BE97F519",
    x"BE97E919",
    x"BE97DD19",
    x"BE97D119",
    x"BE97C518",
    x"BE97B918",
    x"BE97AD17",
    x"BE97A117",
    x"BE979516",
    x"BE978915",
    x"BE977D14",
    x"BE977113",
    x"BE976512",
    x"BE975911",
    x"BE974D10",
    x"BE97410E",
    x"BE97350D",
    x"BE97290B",
    x"BE971D0A",
    x"BE971108",
    x"BE970506",
    x"BE96F904",
    x"BE96ED02",
    x"BE96E100",
    x"BE96D4FE",
    x"BE96C8FC",
    x"BE96BCF9",
    x"BE96B0F7",
    x"BE96A4F4",
    x"BE9698F2",
    x"BE968CEF",
    x"BE9680EC",
    x"BE9674E9",
    x"BE9668E6",
    x"BE965CE3",
    x"BE9650E0",
    x"BE9644DD",
    x"BE9638D9",
    x"BE962CD6",
    x"BE9620D2",
    x"BE9614CF",
    x"BE9608CB",
    x"BE95FCC7",
    x"BE95F0C3",
    x"BE95E4BF",
    x"BE95D8BB",
    x"BE95CCB7",
    x"BE95C0B3",
    x"BE95B4AE",
    x"BE95A8AA",
    x"BE959CA6",
    x"BE9590A1",
    x"BE95849C",
    x"BE957897",
    x"BE956C92",
    x"BE95608D",
    x"BE955488",
    x"BE954883",
    x"BE953C7E",
    x"BE953079",
    x"BE952473",
    x"BE95186E",
    x"BE950C68",
    x"BE950062",
    x"BE94F45D",
    x"BE94E857",
    x"BE94DC51",
    x"BE94D04B",
    x"BE94C444",
    x"BE94B83E",
    x"BE94AC38",
    x"BE94A031",
    x"BE94942B",
    x"BE948824",
    x"BE947C1E",
    x"BE947017",
    x"BE946410",
    x"BE945809",
    x"BE944C02",
    x"BE943FFB",
    x"BE9433F4",
    x"BE9427EC",
    x"BE941BE5",
    x"BE940FDD",
    x"BE9403D6",
    x"BE93F7CE",
    x"BE93EBC6",
    x"BE93DFBF",
    x"BE93D3B7",
    x"BE93C7AF",
    x"BE93BBA6",
    x"BE93AF9E",
    x"BE93A396",
    x"BE93978E",
    x"BE938B85",
    x"BE937F7D",
    x"BE937374",
    x"BE93676B",
    x"BE935B62",
    x"BE934F59",
    x"BE934350",
    x"BE933747",
    x"BE932B3E",
    x"BE931F35",
    x"BE93132B",
    x"BE930722",
    x"BE92FB18",
    x"BE92EF0F",
    x"BE92E305",
    x"BE92D6FB",
    x"BE92CAF1",
    x"BE92BEE7",
    x"BE92B2DD",
    x"BE92A6D3",
    x"BE929AC9",
    x"BE928EBF",
    x"BE9282B4",
    x"BE9276AA",
    x"BE926A9F",
    x"BE925E94",
    x"BE92528A",
    x"BE92467F",
    x"BE923A74",
    x"BE922E69",
    x"BE92225E",
    x"BE921652",
    x"BE920A47",
    x"BE91FE3C",
    x"BE91F230",
    x"BE91E625",
    x"BE91DA19",
    x"BE91CE0D",
    x"BE91C201",
    x"BE91B5F5",
    x"BE91A9E9",
    x"BE919DDD",
    x"BE9191D1",
    x"BE9185C5",
    x"BE9179B9",
    x"BE916DAC",
    x"BE9161A0",
    x"BE915593",
    x"BE914986",
    x"BE913D79",
    x"BE91316D",
    x"BE912560",
    x"BE911953",
    x"BE910D45",
    x"BE910138",
    x"BE90F52B",
    x"BE90E91D",
    x"BE90DD10",
    x"BE90D102",
    x"BE90C4F5",
    x"BE90B8E7",
    x"BE90ACD9",
    x"BE90A0CB",
    x"BE9094BD",
    x"BE9088AF",
    x"BE907CA1",
    x"BE907093",
    x"BE906484",
    x"BE905876",
    x"BE904C67",
    x"BE904059",
    x"BE90344A",
    x"BE90283B",
    x"BE901C2C",
    x"BE90101D",
    x"BE90040E",
    x"BE8FF7FF",
    x"BE8FEBF0",
    x"BE8FDFE0",
    x"BE8FD3D1",
    x"BE8FC7C1",
    x"BE8FBBB2",
    x"BE8FAFA2",
    x"BE8FA392",
    x"BE8F9783",
    x"BE8F8B73",
    x"BE8F7F63",
    x"BE8F7353",
    x"BE8F6742",
    x"BE8F5B32",
    x"BE8F4F22",
    x"BE8F4311",
    x"BE8F3701",
    x"BE8F2AF0",
    x"BE8F1EDF",
    x"BE8F12CF",
    x"BE8F06BE",
    x"BE8EFAAD",
    x"BE8EEE9C",
    x"BE8EE28B",
    x"BE8ED679",
    x"BE8ECA68",
    x"BE8EBE57",
    x"BE8EB245",
    x"BE8EA634",
    x"BE8E9A22",
    x"BE8E8E10",
    x"BE8E81FE",
    x"BE8E75ED",
    x"BE8E69DB",
    x"BE8E5DC8",
    x"BE8E51B6",
    x"BE8E45A4",
    x"BE8E3992",
    x"BE8E2D7F",
    x"BE8E216D",
    x"BE8E155A",
    x"BE8E0947",
    x"BE8DFD35",
    x"BE8DF122",
    x"BE8DE50F",
    x"BE8DD8FC",
    x"BE8DCCE9",
    x"BE8DC0D6",
    x"BE8DB4C2",
    x"BE8DA8AF",
    x"BE8D9C9B",
    x"BE8D9088",
    x"BE8D8474",
    x"BE8D7861",
    x"BE8D6C4D",
    x"BE8D6039",
    x"BE8D5425",
    x"BE8D4811",
    x"BE8D3BFD",
    x"BE8D2FE9",
    x"BE8D23D4",
    x"BE8D17C0",
    x"BE8D0BAB",
    x"BE8CFF97",
    x"BE8CF382",
    x"BE8CE76D",
    x"BE8CDB59",
    x"BE8CCF44",
    x"BE8CC32F",
    x"BE8CB71A",
    x"BE8CAB05",
    x"BE8C9EEF",
    x"BE8C92DA",
    x"BE8C86C5",
    x"BE8C7AAF",
    x"BE8C6E9A",
    x"BE8C6284",
    x"BE8C566E",
    x"BE8C4A58",
    x"BE8C3E42",
    x"BE8C322C",
    x"BE8C2616",
    x"BE8C1A00",
    x"BE8C0DEA",
    x"BE8C01D4",
    x"BE8BF5BD",
    x"BE8BE9A7",
    x"BE8BDD90",
    x"BE8BD179",
    x"BE8BC563",
    x"BE8BB94C",
    x"BE8BAD35",
    x"BE8BA11E",
    x"BE8B9507",
    x"BE8B88F0",
    x"BE8B7CD8",
    x"BE8B70C1",
    x"BE8B64AA",
    x"BE8B5892",
    x"BE8B4C7A",
    x"BE8B4063",
    x"BE8B344B",
    x"BE8B2833",
    x"BE8B1C1B",
    x"BE8B1003",
    x"BE8B03EB",
    x"BE8AF7D3",
    x"BE8AEBBB",
    x"BE8ADFA2",
    x"BE8AD38A",
    x"BE8AC771",
    x"BE8ABB59",
    x"BE8AAF40",
    x"BE8AA327",
    x"BE8A970E",
    x"BE8A8AF5",
    x"BE8A7EDC",
    x"BE8A72C3",
    x"BE8A66AA",
    x"BE8A5A91",
    x"BE8A4E78",
    x"BE8A425E",
    x"BE8A3645",
    x"BE8A2A2B",
    x"BE8A1E11",
    x"BE8A11F7",
    x"BE8A05DE",
    x"BE89F9C4",
    x"BE89EDAA",
    x"BE89E190",
    x"BE89D575",
    x"BE89C95B",
    x"BE89BD41",
    x"BE89B126",
    x"BE89A50C",
    x"BE8998F1",
    x"BE898CD7",
    x"BE8980BC",
    x"BE8974A1",
    x"BE896886",
    x"BE895C6B",
    x"BE895050",
    x"BE894435",
    x"BE893819",
    x"BE892BFE",
    x"BE891FE3",
    x"BE8913C7",
    x"BE8907AC",
    x"BE88FB90",
    x"BE88EF74",
    x"BE88E358",
    x"BE88D73C",
    x"BE88CB20",
    x"BE88BF04",
    x"BE88B2E8",
    x"BE88A6CC",
    x"BE889AB0",
    x"BE888E93",
    x"BE888277",
    x"BE88765A",
    x"BE886A3D",
    x"BE885E21",
    x"BE885204",
    x"BE8845E7",
    x"BE8839CA",
    x"BE882DAD",
    x"BE882190",
    x"BE881572",
    x"BE880955",
    x"BE87FD38",
    x"BE87F11A",
    x"BE87E4FD",
    x"BE87D8DF",
    x"BE87CCC1",
    x"BE87C0A3",
    x"BE87B486",
    x"BE87A868",
    x"BE879C49",
    x"BE87902B",
    x"BE87840D",
    x"BE8777EF",
    x"BE876BD0",
    x"BE875FB2",
    x"BE875393",
    x"BE874775",
    x"BE873B56",
    x"BE872F37",
    x"BE872318",
    x"BE8716F9",
    x"BE870ADA",
    x"BE86FEBB",
    x"BE86F29C",
    x"BE86E67D",
    x"BE86DA5D",
    x"BE86CE3E",
    x"BE86C21F",
    x"BE86B5FF",
    x"BE86A9DF",
    x"BE869DBF",
    x"BE8691A0",
    x"BE868580",
    x"BE867960",
    x"BE866D40",
    x"BE86611F",
    x"BE8654FF",
    x"BE8648DF",
    x"BE863CBE",
    x"BE86309E",
    x"BE86247D",
    x"BE86185D",
    x"BE860C3C",
    x"BE86001B",
    x"BE85F3FA",
    x"BE85E7D9",
    x"BE85DBB8",
    x"BE85CF97",
    x"BE85C376",
    x"BE85B755",
    x"BE85AB33",
    x"BE859F12",
    x"BE8592F0",
    x"BE8586CE",
    x"BE857AAD",
    x"BE856E8B",
    x"BE856269",
    x"BE855647",
    x"BE854A25",
    x"BE853E03",
    x"BE8531E1",
    x"BE8525BF",
    x"BE85199C",
    x"BE850D7A",
    x"BE850157",
    x"BE84F535",
    x"BE84E912",
    x"BE84DCEF",
    x"BE84D0CC",
    x"BE84C4AA",
    x"BE84B887",
    x"BE84AC64",
    x"BE84A040",
    x"BE84941D",
    x"BE8487FA",
    x"BE847BD6",
    x"BE846FB3",
    x"BE84638F",
    x"BE84576C",
    x"BE844B48",
    x"BE843F24",
    x"BE843300",
    x"BE8426DD",
    x"BE841AB8",
    x"BE840E94",
    x"BE840270",
    x"BE83F64C",
    x"BE83EA28",
    x"BE83DE03",
    x"BE83D1DF",
    x"BE83C5BA",
    x"BE83B995",
    x"BE83AD71",
    x"BE83A14C",
    x"BE839527",
    x"BE838902",
    x"BE837CDD",
    x"BE8370B8",
    x"BE836493",
    x"BE83586D",
    x"BE834C48",
    x"BE834022",
    x"BE8333FD",
    x"BE8327D7",
    x"BE831BB2",
    x"BE830F8C",
    x"BE830366",
    x"BE82F740",
    x"BE82EB1A",
    x"BE82DEF4",
    x"BE82D2CE",
    x"BE82C6A8",
    x"BE82BA81",
    x"BE82AE5B",
    x"BE82A234",
    x"BE82960E",
    x"BE8289E7",
    x"BE827DC0",
    x"BE82719A",
    x"BE826573",
    x"BE82594C",
    x"BE824D25",
    x"BE8240FE",
    x"BE8234D7",
    x"BE8228AF",
    x"BE821C88",
    x"BE821060",
    x"BE820439",
    x"BE81F811",
    x"BE81EBEA",
    x"BE81DFC2",
    x"BE81D39A",
    x"BE81C772",
    x"BE81BB4A",
    x"BE81AF22",
    x"BE81A2FA",
    x"BE8196D2",
    x"BE818AAA",
    x"BE817E81",
    x"BE817259",
    x"BE816630",
    x"BE815A08",
    x"BE814DDF",
    x"BE8141B6",
    x"BE81358E",
    x"BE812965",
    x"BE811D3C",
    x"BE811113",
    x"BE8104E9",
    x"BE80F8C0",
    x"BE80EC97",
    x"BE80E06E",
    x"BE80D444",
    x"BE80C81B",
    x"BE80BBF1",
    x"BE80AFC7",
    x"BE80A39E",
    x"BE809774",
    x"BE808B4A",
    x"BE807F20",
    x"BE8072F6",
    x"BE8066CC",
    x"BE805AA1",
    x"BE804E77",
    x"BE80424D",
    x"BE803622",
    x"BE8029F8",
    x"BE801DCD",
    x"BE8011A2",
    x"BE800578",
    x"BE7FF29A",
    x"BE7FDA44",
    x"BE7FC1EE",
    x"BE7FA998",
    x"BE7F9141",
    x"BE7F78EB",
    x"BE7F6094",
    x"BE7F483D",
    x"BE7F2FE7",
    x"BE7F178F",
    x"BE7EFF38",
    x"BE7EE6E1",
    x"BE7ECE89",
    x"BE7EB632",
    x"BE7E9DDA",
    x"BE7E8582",
    x"BE7E6D2A",
    x"BE7E54D1",
    x"BE7E3C79",
    x"BE7E2420",
    x"BE7E0BC8",
    x"BE7DF36F",
    x"BE7DDB16",
    x"BE7DC2BC",
    x"BE7DAA63",
    x"BE7D9209",
    x"BE7D79B0",
    x"BE7D6156",
    x"BE7D48FC",
    x"BE7D30A2",
    x"BE7D1848",
    x"BE7CFFED",
    x"BE7CE793",
    x"BE7CCF38",
    x"BE7CB6DD",
    x"BE7C9E82",
    x"BE7C8627",
    x"BE7C6DCB",
    x"BE7C5570",
    x"BE7C3D14",
    x"BE7C24B8",
    x"BE7C0C5C",
    x"BE7BF400",
    x"BE7BDBA4",
    x"BE7BC348",
    x"BE7BAAEB",
    x"BE7B928E",
    x"BE7B7A31",
    x"BE7B61D4",
    x"BE7B4977",
    x"BE7B311A",
    x"BE7B18BC",
    x"BE7B005F",
    x"BE7AE801",
    x"BE7ACFA3",
    x"BE7AB745",
    x"BE7A9EE7",
    x"BE7A8688",
    x"BE7A6E2A",
    x"BE7A55CB",
    x"BE7A3D6C",
    x"BE7A250D",
    x"BE7A0CAE",
    x"BE79F44F",
    x"BE79DBF0",
    x"BE79C390",
    x"BE79AB30",
    x"BE7992D0",
    x"BE797A70",
    x"BE796210",
    x"BE7949B0",
    x"BE79314F",
    x"BE7918EF",
    x"BE79008E",
    x"BE78E82D",
    x"BE78CFCC",
    x"BE78B76B",
    x"BE789F09",
    x"BE7886A8",
    x"BE786E46",
    x"BE7855E4",
    x"BE783D82",
    x"BE782520",
    x"BE780CBE",
    x"BE77F45B",
    x"BE77DBF9",
    x"BE77C396",
    x"BE77AB33",
    x"BE7792D0",
    x"BE777A6D",
    x"BE77620A",
    x"BE7749A6",
    x"BE773142",
    x"BE7718DF",
    x"BE77007B",
    x"BE76E817",
    x"BE76CFB2",
    x"BE76B74E",
    x"BE769EEA",
    x"BE768685",
    x"BE766E20",
    x"BE7655BB",
    x"BE763D56",
    x"BE7624F1",
    x"BE760C8B",
    x"BE75F426",
    x"BE75DBC0",
    x"BE75C35A",
    x"BE75AAF4",
    x"BE75928E",
    x"BE757A28",
    x"BE7561C1",
    x"BE75495B",
    x"BE7530F4",
    x"BE75188D",
    x"BE750026",
    x"BE74E7BF",
    x"BE74CF57",
    x"BE74B6F0",
    x"BE749E88",
    x"BE748621",
    x"BE746DB9",
    x"BE745551",
    x"BE743CE8",
    x"BE742480",
    x"BE740C18",
    x"BE73F3AF",
    x"BE73DB46",
    x"BE73C2DD",
    x"BE73AA74",
    x"BE73920B",
    x"BE7379A1",
    x"BE736138",
    x"BE7348CE",
    x"BE733064",
    x"BE7317FA",
    x"BE72FF90",
    x"BE72E726",
    x"BE72CEBC",
    x"BE72B651",
    x"BE729DE6",
    x"BE72857B",
    x"BE726D10",
    x"BE7254A5",
    x"BE723C3A",
    x"BE7223CE",
    x"BE720B63",
    x"BE71F2F7",
    x"BE71DA8B",
    x"BE71C21F",
    x"BE71A9B3",
    x"BE719147",
    x"BE7178DA",
    x"BE71606E",
    x"BE714801",
    x"BE712F94",
    x"BE711727",
    x"BE70FEBA",
    x"BE70E64C",
    x"BE70CDDF",
    x"BE70B571",
    x"BE709D04",
    x"BE708496",
    x"BE706C28",
    x"BE7053B9",
    x"BE703B4B",
    x"BE7022DD",
    x"BE700A6E",
    x"BE6FF1FF",
    x"BE6FD990",
    x"BE6FC121",
    x"BE6FA8B2",
    x"BE6F9043",
    x"BE6F77D3",
    x"BE6F5F63",
    x"BE6F46F4",
    x"BE6F2E84",
    x"BE6F1614",
    x"BE6EFDA3",
    x"BE6EE533",
    x"BE6ECCC3",
    x"BE6EB452",
    x"BE6E9BE1",
    x"BE6E8370",
    x"BE6E6AFF",
    x"BE6E528E",
    x"BE6E3A1C",
    x"BE6E21AB",
    x"BE6E0939",
    x"BE6DF0C7",
    x"BE6DD856",
    x"BE6DBFE3",
    x"BE6DA771",
    x"BE6D8EFF",
    x"BE6D768C",
    x"BE6D5E1A",
    x"BE6D45A7",
    x"BE6D2D34",
    x"BE6D14C1",
    x"BE6CFC4E",
    x"BE6CE3DA",
    x"BE6CCB67",
    x"BE6CB2F3",
    x"BE6C9A7F",
    x"BE6C820B",
    x"BE6C6997",
    x"BE6C5123",
    x"BE6C38AF",
    x"BE6C203A",
    x"BE6C07C5",
    x"BE6BEF51",
    x"BE6BD6DC",
    x"BE6BBE66",
    x"BE6BA5F1",
    x"BE6B8D7C",
    x"BE6B7506",
    x"BE6B5C91",
    x"BE6B441B",
    x"BE6B2BA5",
    x"BE6B132F",
    x"BE6AFAB9",
    x"BE6AE242",
    x"BE6AC9CC",
    x"BE6AB155",
    x"BE6A98DE",
    x"BE6A8067",
    x"BE6A67F0",
    x"BE6A4F79",
    x"BE6A3702",
    x"BE6A1E8A",
    x"BE6A0613",
    x"BE69ED9B",
    x"BE69D523",
    x"BE69BCAB",
    x"BE69A433",
    x"BE698BBA",
    x"BE697342",
    x"BE695AC9",
    x"BE694251",
    x"BE6929D8",
    x"BE69115F",
    x"BE68F8E5",
    x"BE68E06C",
    x"BE68C7F3",
    x"BE68AF79",
    x"BE6896FF",
    x"BE687E85",
    x"BE68660B",
    x"BE684D91",
    x"BE683517",
    x"BE681C9C",
    x"BE680422",
    x"BE67EBA7",
    x"BE67D32C",
    x"BE67BAB1",
    x"BE67A236",
    x"BE6789BB",
    x"BE67713F",
    x"BE6758C4",
    x"BE674048",
    x"BE6727CC",
    x"BE670F50",
    x"BE66F6D4",
    x"BE66DE58",
    x"BE66C5DC",
    x"BE66AD5F",
    x"BE6694E2",
    x"BE667C66",
    x"BE6663E9",
    x"BE664B6C",
    x"BE6632EE",
    x"BE661A71",
    x"BE6601F3",
    x"BE65E976",
    x"BE65D0F8",
    x"BE65B87A",
    x"BE659FFC",
    x"BE65877E",
    x"BE656F00",
    x"BE655681",
    x"BE653E02",
    x"BE652584",
    x"BE650D05",
    x"BE64F486",
    x"BE64DC07",
    x"BE64C387",
    x"BE64AB08",
    x"BE649288",
    x"BE647A09",
    x"BE646189",
    x"BE644909",
    x"BE643089",
    x"BE641808",
    x"BE63FF88",
    x"BE63E707",
    x"BE63CE87",
    x"BE63B606",
    x"BE639D85",
    x"BE638504",
    x"BE636C83",
    x"BE635401",
    x"BE633B80",
    x"BE6322FE",
    x"BE630A7C",
    x"BE62F1FA",
    x"BE62D978",
    x"BE62C0F6",
    x"BE62A874",
    x"BE628FF1",
    x"BE62776F",
    x"BE625EEC",
    x"BE624669",
    x"BE622DE6",
    x"BE621563",
    x"BE61FCE0",
    x"BE61E45C",
    x"BE61CBD9",
    x"BE61B355",
    x"BE619AD1",
    x"BE61824D",
    x"BE6169C9",
    x"BE615145",
    x"BE6138C1",
    x"BE61203C",
    x"BE6107B8",
    x"BE60EF33",
    x"BE60D6AE",
    x"BE60BE29",
    x"BE60A5A4",
    x"BE608D1E",
    x"BE607499",
    x"BE605C13",
    x"BE60438E",
    x"BE602B08",
    x"BE601282",
    x"BE5FF9FC",
    x"BE5FE175",
    x"BE5FC8EF",
    x"BE5FB068",
    x"BE5F97E2",
    x"BE5F7F5B",
    x"BE5F66D4",
    x"BE5F4E4D",
    x"BE5F35C6",
    x"BE5F1D3E",
    x"BE5F04B7",
    x"BE5EEC2F",
    x"BE5ED3A8",
    x"BE5EBB20",
    x"BE5EA298",
    x"BE5E8A10",
    x"BE5E7187",
    x"BE5E58FF",
    x"BE5E4076",
    x"BE5E27EE",
    x"BE5E0F65",
    x"BE5DF6DC",
    x"BE5DDE53",
    x"BE5DC5CA",
    x"BE5DAD40",
    x"BE5D94B7",
    x"BE5D7C2D",
    x"BE5D63A4",
    x"BE5D4B1A",
    x"BE5D3290",
    x"BE5D1A05",
    x"BE5D017B",
    x"BE5CE8F1",
    x"BE5CD066",
    x"BE5CB7DC",
    x"BE5C9F51",
    x"BE5C86C6",
    x"BE5C6E3B",
    x"BE5C55B0",
    x"BE5C3D24",
    x"BE5C2499",
    x"BE5C0C0D",
    x"BE5BF381",
    x"BE5BDAF6",
    x"BE5BC26A",
    x"BE5BA9DD",
    x"BE5B9151",
    x"BE5B78C5",
    x"BE5B6038",
    x"BE5B47AC",
    x"BE5B2F1F",
    x"BE5B1692",
    x"BE5AFE05",
    x"BE5AE578",
    x"BE5ACCEA",
    x"BE5AB45D",
    x"BE5A9BCF",
    x"BE5A8341",
    x"BE5A6AB4",
    x"BE5A5226",
    x"BE5A3997",
    x"BE5A2109",
    x"BE5A087B",
    x"BE59EFEC",
    x"BE59D75E",
    x"BE59BECF",
    x"BE59A640",
    x"BE598DB1",
    x"BE597522",
    x"BE595C93",
    x"BE594403",
    x"BE592B74",
    x"BE5912E4",
    x"BE58FA54",
    x"BE58E1C4",
    x"BE58C934",
    x"BE58B0A4",
    x"BE589813",
    x"BE587F83",
    x"BE5866F2",
    x"BE584E62",
    x"BE5835D1",
    x"BE581D40",
    x"BE5804AF",
    x"BE57EC1D",
    x"BE57D38C",
    x"BE57BAFB",
    x"BE57A269",
    x"BE5789D7",
    x"BE577145",
    x"BE5758B3",
    x"BE574021",
    x"BE57278F",
    x"BE570EFC",
    x"BE56F66A",
    x"BE56DDD7",
    x"BE56C544",
    x"BE56ACB1",
    x"BE56941E",
    x"BE567B8B",
    x"BE5662F8",
    x"BE564A64",
    x"BE5631D1",
    x"BE56193D",
    x"BE5600A9",
    x"BE55E815",
    x"BE55CF81",
    x"BE55B6ED",
    x"BE559E58",
    x"BE5585C4",
    x"BE556D2F",
    x"BE55549B",
    x"BE553C06",
    x"BE552371",
    x"BE550ADC",
    x"BE54F246",
    x"BE54D9B1",
    x"BE54C11B",
    x"BE54A886",
    x"BE548FF0",
    x"BE54775A",
    x"BE545EC4",
    x"BE54462E",
    x"BE542D98",
    x"BE541501",
    x"BE53FC6B",
    x"BE53E3D4",
    x"BE53CB3D",
    x"BE53B2A6",
    x"BE539A0F",
    x"BE538178",
    x"BE5368E1",
    x"BE535049",
    x"BE5337B2",
    x"BE531F1A",
    x"BE530682",
    x"BE52EDEA",
    x"BE52D552",
    x"BE52BCBA",
    x"BE52A422",
    x"BE528B89",
    x"BE5272F1",
    x"BE525A58",
    x"BE5241BF",
    x"BE522926",
    x"BE52108D",
    x"BE51F7F4",
    x"BE51DF5B",
    x"BE51C6C1",
    x"BE51AE28",
    x"BE51958E",
    x"BE517CF4",
    x"BE51645A",
    x"BE514BC0",
    x"BE513326",
    x"BE511A8B",
    x"BE5101F1",
    x"BE50E956",
    x"BE50D0BC",
    x"BE50B821",
    x"BE509F86",
    x"BE5086EB",
    x"BE506E4F",
    x"BE5055B4",
    x"BE503D19",
    x"BE50247D",
    x"BE500BE1",
    x"BE4FF345",
    x"BE4FDAA9",
    x"BE4FC20D",
    x"BE4FA971",
    x"BE4F90D5",
    x"BE4F7838",
    x"BE4F5F9C",
    x"BE4F46FF",
    x"BE4F2E62",
    x"BE4F15C5",
    x"BE4EFD28",
    x"BE4EE48B",
    x"BE4ECBED",
    x"BE4EB350",
    x"BE4E9AB2",
    x"BE4E8215",
    x"BE4E6977",
    x"BE4E50D9",
    x"BE4E383B",
    x"BE4E1F9C",
    x"BE4E06FE",
    x"BE4DEE60",
    x"BE4DD5C1",
    x"BE4DBD22",
    x"BE4DA483",
    x"BE4D8BE4",
    x"BE4D7345",
    x"BE4D5AA6",
    x"BE4D4207",
    x"BE4D2967",
    x"BE4D10C8",
    x"BE4CF828",
    x"BE4CDF88",
    x"BE4CC6E8",
    x"BE4CAE48",
    x"BE4C95A8",
    x"BE4C7D08",
    x"BE4C6467",
    x"BE4C4BC7",
    x"BE4C3326",
    x"BE4C1A85",
    x"BE4C01E4",
    x"BE4BE943",
    x"BE4BD0A2",
    x"BE4BB801",
    x"BE4B9F5F",
    x"BE4B86BE",
    x"BE4B6E1C",
    x"BE4B557A",
    x"BE4B3CD8",
    x"BE4B2436",
    x"BE4B0B94",
    x"BE4AF2F2",
    x"BE4ADA4F",
    x"BE4AC1AD",
    x"BE4AA90A",
    x"BE4A9067",
    x"BE4A77C4",
    x"BE4A5F21",
    x"BE4A467E",
    x"BE4A2DDB",
    x"BE4A1538",
    x"BE49FC94",
    x"BE49E3F0",
    x"BE49CB4D",
    x"BE49B2A9",
    x"BE499A05",
    x"BE498161",
    x"BE4968BC",
    x"BE495018",
    x"BE493774",
    x"BE491ECF",
    x"BE49062A",
    x"BE48ED85",
    x"BE48D4E0",
    x"BE48BC3B",
    x"BE48A396",
    x"BE488AF1",
    x"BE48724B",
    x"BE4859A6",
    x"BE484100",
    x"BE48285A",
    x"BE480FB4",
    x"BE47F70E",
    x"BE47DE68",
    x"BE47C5C2",
    x"BE47AD1B",
    x"BE479475",
    x"BE477BCE",
    x"BE476328",
    x"BE474A81",
    x"BE4731DA",
    x"BE471932",
    x"BE47008B",
    x"BE46E7E4",
    x"BE46CF3C",
    x"BE46B695",
    x"BE469DED",
    x"BE468545",
    x"BE466C9D",
    x"BE4653F5",
    x"BE463B4D",
    x"BE4622A5",
    x"BE4609FC",
    x"BE45F153",
    x"BE45D8AB",
    x"BE45C002",
    x"BE45A759",
    x"BE458EB0",
    x"BE457607",
    x"BE455D5E",
    x"BE4544B4",
    x"BE452C0B",
    x"BE451361",
    x"BE44FAB7",
    x"BE44E20D",
    x"BE44C963",
    x"BE44B0B9",
    x"BE44980F",
    x"BE447F65",
    x"BE4466BA",
    x"BE444E10",
    x"BE443565",
    x"BE441CBA",
    x"BE44040F",
    x"BE43EB64",
    x"BE43D2B9",
    x"BE43BA0E",
    x"BE43A162",
    x"BE4388B7",
    x"BE43700B",
    x"BE43575F",
    x"BE433EB3",
    x"BE432607",
    x"BE430D5B",
    x"BE42F4AF",
    x"BE42DC03",
    x"BE42C356",
    x"BE42AAAA",
    x"BE4291FD",
    x"BE427950",
    x"BE4260A3",
    x"BE4247F6",
    x"BE422F49",
    x"BE42169B",
    x"BE41FDEE",
    x"BE41E541",
    x"BE41CC93",
    x"BE41B3E5",
    x"BE419B37",
    x"BE418289",
    x"BE4169DB",
    x"BE41512D",
    x"BE41387F",
    x"BE411FD0",
    x"BE410722",
    x"BE40EE73",
    x"BE40D5C4",
    x"BE40BD15",
    x"BE40A466",
    x"BE408BB7",
    x"BE407308",
    x"BE405A58",
    x"BE4041A9",
    x"BE4028F9",
    x"BE401049",
    x"BE3FF79A",
    x"BE3FDEEA",
    x"BE3FC639",
    x"BE3FAD89",
    x"BE3F94D9",
    x"BE3F7C29",
    x"BE3F6378",
    x"BE3F4AC7",
    x"BE3F3217",
    x"BE3F1966",
    x"BE3F00B5",
    x"BE3EE804",
    x"BE3ECF52",
    x"BE3EB6A1",
    x"BE3E9DEF",
    x"BE3E853E",
    x"BE3E6C8C",
    x"BE3E53DA",
    x"BE3E3B28",
    x"BE3E2276",
    x"BE3E09C4",
    x"BE3DF112",
    x"BE3DD860",
    x"BE3DBFAD",
    x"BE3DA6FA",
    x"BE3D8E48",
    x"BE3D7595",
    x"BE3D5CE2",
    x"BE3D442F",
    x"BE3D2B7C",
    x"BE3D12C8",
    x"BE3CFA15",
    x"BE3CE161",
    x"BE3CC8AE",
    x"BE3CAFFA",
    x"BE3C9746",
    x"BE3C7E92",
    x"BE3C65DE",
    x"BE3C4D2A",
    x"BE3C3476",
    x"BE3C1BC1",
    x"BE3C030D",
    x"BE3BEA58",
    x"BE3BD1A3",
    x"BE3BB8EE",
    x"BE3BA039",
    x"BE3B8784",
    x"BE3B6ECF",
    x"BE3B561A",
    x"BE3B3D64",
    x"BE3B24AF",
    x"BE3B0BF9",
    x"BE3AF343",
    x"BE3ADA8D",
    x"BE3AC1D7",
    x"BE3AA921",
    x"BE3A906B",
    x"BE3A77B4",
    x"BE3A5EFE",
    x"BE3A4647",
    x"BE3A2D91",
    x"BE3A14DA",
    x"BE39FC23",
    x"BE39E36C",
    x"BE39CAB5",
    x"BE39B1FE",
    x"BE399946",
    x"BE39808F",
    x"BE3967D7",
    x"BE394F20",
    x"BE393668",
    x"BE391DB0",
    x"BE3904F8",
    x"BE38EC40",
    x"BE38D387",
    x"BE38BACF",
    x"BE38A217",
    x"BE38895E",
    x"BE3870A5",
    x"BE3857EC",
    x"BE383F33",
    x"BE38267A",
    x"BE380DC1",
    x"BE37F508",
    x"BE37DC4F",
    x"BE37C395",
    x"BE37AADC",
    x"BE379222",
    x"BE377968",
    x"BE3760AE",
    x"BE3747F4",
    x"BE372F3A",
    x"BE371680",
    x"BE36FDC5",
    x"BE36E50B",
    x"BE36CC50",
    x"BE36B396",
    x"BE369ADB",
    x"BE368220",
    x"BE366965",
    x"BE3650AA",
    x"BE3637EF",
    x"BE361F33",
    x"BE360678",
    x"BE35EDBC",
    x"BE35D501",
    x"BE35BC45",
    x"BE35A389",
    x"BE358ACD",
    x"BE357211",
    x"BE355954",
    x"BE354098",
    x"BE3527DC",
    x"BE350F1F",
    x"BE34F662",
    x"BE34DDA6",
    x"BE34C4E9",
    x"BE34AC2C",
    x"BE34936F",
    x"BE347AB2",
    x"BE3461F4",
    x"BE344937",
    x"BE343079",
    x"BE3417BC",
    x"BE33FEFE",
    x"BE33E640",
    x"BE33CD82",
    x"BE33B4C4",
    x"BE339C06",
    x"BE338348",
    x"BE336A89",
    x"BE3351CB",
    x"BE33390C",
    x"BE33204D",
    x"BE33078E",
    x"BE32EECF",
    x"BE32D610",
    x"BE32BD51",
    x"BE32A492",
    x"BE328BD3",
    x"BE327313",
    x"BE325A54",
    x"BE324194",
    x"BE3228D4",
    x"BE321014",
    x"BE31F754",
    x"BE31DE94",
    x"BE31C5D4",
    x"BE31AD13",
    x"BE319453",
    x"BE317B92",
    x"BE3162D2",
    x"BE314A11",
    x"BE313150",
    x"BE31188F",
    x"BE30FFCE",
    x"BE30E70D",
    x"BE30CE4C",
    x"BE30B58A",
    x"BE309CC9",
    x"BE308407",
    x"BE306B45",
    x"BE305284",
    x"BE3039C2",
    x"BE302100",
    x"BE30083D",
    x"BE2FEF7B",
    x"BE2FD6B9",
    x"BE2FBDF6",
    x"BE2FA534",
    x"BE2F8C71",
    x"BE2F73AE",
    x"BE2F5AEB",
    x"BE2F4228",
    x"BE2F2965",
    x"BE2F10A2",
    x"BE2EF7DF",
    x"BE2EDF1B",
    x"BE2EC658",
    x"BE2EAD94",
    x"BE2E94D1",
    x"BE2E7C0D",
    x"BE2E6349",
    x"BE2E4A85",
    x"BE2E31C1",
    x"BE2E18FC",
    x"BE2E0038",
    x"BE2DE773",
    x"BE2DCEAF",
    x"BE2DB5EA",
    x"BE2D9D25",
    x"BE2D8461",
    x"BE2D6B9C",
    x"BE2D52D6",
    x"BE2D3A11",
    x"BE2D214C",
    x"BE2D0887",
    x"BE2CEFC1",
    x"BE2CD6FB",
    x"BE2CBE36",
    x"BE2CA570",
    x"BE2C8CAA",
    x"BE2C73E4",
    x"BE2C5B1E",
    x"BE2C4258",
    x"BE2C2991",
    x"BE2C10CB",
    x"BE2BF804",
    x"BE2BDF3E",
    x"BE2BC677",
    x"BE2BADB0",
    x"BE2B94E9",
    x"BE2B7C22",
    x"BE2B635B",
    x"BE2B4A93",
    x"BE2B31CC",
    x"BE2B1905",
    x"BE2B003D",
    x"BE2AE775",
    x"BE2ACEAE",
    x"BE2AB5E6",
    x"BE2A9D1E",
    x"BE2A8456",
    x"BE2A6B8D",
    x"BE2A52C5",
    x"BE2A39FD",
    x"BE2A2134",
    x"BE2A086B",
    x"BE29EFA3",
    x"BE29D6DA",
    x"BE29BE11",
    x"BE29A548",
    x"BE298C7F",
    x"BE2973B6",
    x"BE295AEC",
    x"BE294223",
    x"BE292959",
    x"BE291090",
    x"BE28F7C6",
    x"BE28DEFC",
    x"BE28C632",
    x"BE28AD68",
    x"BE28949E",
    x"BE287BD4",
    x"BE286309",
    x"BE284A3F",
    x"BE283174",
    x"BE2818AA",
    x"BE27FFDF",
    x"BE27E714",
    x"BE27CE49",
    x"BE27B57E",
    x"BE279CB3",
    x"BE2783E8",
    x"BE276B1C",
    x"BE275251",
    x"BE273985",
    x"BE2720BA",
    x"BE2707EE",
    x"BE26EF22",
    x"BE26D656",
    x"BE26BD8A",
    x"BE26A4BE",
    x"BE268BF2",
    x"BE267325",
    x"BE265A59",
    x"BE26418C",
    x"BE2628C0",
    x"BE260FF3",
    x"BE25F726",
    x"BE25DE59",
    x"BE25C58C",
    x"BE25ACBF",
    x"BE2593F2",
    x"BE257B24",
    x"BE256257",
    x"BE254989",
    x"BE2530BC",
    x"BE2517EE",
    x"BE24FF20",
    x"BE24E652",
    x"BE24CD84",
    x"BE24B4B6",
    x"BE249BE7",
    x"BE248319",
    x"BE246A4B",
    x"BE24517C",
    x"BE2438AD",
    x"BE241FDF",
    x"BE240710",
    x"BE23EE41",
    x"BE23D572",
    x"BE23BCA3",
    x"BE23A3D3",
    x"BE238B04",
    x"BE237235",
    x"BE235965",
    x"BE234095",
    x"BE2327C6",
    x"BE230EF6",
    x"BE22F626",
    x"BE22DD56",
    x"BE22C486",
    x"BE22ABB6",
    x"BE2292E5",
    x"BE227A15",
    x"BE226144",
    x"BE224874",
    x"BE222FA3",
    x"BE2216D2",
    x"BE21FE01",
    x"BE21E530",
    x"BE21CC5F",
    x"BE21B38E",
    x"BE219ABD",
    x"BE2181EB",
    x"BE21691A",
    x"BE215048",
    x"BE213776",
    x"BE211EA5",
    x"BE2105D3",
    x"BE20ED01",
    x"BE20D42F",
    x"BE20BB5C",
    x"BE20A28A",
    x"BE2089B8",
    x"BE2070E5",
    x"BE205813",
    x"BE203F40",
    x"BE20266D",
    x"BE200D9A",
    x"BE1FF4C8",
    x"BE1FDBF4",
    x"BE1FC321",
    x"BE1FAA4E",
    x"BE1F917B",
    x"BE1F78A7",
    x"BE1F5FD4",
    x"BE1F4700",
    x"BE1F2E2C",
    x"BE1F1559",
    x"BE1EFC85",
    x"BE1EE3B1",
    x"BE1ECADD",
    x"BE1EB208",
    x"BE1E9934",
    x"BE1E8060",
    x"BE1E678B",
    x"BE1E4EB7",
    x"BE1E35E2",
    x"BE1E1D0D",
    x"BE1E0438",
    x"BE1DEB63",
    x"BE1DD28E",
    x"BE1DB9B9",
    x"BE1DA0E4",
    x"BE1D880F",
    x"BE1D6F39",
    x"BE1D5664",
    x"BE1D3D8E",
    x"BE1D24B8",
    x"BE1D0BE2",
    x"BE1CF30D",
    x"BE1CDA36",
    x"BE1CC160",
    x"BE1CA88A",
    x"BE1C8FB4",
    x"BE1C76DE",
    x"BE1C5E07",
    x"BE1C4530",
    x"BE1C2C5A",
    x"BE1C1383",
    x"BE1BFAAC",
    x"BE1BE1D5",
    x"BE1BC8FE",
    x"BE1BB027",
    x"BE1B9750",
    x"BE1B7E79",
    x"BE1B65A1",
    x"BE1B4CCA",
    x"BE1B33F2",
    x"BE1B1B1A",
    x"BE1B0242",
    x"BE1AE96B",
    x"BE1AD093",
    x"BE1AB7BB",
    x"BE1A9EE2",
    x"BE1A860A",
    x"BE1A6D32",
    x"BE1A5459",
    x"BE1A3B81",
    x"BE1A22A8",
    x"BE1A09CF",
    x"BE19F0F7",
    x"BE19D81E",
    x"BE19BF45",
    x"BE19A66C",
    x"BE198D92",
    x"BE1974B9",
    x"BE195BE0",
    x"BE194306",
    x"BE192A2D",
    x"BE191153",
    x"BE18F879",
    x"BE18DFA0",
    x"BE18C6C6",
    x"BE18ADEC",
    x"BE189511",
    x"BE187C37",
    x"BE18635D",
    x"BE184A83",
    x"BE1831A8",
    x"BE1818CE",
    x"BE17FFF3",
    x"BE17E718",
    x"BE17CE3D",
    x"BE17B562",
    x"BE179C87",
    x"BE1783AC",
    x"BE176AD1",
    x"BE1751F6",
    x"BE17391A",
    x"BE17203F",
    x"BE170763",
    x"BE16EE88",
    x"BE16D5AC",
    x"BE16BCD0",
    x"BE16A3F4",
    x"BE168B18",
    x"BE16723C",
    x"BE165960",
    x"BE164083",
    x"BE1627A7",
    x"BE160ECB",
    x"BE15F5EE",
    x"BE15DD11",
    x"BE15C435",
    x"BE15AB58",
    x"BE15927B",
    x"BE15799E",
    x"BE1560C1",
    x"BE1547E4",
    x"BE152F06",
    x"BE151629",
    x"BE14FD4B",
    x"BE14E46E",
    x"BE14CB90",
    x"BE14B2B2",
    x"BE1499D5",
    x"BE1480F7",
    x"BE146819",
    x"BE144F3B",
    x"BE14365C",
    x"BE141D7E",
    x"BE1404A0",
    x"BE13EBC1",
    x"BE13D2E3",
    x"BE13BA04",
    x"BE13A125",
    x"BE138847",
    x"BE136F68",
    x"BE135689",
    x"BE133DAA",
    x"BE1324CA",
    x"BE130BEB",
    x"BE12F30C",
    x"BE12DA2C",
    x"BE12C14D",
    x"BE12A86D",
    x"BE128F8E",
    x"BE1276AE",
    x"BE125DCE",
    x"BE1244EE",
    x"BE122C0E",
    x"BE12132E",
    x"BE11FA4E",
    x"BE11E16D",
    x"BE11C88D",
    x"BE11AFAC",
    x"BE1196CC",
    x"BE117DEB",
    x"BE11650A",
    x"BE114C2A",
    x"BE113349",
    x"BE111A68",
    x"BE110186",
    x"BE10E8A5",
    x"BE10CFC4",
    x"BE10B6E3",
    x"BE109E01",
    x"BE108520",
    x"BE106C3E",
    x"BE10535C",
    x"BE103A7B",
    x"BE102199",
    x"BE1008B7",
    x"BE0FEFD5",
    x"BE0FD6F2",
    x"BE0FBE10",
    x"BE0FA52E",
    x"BE0F8C4B",
    x"BE0F7369",
    x"BE0F5A86",
    x"BE0F41A4",
    x"BE0F28C1",
    x"BE0F0FDE",
    x"BE0EF6FB",
    x"BE0EDE18",
    x"BE0EC535",
    x"BE0EAC52",
    x"BE0E936F",
    x"BE0E7A8B",
    x"BE0E61A8",
    x"BE0E48C4",
    x"BE0E2FE1",
    x"BE0E16FD",
    x"BE0DFE19",
    x"BE0DE535",
    x"BE0DCC51",
    x"BE0DB36D",
    x"BE0D9A89",
    x"BE0D81A5",
    x"BE0D68C1",
    x"BE0D4FDC",
    x"BE0D36F8",
    x"BE0D1E13",
    x"BE0D052F",
    x"BE0CEC4A",
    x"BE0CD365",
    x"BE0CBA80",
    x"BE0CA19B",
    x"BE0C88B6",
    x"BE0C6FD1",
    x"BE0C56EC",
    x"BE0C3E07",
    x"BE0C2521",
    x"BE0C0C3C",
    x"BE0BF356",
    x"BE0BDA71",
    x"BE0BC18B",
    x"BE0BA8A5",
    x"BE0B8FBF",
    x"BE0B76D9",
    x"BE0B5DF3",
    x"BE0B450D",
    x"BE0B2C27",
    x"BE0B1340",
    x"BE0AFA5A",
    x"BE0AE173",
    x"BE0AC88D",
    x"BE0AAFA6",
    x"BE0A96BF",
    x"BE0A7DD9",
    x"BE0A64F2",
    x"BE0A4C0B",
    x"BE0A3324",
    x"BE0A1A3C",
    x"BE0A0155",
    x"BE09E86E",
    x"BE09CF86",
    x"BE09B69F",
    x"BE099DB7",
    x"BE0984D0",
    x"BE096BE8",
    x"BE095300",
    x"BE093A18",
    x"BE092130",
    x"BE090848",
    x"BE08EF60",
    x"BE08D678",
    x"BE08BD90",
    x"BE08A4A7",
    x"BE088BBF",
    x"BE0872D6",
    x"BE0859ED",
    x"BE084105",
    x"BE08281C",
    x"BE080F33",
    x"BE07F64A",
    x"BE07DD61",
    x"BE07C478",
    x"BE07AB8F",
    x"BE0792A5",
    x"BE0779BC",
    x"BE0760D2",
    x"BE0747E9",
    x"BE072EFF",
    x"BE071616",
    x"BE06FD2C",
    x"BE06E442",
    x"BE06CB58",
    x"BE06B26E",
    x"BE069984",
    x"BE06809A",
    x"BE0667AF",
    x"BE064EC5",
    x"BE0635DB",
    x"BE061CF0",
    x"BE060405",
    x"BE05EB1B",
    x"BE05D230",
    x"BE05B945",
    x"BE05A05A",
    x"BE05876F",
    x"BE056E84",
    x"BE055599",
    x"BE053CAE",
    x"BE0523C2",
    x"BE050AD7",
    x"BE04F1EB",
    x"BE04D900",
    x"BE04C014",
    x"BE04A729",
    x"BE048E3D",
    x"BE047551",
    x"BE045C65",
    x"BE044379",
    x"BE042A8D",
    x"BE0411A0",
    x"BE03F8B4",
    x"BE03DFC8",
    x"BE03C6DB",
    x"BE03ADEF",
    x"BE039502",
    x"BE037C16",
    x"BE036329",
    x"BE034A3C",
    x"BE03314F",
    x"BE031862",
    x"BE02FF75",
    x"BE02E688",
    x"BE02CD9B",
    x"BE02B4AD",
    x"BE029BC0",
    x"BE0282D2",
    x"BE0269E5",
    x"BE0250F7",
    x"BE02380A",
    x"BE021F1C",
    x"BE02062E",
    x"BE01ED40",
    x"BE01D452",
    x"BE01BB64",
    x"BE01A276",
    x"BE018987",
    x"BE017099",
    x"BE0157AB",
    x"BE013EBC",
    x"BE0125CE",
    x"BE010CDF",
    x"BE00F3F0",
    x"BE00DB01",
    x"BE00C213",
    x"BE00A924",
    x"BE009035",
    x"BE007745",
    x"BE005E56",
    x"BE004567",
    x"BE002C78",
    x"BE001388",
    x"BDFFF531",
    x"BDFFC352",
    x"BDFF9173",
    x"BDFF5F94",
    x"BDFF2DB4",
    x"BDFEFBD4",
    x"BDFEC9F4",
    x"BDFE9814",
    x"BDFE6634",
    x"BDFE3454",
    x"BDFE0273",
    x"BDFDD092",
    x"BDFD9EB2",
    x"BDFD6CD1",
    x"BDFD3AEF",
    x"BDFD090E",
    x"BDFCD72D",
    x"BDFCA54B",
    x"BDFC7369",
    x"BDFC4187",
    x"BDFC0FA5",
    x"BDFBDDC3",
    x"BDFBABE1",
    x"BDFB79FE",
    x"BDFB481C",
    x"BDFB1639",
    x"BDFAE456",
    x"BDFAB273",
    x"BDFA808F",
    x"BDFA4EAC",
    x"BDFA1CC8",
    x"BDF9EAE5",
    x"BDF9B901",
    x"BDF9871D",
    x"BDF95539",
    x"BDF92354",
    x"BDF8F170",
    x"BDF8BF8B",
    x"BDF88DA7",
    x"BDF85BC2",
    x"BDF829DD",
    x"BDF7F7F7",
    x"BDF7C612",
    x"BDF7942C",
    x"BDF76247",
    x"BDF73061",
    x"BDF6FE7B",
    x"BDF6CC95",
    x"BDF69AAF",
    x"BDF668C8",
    x"BDF636E2",
    x"BDF604FB",
    x"BDF5D314",
    x"BDF5A12D",
    x"BDF56F46",
    x"BDF53D5F",
    x"BDF50B77",
    x"BDF4D990",
    x"BDF4A7A8",
    x"BDF475C0",
    x"BDF443D8",
    x"BDF411F0",
    x"BDF3E007",
    x"BDF3AE1F",
    x"BDF37C36",
    x"BDF34A4E",
    x"BDF31865",
    x"BDF2E67C",
    x"BDF2B492",
    x"BDF282A9",
    x"BDF250BF",
    x"BDF21ED6",
    x"BDF1ECEC",
    x"BDF1BB02",
    x"BDF18918",
    x"BDF1572E",
    x"BDF12543",
    x"BDF0F359",
    x"BDF0C16E",
    x"BDF08F83",
    x"BDF05D98",
    x"BDF02BAD",
    x"BDEFF9C2",
    x"BDEFC7D7",
    x"BDEF95EB",
    x"BDEF63FF",
    x"BDEF3214",
    x"BDEF0028",
    x"BDEECE3C",
    x"BDEE9C4F",
    x"BDEE6A63",
    x"BDEE3876",
    x"BDEE068A",
    x"BDEDD49D",
    x"BDEDA2B0",
    x"BDED70C3",
    x"BDED3ED5",
    x"BDED0CE8",
    x"BDECDAFB",
    x"BDECA90D",
    x"BDEC771F",
    x"BDEC4531",
    x"BDEC1343",
    x"BDEBE155",
    x"BDEBAF66",
    x"BDEB7D78",
    x"BDEB4B89",
    x"BDEB199A",
    x"BDEAE7AB",
    x"BDEAB5BC",
    x"BDEA83CD",
    x"BDEA51DE",
    x"BDEA1FEE",
    x"BDE9EDFE",
    x"BDE9BC0E",
    x"BDE98A1F",
    x"BDE9582E",
    x"BDE9263E",
    x"BDE8F44E",
    x"BDE8C25D",
    x"BDE8906D",
    x"BDE85E7C",
    x"BDE82C8B",
    x"BDE7FA9A",
    x"BDE7C8A9",
    x"BDE796B7",
    x"BDE764C6",
    x"BDE732D4",
    x"BDE700E2",
    x"BDE6CEF0",
    x"BDE69CFE",
    x"BDE66B0C",
    x"BDE6391A",
    x"BDE60727",
    x"BDE5D535",
    x"BDE5A342",
    x"BDE5714F",
    x"BDE53F5C",
    x"BDE50D69",
    x"BDE4DB76",
    x"BDE4A982",
    x"BDE4778F",
    x"BDE4459B",
    x"BDE413A7",
    x"BDE3E1B3",
    x"BDE3AFBF",
    x"BDE37DCB",
    x"BDE34BD6",
    x"BDE319E2",
    x"BDE2E7ED",
    x"BDE2B5F8",
    x"BDE28403",
    x"BDE2520E",
    x"BDE22019",
    x"BDE1EE24",
    x"BDE1BC2E",
    x"BDE18A39",
    x"BDE15843",
    x"BDE1264D",
    x"BDE0F457",
    x"BDE0C261",
    x"BDE0906A",
    x"BDE05E74",
    x"BDE02C7D",
    x"BDDFFA87",
    x"BDDFC890",
    x"BDDF9699",
    x"BDDF64A2",
    x"BDDF32AB",
    x"BDDF00B3",
    x"BDDECEBC",
    x"BDDE9CC4",
    x"BDDE6ACC",
    x"BDDE38D4",
    x"BDDE06DC",
    x"BDDDD4E4",
    x"BDDDA2EC",
    x"BDDD70F3",
    x"BDDD3EFB",
    x"BDDD0D02",
    x"BDDCDB09",
    x"BDDCA910",
    x"BDDC7717",
    x"BDDC451E",
    x"BDDC1324",
    x"BDDBE12B",
    x"BDDBAF31",
    x"BDDB7D37",
    x"BDDB4B3D",
    x"BDDB1943",
    x"BDDAE749",
    x"BDDAB54F",
    x"BDDA8354",
    x"BDDA515A",
    x"BDDA1F5F",
    x"BDD9ED64",
    x"BDD9BB69",
    x"BDD9896E",
    x"BDD95773",
    x"BDD92578",
    x"BDD8F37C",
    x"BDD8C181",
    x"BDD88F85",
    x"BDD85D89",
    x"BDD82B8D",
    x"BDD7F991",
    x"BDD7C795",
    x"BDD79598",
    x"BDD7639C",
    x"BDD7319F",
    x"BDD6FFA2",
    x"BDD6CDA5",
    x"BDD69BA8",
    x"BDD669AB",
    x"BDD637AE",
    x"BDD605B0",
    x"BDD5D3B3",
    x"BDD5A1B5",
    x"BDD56FB7",
    x"BDD53DB9",
    x"BDD50BBB",
    x"BDD4D9BD",
    x"BDD4A7BE",
    x"BDD475C0",
    x"BDD443C1",
    x"BDD411C3",
    x"BDD3DFC4",
    x"BDD3ADC5",
    x"BDD37BC6",
    x"BDD349C7",
    x"BDD317C7",
    x"BDD2E5C8",
    x"BDD2B3C8",
    x"BDD281C8",
    x"BDD24FC8",
    x"BDD21DC8",
    x"BDD1EBC8",
    x"BDD1B9C8",
    x"BDD187C8",
    x"BDD155C7",
    x"BDD123C7",
    x"BDD0F1C6",
    x"BDD0BFC5",
    x"BDD08DC4",
    x"BDD05BC3",
    x"BDD029C2",
    x"BDCFF7C0",
    x"BDCFC5BF",
    x"BDCF93BD",
    x"BDCF61BB",
    x"BDCF2FB9",
    x"BDCEFDB7",
    x"BDCECBB5",
    x"BDCE99B3",
    x"BDCE67B1",
    x"BDCE35AE",
    x"BDCE03AB",
    x"BDCDD1A9",
    x"BDCD9FA6",
    x"BDCD6DA3",
    x"BDCD3BA0",
    x"BDCD099C",
    x"BDCCD799",
    x"BDCCA596",
    x"BDCC7392",
    x"BDCC418E",
    x"BDCC0F8A",
    x"BDCBDD86",
    x"BDCBAB82",
    x"BDCB797E",
    x"BDCB477A",
    x"BDCB1575",
    x"BDCAE371",
    x"BDCAB16C",
    x"BDCA7F67",
    x"BDCA4D62",
    x"BDCA1B5D",
    x"BDC9E958",
    x"BDC9B752",
    x"BDC9854D",
    x"BDC95347",
    x"BDC92142",
    x"BDC8EF3C",
    x"BDC8BD36",
    x"BDC88B30",
    x"BDC8592A",
    x"BDC82723",
    x"BDC7F51D",
    x"BDC7C316",
    x"BDC79110",
    x"BDC75F09",
    x"BDC72D02",
    x"BDC6FAFB",
    x"BDC6C8F4",
    x"BDC696ED",
    x"BDC664E5",
    x"BDC632DE",
    x"BDC600D6",
    x"BDC5CECE",
    x"BDC59CC6",
    x"BDC56ABE",
    x"BDC538B6",
    x"BDC506AE",
    x"BDC4D4A6",
    x"BDC4A29D",
    x"BDC47095",
    x"BDC43E8C",
    x"BDC40C83",
    x"BDC3DA7A",
    x"BDC3A871",
    x"BDC37668",
    x"BDC3445F",
    x"BDC31255",
    x"BDC2E04C",
    x"BDC2AE42",
    x"BDC27C39",
    x"BDC24A2F",
    x"BDC21825",
    x"BDC1E61B",
    x"BDC1B410",
    x"BDC18206",
    x"BDC14FFC",
    x"BDC11DF1",
    x"BDC0EBE6",
    x"BDC0B9DC",
    x"BDC087D1",
    x"BDC055C6",
    x"BDC023BA",
    x"BDBFF1AF",
    x"BDBFBFA4",
    x"BDBF8D98",
    x"BDBF5B8D",
    x"BDBF2981",
    x"BDBEF775",
    x"BDBEC569",
    x"BDBE935D",
    x"BDBE6151",
    x"BDBE2F45",
    x"BDBDFD38",
    x"BDBDCB2C",
    x"BDBD991F",
    x"BDBD6712",
    x"BDBD3505",
    x"BDBD02F8",
    x"BDBCD0EB",
    x"BDBC9EDE",
    x"BDBC6CD1",
    x"BDBC3AC3",
    x"BDBC08B6",
    x"BDBBD6A8",
    x"BDBBA49A",
    x"BDBB728C",
    x"BDBB407E",
    x"BDBB0E70",
    x"BDBADC62",
    x"BDBAAA54",
    x"BDBA7845",
    x"BDBA4637",
    x"BDBA1428",
    x"BDB9E219",
    x"BDB9B00A",
    x"BDB97DFB",
    x"BDB94BEC",
    x"BDB919DD",
    x"BDB8E7CE",
    x"BDB8B5BE",
    x"BDB883AF",
    x"BDB8519F",
    x"BDB81F8F",
    x"BDB7ED7F",
    x"BDB7BB6F",
    x"BDB7895F",
    x"BDB7574F",
    x"BDB7253E",
    x"BDB6F32E",
    x"BDB6C11D",
    x"BDB68F0D",
    x"BDB65CFC",
    x"BDB62AEB",
    x"BDB5F8DA",
    x"BDB5C6C9",
    x"BDB594B8",
    x"BDB562A6",
    x"BDB53095",
    x"BDB4FE83",
    x"BDB4CC72",
    x"BDB49A60",
    x"BDB4684E",
    x"BDB4363C",
    x"BDB4042A",
    x"BDB3D218",
    x"BDB3A005",
    x"BDB36DF3",
    x"BDB33BE0",
    x"BDB309CE",
    x"BDB2D7BB",
    x"BDB2A5A8",
    x"BDB27395",
    x"BDB24182",
    x"BDB20F6F",
    x"BDB1DD5C",
    x"BDB1AB48",
    x"BDB17935",
    x"BDB14721",
    x"BDB1150D",
    x"BDB0E2FA",
    x"BDB0B0E6",
    x"BDB07ED2",
    x"BDB04CBD",
    x"BDB01AA9",
    x"BDAFE895",
    x"BDAFB680",
    x"BDAF846C",
    x"BDAF5257",
    x"BDAF2042",
    x"BDAEEE2D",
    x"BDAEBC18",
    x"BDAE8A03",
    x"BDAE57EE",
    x"BDAE25D9",
    x"BDADF3C3",
    x"BDADC1AE",
    x"BDAD8F98",
    x"BDAD5D83",
    x"BDAD2B6D",
    x"BDACF957",
    x"BDACC741",
    x"BDAC952B",
    x"BDAC6314",
    x"BDAC30FE",
    x"BDABFEE8",
    x"BDABCCD1",
    x"BDAB9ABA",
    x"BDAB68A4",
    x"BDAB368D",
    x"BDAB0476",
    x"BDAAD25F",
    x"BDAAA048",
    x"BDAA6E30",
    x"BDAA3C19",
    x"BDAA0A01",
    x"BDA9D7EA",
    x"BDA9A5D2",
    x"BDA973BA",
    x"BDA941A2",
    x"BDA90F8A",
    x"BDA8DD72",
    x"BDA8AB5A",
    x"BDA87942",
    x"BDA84729",
    x"BDA81511",
    x"BDA7E2F8",
    x"BDA7B0E0",
    x"BDA77EC7",
    x"BDA74CAE",
    x"BDA71A95",
    x"BDA6E87C",
    x"BDA6B663",
    x"BDA68449",
    x"BDA65230",
    x"BDA62016",
    x"BDA5EDFD",
    x"BDA5BBE3",
    x"BDA589C9",
    x"BDA557AF",
    x"BDA52595",
    x"BDA4F37B",
    x"BDA4C161",
    x"BDA48F47",
    x"BDA45D2C",
    x"BDA42B12",
    x"BDA3F8F7",
    x"BDA3C6DC",
    x"BDA394C2",
    x"BDA362A7",
    x"BDA3308C",
    x"BDA2FE71",
    x"BDA2CC55",
    x"BDA29A3A",
    x"BDA2681F",
    x"BDA23603",
    x"BDA203E8",
    x"BDA1D1CC",
    x"BDA19FB0",
    x"BDA16D94",
    x"BDA13B78",
    x"BDA1095C",
    x"BDA0D740",
    x"BDA0A524",
    x"BDA07308",
    x"BDA040EB",
    x"BDA00ECF",
    x"BD9FDCB2",
    x"BD9FAA95",
    x"BD9F7878",
    x"BD9F465B",
    x"BD9F143E",
    x"BD9EE221",
    x"BD9EB004",
    x"BD9E7DE7",
    x"BD9E4BC9",
    x"BD9E19AC",
    x"BD9DE78E",
    x"BD9DB570",
    x"BD9D8353",
    x"BD9D5135",
    x"BD9D1F17",
    x"BD9CECF9",
    x"BD9CBADA",
    x"BD9C88BC",
    x"BD9C569E",
    x"BD9C247F",
    x"BD9BF261",
    x"BD9BC042",
    x"BD9B8E23",
    x"BD9B5C05",
    x"BD9B29E6",
    x"BD9AF7C7",
    x"BD9AC5A7",
    x"BD9A9388",
    x"BD9A6169",
    x"BD9A2F4A",
    x"BD99FD2A",
    x"BD99CB0A",
    x"BD9998EB",
    x"BD9966CB",
    x"BD9934AB",
    x"BD99028B",
    x"BD98D06B",
    x"BD989E4B",
    x"BD986C2B",
    x"BD983A0A",
    x"BD9807EA",
    x"BD97D5CA",
    x"BD97A3A9",
    x"BD977188",
    x"BD973F67",
    x"BD970D47",
    x"BD96DB26",
    x"BD96A905",
    x"BD9676E3",
    x"BD9644C2",
    x"BD9612A1",
    x"BD95E07F",
    x"BD95AE5E",
    x"BD957C3C",
    x"BD954A1B",
    x"BD9517F9",
    x"BD94E5D7",
    x"BD94B3B5",
    x"BD948193",
    x"BD944F71",
    x"BD941D4F",
    x"BD93EB2C",
    x"BD93B90A",
    x"BD9386E7",
    x"BD9354C5",
    x"BD9322A2",
    x"BD92F07F",
    x"BD92BE5D",
    x"BD928C3A",
    x"BD925A17",
    x"BD9227F4",
    x"BD91F5D0",
    x"BD91C3AD",
    x"BD91918A",
    x"BD915F66",
    x"BD912D43",
    x"BD90FB1F",
    x"BD90C8FB",
    x"BD9096D8",
    x"BD9064B4",
    x"BD903290",
    x"BD90006C",
    x"BD8FCE47",
    x"BD8F9C23",
    x"BD8F69FF",
    x"BD8F37DA",
    x"BD8F05B6",
    x"BD8ED391",
    x"BD8EA16D",
    x"BD8E6F48",
    x"BD8E3D23",
    x"BD8E0AFE",
    x"BD8DD8D9",
    x"BD8DA6B4",
    x"BD8D748F",
    x"BD8D426A",
    x"BD8D1044",
    x"BD8CDE1F",
    x"BD8CABF9",
    x"BD8C79D4",
    x"BD8C47AE",
    x"BD8C1588",
    x"BD8BE362",
    x"BD8BB13C",
    x"BD8B7F16",
    x"BD8B4CF0",
    x"BD8B1ACA",
    x"BD8AE8A4",
    x"BD8AB67D",
    x"BD8A8457",
    x"BD8A5230",
    x"BD8A200A",
    x"BD89EDE3",
    x"BD89BBBC",
    x"BD898995",
    x"BD89576E",
    x"BD892547",
    x"BD88F320",
    x"BD88C0F9",
    x"BD888ED2",
    x"BD885CAA",
    x"BD882A83",
    x"BD87F85B",
    x"BD87C634",
    x"BD87940C",
    x"BD8761E4",
    x"BD872FBC",
    x"BD86FD94",
    x"BD86CB6C",
    x"BD869944",
    x"BD86671C",
    x"BD8634F4",
    x"BD8602CC",
    x"BD85D0A3",
    x"BD859E7B",
    x"BD856C52",
    x"BD853A29",
    x"BD850801",
    x"BD84D5D8",
    x"BD84A3AF",
    x"BD847186",
    x"BD843F5D",
    x"BD840D34",
    x"BD83DB0A",
    x"BD83A8E1",
    x"BD8376B8",
    x"BD83448E",
    x"BD831265",
    x"BD82E03B",
    x"BD82AE11",
    x"BD827BE8",
    x"BD8249BE",
    x"BD821794",
    x"BD81E56A",
    x"BD81B340",
    x"BD818116",
    x"BD814EEB",
    x"BD811CC1",
    x"BD80EA97",
    x"BD80B86C",
    x"BD808642",
    x"BD805417",
    x"BD8021EC",
    x"BD7FDF83",
    x"BD7F7B2D",
    x"BD7F16D7",
    x"BD7EB281",
    x"BD7E4E2B",
    x"BD7DE9D5",
    x"BD7D857E",
    x"BD7D2127",
    x"BD7CBCD1",
    x"BD7C587A",
    x"BD7BF422",
    x"BD7B8FCB",
    x"BD7B2B74",
    x"BD7AC71C",
    x"BD7A62C5",
    x"BD79FE6D",
    x"BD799A15",
    x"BD7935BC",
    x"BD78D164",
    x"BD786D0C",
    x"BD7808B3",
    x"BD77A45A",
    x"BD774001",
    x"BD76DBA8",
    x"BD76774F",
    x"BD7612F6",
    x"BD75AE9C",
    x"BD754A42",
    x"BD74E5E9",
    x"BD74818F",
    x"BD741D35",
    x"BD73B8DA",
    x"BD735480",
    x"BD72F025",
    x"BD728BCB",
    x"BD722770",
    x"BD71C315",
    x"BD715EBA",
    x"BD70FA5E",
    x"BD709603",
    x"BD7031A8",
    x"BD6FCD4C",
    x"BD6F68F0",
    x"BD6F0494",
    x"BD6EA038",
    x"BD6E3BDC",
    x"BD6DD77F",
    x"BD6D7323",
    x"BD6D0EC6",
    x"BD6CAA69",
    x"BD6C460C",
    x"BD6BE1AF",
    x"BD6B7D51",
    x"BD6B18F4",
    x"BD6AB496",
    x"BD6A5039",
    x"BD69EBDB",
    x"BD69877D",
    x"BD69231F",
    x"BD68BEC1",
    x"BD685A62",
    x"BD67F604",
    x"BD6791A5",
    x"BD672D46",
    x"BD66C8E7",
    x"BD666488",
    x"BD660029",
    x"BD659BC9",
    x"BD65376A",
    x"BD64D30A",
    x"BD646EAA",
    x"BD640A4A",
    x"BD63A5EA",
    x"BD63418A",
    x"BD62DD2A",
    x"BD6278C9",
    x"BD621469",
    x"BD61B008",
    x"BD614BA7",
    x"BD60E746",
    x"BD6082E5",
    x"BD601E83",
    x"BD5FBA22",
    x"BD5F55C0",
    x"BD5EF15F",
    x"BD5E8CFD",
    x"BD5E289B",
    x"BD5DC439",
    x"BD5D5FD7",
    x"BD5CFB74",
    x"BD5C9712",
    x"BD5C32AF",
    x"BD5BCE4C",
    x"BD5B69E9",
    x"BD5B0586",
    x"BD5AA123",
    x"BD5A3CC0",
    x"BD59D85C",
    x"BD5973F9",
    x"BD590F95",
    x"BD58AB31",
    x"BD5846CD",
    x"BD57E269",
    x"BD577E05",
    x"BD5719A1",
    x"BD56B53C",
    x"BD5650D8",
    x"BD55EC73",
    x"BD55880E",
    x"BD5523A9",
    x"BD54BF44",
    x"BD545ADF",
    x"BD53F679",
    x"BD539214",
    x"BD532DAE",
    x"BD52C948",
    x"BD5264E2",
    x"BD52007C",
    x"BD519C16",
    x"BD5137B0",
    x"BD50D34A",
    x"BD506EE3",
    x"BD500A7C",
    x"BD4FA616",
    x"BD4F41AF",
    x"BD4EDD48",
    x"BD4E78E1",
    x"BD4E1479",
    x"BD4DB012",
    x"BD4D4BAA",
    x"BD4CE743",
    x"BD4C82DB",
    x"BD4C1E73",
    x"BD4BBA0B",
    x"BD4B55A3",
    x"BD4AF13B",
    x"BD4A8CD2",
    x"BD4A286A",
    x"BD49C401",
    x"BD495F98",
    x"BD48FB30",
    x"BD4896C7",
    x"BD48325D",
    x"BD47CDF4",
    x"BD47698B",
    x"BD470521",
    x"BD46A0B8",
    x"BD463C4E",
    x"BD45D7E4",
    x"BD45737A",
    x"BD450F10",
    x"BD44AAA6",
    x"BD44463C",
    x"BD43E1D1",
    x"BD437D67",
    x"BD4318FC",
    x"BD42B491",
    x"BD425026",
    x"BD41EBBB",
    x"BD418750",
    x"BD4122E5",
    x"BD40BE7A",
    x"BD405A0E",
    x"BD3FF5A3",
    x"BD3F9137",
    x"BD3F2CCB",
    x"BD3EC85F",
    x"BD3E63F3",
    x"BD3DFF87",
    x"BD3D9B1B",
    x"BD3D36AE",
    x"BD3CD242",
    x"BD3C6DD5",
    x"BD3C0968",
    x"BD3BA4FC",
    x"BD3B408F",
    x"BD3ADC22",
    x"BD3A77B4",
    x"BD3A1347",
    x"BD39AEDA",
    x"BD394A6C",
    x"BD38E5FE",
    x"BD388191",
    x"BD381D23",
    x"BD37B8B5",
    x"BD375447",
    x"BD36EFD9",
    x"BD368B6A",
    x"BD3626FC",
    x"BD35C28D",
    x"BD355E1F",
    x"BD34F9B0",
    x"BD349541",
    x"BD3430D2",
    x"BD33CC63",
    x"BD3367F4",
    x"BD330385",
    x"BD329F15",
    x"BD323AA6",
    x"BD31D636",
    x"BD3171C6",
    x"BD310D57",
    x"BD30A8E7",
    x"BD304477",
    x"BD2FE007",
    x"BD2F7B96",
    x"BD2F1726",
    x"BD2EB2B6",
    x"BD2E4E45",
    x"BD2DE9D4",
    x"BD2D8564",
    x"BD2D20F3",
    x"BD2CBC82",
    x"BD2C5811",
    x"BD2BF39F",
    x"BD2B8F2E",
    x"BD2B2ABD",
    x"BD2AC64B",
    x"BD2A61DA",
    x"BD29FD68",
    x"BD2998F6",
    x"BD293484",
    x"BD28D012",
    x"BD286BA0",
    x"BD28072E",
    x"BD27A2BC",
    x"BD273E49",
    x"BD26D9D7",
    x"BD267564",
    x"BD2610F1",
    x"BD25AC7E",
    x"BD25480C",
    x"BD24E399",
    x"BD247F25",
    x"BD241AB2",
    x"BD23B63F",
    x"BD2351CB",
    x"BD22ED58",
    x"BD2288E4",
    x"BD222471",
    x"BD21BFFD",
    x"BD215B89",
    x"BD20F715",
    x"BD2092A1",
    x"BD202E2D",
    x"BD1FC9B8",
    x"BD1F6544",
    x"BD1F00D0",
    x"BD1E9C5B",
    x"BD1E37E6",
    x"BD1DD372",
    x"BD1D6EFD",
    x"BD1D0A88",
    x"BD1CA613",
    x"BD1C419D",
    x"BD1BDD28",
    x"BD1B78B3",
    x"BD1B143D",
    x"BD1AAFC8",
    x"BD1A4B52",
    x"BD19E6DD",
    x"BD198267",
    x"BD191DF1",
    x"BD18B97B",
    x"BD185505",
    x"BD17F08F",
    x"BD178C18",
    x"BD1727A2",
    x"BD16C32C",
    x"BD165EB5",
    x"BD15FA3F",
    x"BD1595C8",
    x"BD153151",
    x"BD14CCDA",
    x"BD146863",
    x"BD1403EC",
    x"BD139F75",
    x"BD133AFE",
    x"BD12D686",
    x"BD12720F",
    x"BD120D97",
    x"BD11A920",
    x"BD1144A8",
    x"BD10E030",
    x"BD107BB8",
    x"BD101740",
    x"BD0FB2C8",
    x"BD0F4E50",
    x"BD0EE9D8",
    x"BD0E8560",
    x"BD0E20E7",
    x"BD0DBC6F",
    x"BD0D57F6",
    x"BD0CF37E",
    x"BD0C8F05",
    x"BD0C2A8C",
    x"BD0BC613",
    x"BD0B619A",
    x"BD0AFD21",
    x"BD0A98A8",
    x"BD0A342F",
    x"BD09CFB6",
    x"BD096B3C",
    x"BD0906C3",
    x"BD08A249",
    x"BD083DCF",
    x"BD07D956",
    x"BD0774DC",
    x"BD071062",
    x"BD06ABE8",
    x"BD06476E",
    x"BD05E2F4",
    x"BD057E7A",
    x"BD0519FF",
    x"BD04B585",
    x"BD04510B",
    x"BD03EC90",
    x"BD038815",
    x"BD03239B",
    x"BD02BF20",
    x"BD025AA5",
    x"BD01F62A",
    x"BD0191AF",
    x"BD012D34",
    x"BD00C8B9",
    x"BD00643E",
    x"BCFFFF85",
    x"BCFF368E",
    x"BCFE6D97",
    x"BCFDA4A0",
    x"BCFCDBA9",
    x"BCFC12B1",
    x"BCFB49BA",
    x"BCFA80C2",
    x"BCF9B7CA",
    x"BCF8EED2",
    x"BCF825DA",
    x"BCF75CE2",
    x"BCF693E9",
    x"BCF5CAF0",
    x"BCF501F8",
    x"BCF438FF",
    x"BCF37006",
    x"BCF2A70D",
    x"BCF1DE13",
    x"BCF1151A",
    x"BCF04C20",
    x"BCEF8326",
    x"BCEEBA2C",
    x"BCEDF132",
    x"BCED2838",
    x"BCEC5F3E",
    x"BCEB9643",
    x"BCEACD49",
    x"BCEA044E",
    x"BCE93B53",
    x"BCE87258",
    x"BCE7A95D",
    x"BCE6E061",
    x"BCE61766",
    x"BCE54E6A",
    x"BCE4856E",
    x"BCE3BC73",
    x"BCE2F377",
    x"BCE22A7A",
    x"BCE1617E",
    x"BCE09882",
    x"BCDFCF85",
    x"BCDF0688",
    x"BCDE3D8C",
    x"BCDD748F",
    x"BCDCAB91",
    x"BCDBE294",
    x"BCDB1997",
    x"BCDA5099",
    x"BCD9879C",
    x"BCD8BE9E",
    x"BCD7F5A0",
    x"BCD72CA2",
    x"BCD663A4",
    x"BCD59AA6",
    x"BCD4D1A7",
    x"BCD408A9",
    x"BCD33FAA",
    x"BCD276AB",
    x"BCD1ADAC",
    x"BCD0E4AD",
    x"BCD01BAE",
    x"BCCF52AF",
    x"BCCE89AF",
    x"BCCDC0B0",
    x"BCCCF7B0",
    x"BCCC2EB0",
    x"BCCB65B0",
    x"BCCA9CB0",
    x"BCC9D3B0",
    x"BCC90AB0",
    x"BCC841AF",
    x"BCC778AF",
    x"BCC6AFAE",
    x"BCC5E6AD",
    x"BCC51DAC",
    x"BCC454AB",
    x"BCC38BAA",
    x"BCC2C2A9",
    x"BCC1F9A8",
    x"BCC130A6",
    x"BCC067A5",
    x"BCBF9EA3",
    x"BCBED5A1",
    x"BCBE0C9F",
    x"BCBD439D",
    x"BCBC7A9B",
    x"BCBBB199",
    x"BCBAE896",
    x"BCBA1F94",
    x"BCB95691",
    x"BCB88D8E",
    x"BCB7C48C",
    x"BCB6FB89",
    x"BCB63286",
    x"BCB56982",
    x"BCB4A07F",
    x"BCB3D77C",
    x"BCB30E78",
    x"BCB24575",
    x"BCB17C71",
    x"BCB0B36D",
    x"BCAFEA69",
    x"BCAF2165",
    x"BCAE5861",
    x"BCAD8F5D",
    x"BCACC658",
    x"BCABFD54",
    x"BCAB344F",
    x"BCAA6B4B",
    x"BCA9A246",
    x"BCA8D941",
    x"BCA8103C",
    x"BCA74737",
    x"BCA67E32",
    x"BCA5B52C",
    x"BCA4EC27",
    x"BCA42322",
    x"BCA35A1C",
    x"BCA29116",
    x"BCA1C811",
    x"BCA0FF0B",
    x"BCA03605",
    x"BC9F6CFF",
    x"BC9EA3F9",
    x"BC9DDAF2",
    x"BC9D11EC",
    x"BC9C48E6",
    x"BC9B7FDF",
    x"BC9AB6D8",
    x"BC99EDD2",
    x"BC9924CB",
    x"BC985BC4",
    x"BC9792BD",
    x"BC96C9B6",
    x"BC9600AF",
    x"BC9537A7",
    x"BC946EA0",
    x"BC93A599",
    x"BC92DC91",
    x"BC921389",
    x"BC914A82",
    x"BC90817A",
    x"BC8FB872",
    x"BC8EEF6A",
    x"BC8E2662",
    x"BC8D5D5A",
    x"BC8C9452",
    x"BC8BCB49",
    x"BC8B0241",
    x"BC8A3938",
    x"BC897030",
    x"BC88A727",
    x"BC87DE1E",
    x"BC871516",
    x"BC864C0D",
    x"BC858304",
    x"BC84B9FB",
    x"BC83F0F2",
    x"BC8327E8",
    x"BC825EDF",
    x"BC8195D6",
    x"BC80CCCC",
    x"BC8003C3",
    x"BC7E7572",
    x"BC7CE35F",
    x"BC7B514B",
    x"BC79BF38",
    x"BC782D24",
    x"BC769B10",
    x"BC7508FC",
    x"BC7376E7",
    x"BC71E4D3",
    x"BC7052BF",
    x"BC6EC0AA",
    x"BC6D2E95",
    x"BC6B9C80",
    x"BC6A0A6B",
    x"BC687856",
    x"BC66E640",
    x"BC65542B",
    x"BC63C215",
    x"BC622FFF",
    x"BC609DE9",
    x"BC5F0BD3",
    x"BC5D79BD",
    x"BC5BE7A6",
    x"BC5A5590",
    x"BC58C379",
    x"BC573162",
    x"BC559F4C",
    x"BC540D35",
    x"BC527B1D",
    x"BC50E906",
    x"BC4F56EF",
    x"BC4DC4D7",
    x"BC4C32C0",
    x"BC4AA0A8",
    x"BC490E90",
    x"BC477C78",
    x"BC45EA60",
    x"BC445847",
    x"BC42C62F",
    x"BC413417",
    x"BC3FA1FE",
    x"BC3E0FE5",
    x"BC3C7DCC",
    x"BC3AEBB4",
    x"BC39599A",
    x"BC37C781",
    x"BC363568",
    x"BC34A34F",
    x"BC331135",
    x"BC317F1B",
    x"BC2FED02",
    x"BC2E5AE8",
    x"BC2CC8CE",
    x"BC2B36B4",
    x"BC29A49A",
    x"BC281280",
    x"BC268065",
    x"BC24EE4B",
    x"BC235C30",
    x"BC21CA16",
    x"BC2037FB",
    x"BC1EA5E0",
    x"BC1D13C5",
    x"BC1B81AA",
    x"BC19EF8F",
    x"BC185D74",
    x"BC16CB58",
    x"BC15393D",
    x"BC13A722",
    x"BC121506",
    x"BC1082EA",
    x"BC0EF0CF",
    x"BC0D5EB3",
    x"BC0BCC97",
    x"BC0A3A7B",
    x"BC08A85F",
    x"BC071643",
    x"BC058426",
    x"BC03F20A",
    x"BC025FEE",
    x"BC00CDD1",
    x"BBFE7769",
    x"BBFB5330",
    x"BBF82EF6",
    x"BBF50ABD",
    x"BBF1E683",
    x"BBEEC249",
    x"BBEB9E0F",
    x"BBE879D5",
    x"BBE5559B",
    x"BBE23160",
    x"BBDF0D26",
    x"BBDBE8EB",
    x"BBD8C4B0",
    x"BBD5A075",
    x"BBD27C3A",
    x"BBCF57FF",
    x"BBCC33C3",
    x"BBC90F88",
    x"BBC5EB4C",
    x"BBC2C711",
    x"BBBFA2D5",
    x"BBBC7E99",
    x"BBB95A5D",
    x"BBB63621",
    x"BBB311E4",
    x"BBAFEDA8",
    x"BBACC96B",
    x"BBA9A52F",
    x"BBA680F2",
    x"BBA35CB5",
    x"BBA03878",
    x"BB9D143B",
    x"BB99EFFE",
    x"BB96CBC1",
    x"BB93A784",
    x"BB908346",
    x"BB8D5F09",
    x"BB8A3ACB",
    x"BB87168E",
    x"BB83F250",
    x"BB80CE12",
    x"BB7B53A9",
    x"BB750B2D",
    x"BB6EC2B1",
    x"BB687A35",
    x"BB6231B9",
    x"BB5BE93C",
    x"BB55A0C0",
    x"BB4F5843",
    x"BB490FC6",
    x"BB42C749",
    x"BB3C7ECC",
    x"BB36364F",
    x"BB2FEDD1",
    x"BB29A554",
    x"BB235CD7",
    x"BB1D1459",
    x"BB16CBDB",
    x"BB10835D",
    x"BB0A3AE0",
    x"BB03F262",
    x"BAFB53C7",
    x"BAEEC2CB",
    x"BAE231CF",
    x"BAD5A0D2",
    x"BAC90FD5",
    x"BABC7ED9",
    x"BAAFEDDC",
    x"BAA35CDF",
    x"BA96CBE2",
    x"BA8A3AE5",
    x"BA7B53CF",
    x"BA6231D4",
    x"BA490FD9",
    x"BA2FEDDE",
    x"BA16CBE3",
    x"B9FB53D1",
    x"B9C90FDA",
    x"B996CBE4",
    x"B9490FDB",
    x"B8C90FDB"
  );

begin

  p_mem_read : process (clk) begin
    if rising_edge(clk) then
      data_out <= mem(to_integer(unsigned(address)));
    end if;
  end process;

end architecture;
