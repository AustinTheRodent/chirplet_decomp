
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity exponential_rom is
  port
  (
    clk       : in  std_logic;
    address   : in  std_logic_vector(15 downto 0);
    data_out  : out std_logic_vector(31 downto 0)
  );
end entity;

architecture rtl of exponential_rom is

  constant C_DATA_WIDTH  : integer := 32;
  constant C_ADDR_WIDTH  : integer := 16;

  constant RAM_DEPTH :integer := 2**C_ADDR_WIDTH;

  type RAM is array (integer range <>) of std_logic_vector (C_DATA_WIDTH-1 downto 0);
  signal mem : RAM (0 to RAM_DEPTH-1) :=
  (
    x"3F80000",
    x"3F7FC00",
    x"3F7F802",
    x"3F7F404",
    x"3F7F008",
    x"3F7EC0C",
    x"3F7E811",
    x"3F7E418",
    x"3F7E01F",
    x"3F7DC28",
    x"3F7D831",
    x"3F7D43C",
    x"3F7D047",
    x"3F7CC54",
    x"3F7C861",
    x"3F7C46F",
    x"3F7C07F",
    x"3F7BC8F",
    x"3F7B8A1",
    x"3F7B4B3",
    x"3F7B0C6",
    x"3F7ACDB",
    x"3F7A8F0",
    x"3F7A506",
    x"3F7A11D",
    x"3F79D36",
    x"3F7994F",
    x"3F79569",
    x"3F79184",
    x"3F78DA0",
    x"3F789BD",
    x"3F785DB",
    x"3F781FA",
    x"3F77E1A",
    x"3F77A3B",
    x"3F7765D",
    x"3F77280",
    x"3F76EA4",
    x"3F76AC9",
    x"3F766EE",
    x"3F76315",
    x"3F75F3D",
    x"3F75B66",
    x"3F7578F",
    x"3F753BA",
    x"3F74FE5",
    x"3F74C12",
    x"3F7483F",
    x"3F7446E",
    x"3F7409D",
    x"3F73CCD",
    x"3F738FF",
    x"3F73531",
    x"3F73164",
    x"3F72D98",
    x"3F729CD",
    x"3F72603",
    x"3F7223A",
    x"3F71E72",
    x"3F71AAB",
    x"3F716E5",
    x"3F71320",
    x"3F70F5B",
    x"3F70B98",
    x"3F707D6",
    x"3F70414",
    x"3F70053",
    x"3F6FC94",
    x"3F6F8D5",
    x"3F6F517",
    x"3F6F15B",
    x"3F6ED9F",
    x"3F6E9E4",
    x"3F6E62A",
    x"3F6E271",
    x"3F6DEB9",
    x"3F6DB01",
    x"3F6D74B",
    x"3F6D396",
    x"3F6CFE1",
    x"3F6CC2E",
    x"3F6C87B",
    x"3F6C4CA",
    x"3F6C119",
    x"3F6BD69",
    x"3F6B9BA",
    x"3F6B60C",
    x"3F6B25F",
    x"3F6AEB3",
    x"3F6AB08",
    x"3F6A75D",
    x"3F6A3B4",
    x"3F6A00C",
    x"3F69C64",
    x"3F698BD",
    x"3F69518",
    x"3F69173",
    x"3F68DCF",
    x"3F68A2C",
    x"3F6868A",
    x"3F682E9",
    x"3F67F48",
    x"3F67BA9",
    x"3F6780B",
    x"3F6746D",
    x"3F670D0",
    x"3F66D35",
    x"3F6699A",
    x"3F66600",
    x"3F66267",
    x"3F65ECF",
    x"3F65B37",
    x"3F657A1",
    x"3F6540C",
    x"3F65077",
    x"3F64CE3",
    x"3F64951",
    x"3F645BF",
    x"3F6422E",
    x"3F63E9E",
    x"3F63B0E",
    x"3F63780",
    x"3F633F3",
    x"3F63066",
    x"3F62CDA",
    x"3F62950",
    x"3F625C6",
    x"3F6223D",
    x"3F61EB5",
    x"3F61B2D",
    x"3F617A7",
    x"3F61422",
    x"3F6109D",
    x"3F60D19",
    x"3F60996",
    x"3F60614",
    x"3F60293",
    x"3F5FF13",
    x"3F5FB94",
    x"3F5F815",
    x"3F5F498",
    x"3F5F11B",
    x"3F5ED9F",
    x"3F5EA24",
    x"3F5E6AA",
    x"3F5E331",
    x"3F5DFB9",
    x"3F5DC41",
    x"3F5D8CA",
    x"3F5D555",
    x"3F5D1E0",
    x"3F5CE6C",
    x"3F5CAF9",
    x"3F5C786",
    x"3F5C415",
    x"3F5C0A4",
    x"3F5BD34",
    x"3F5B9C6",
    x"3F5B658",
    x"3F5B2EA",
    x"3F5AF7E",
    x"3F5AC13",
    x"3F5A8A8",
    x"3F5A53E",
    x"3F5A1D5",
    x"3F59E6D",
    x"3F59B06",
    x"3F597A0",
    x"3F5943A",
    x"3F590D6",
    x"3F58D72",
    x"3F58A0F",
    x"3F586AD",
    x"3F5834C",
    x"3F57FEB",
    x"3F57C8C",
    x"3F5792D",
    x"3F575CF",
    x"3F57272",
    x"3F56F16",
    x"3F56BBB",
    x"3F56860",
    x"3F56506",
    x"3F561AE",
    x"3F55E56",
    x"3F55AFE",
    x"3F557A8",
    x"3F55453",
    x"3F550FE",
    x"3F54DAA",
    x"3F54A57",
    x"3F54705",
    x"3F543B4",
    x"3F54063",
    x"3F53D13",
    x"3F539C5",
    x"3F53676",
    x"3F53329",
    x"3F52FDD",
    x"3F52C91",
    x"3F52947",
    x"3F525FD",
    x"3F522B4",
    x"3F51F6B",
    x"3F51C24",
    x"3F518DD",
    x"3F51597",
    x"3F51252",
    x"3F50F0E",
    x"3F50BCB",
    x"3F50888",
    x"3F50547",
    x"3F50206",
    x"3F4FEC6",
    x"3F4FB86",
    x"3F4F848",
    x"3F4F50A",
    x"3F4F1CD",
    x"3F4EE91",
    x"3F4EB56",
    x"3F4E81C",
    x"3F4E4E2",
    x"3F4E1A9",
    x"3F4DE71",
    x"3F4DB3A",
    x"3F4D804",
    x"3F4D4CE",
    x"3F4D199",
    x"3F4CE65",
    x"3F4CB32",
    x"3F4C800",
    x"3F4C4CE",
    x"3F4C19D",
    x"3F4BE6D",
    x"3F4BB3E",
    x"3F4B810",
    x"3F4B4E2",
    x"3F4B1B5",
    x"3F4AE89",
    x"3F4AB5E",
    x"3F4A833",
    x"3F4A50A",
    x"3F4A1E1",
    x"3F49EB9",
    x"3F49B92",
    x"3F4986B",
    x"3F49545",
    x"3F49220",
    x"3F48EFC",
    x"3F48BD9",
    x"3F488B6",
    x"3F48595",
    x"3F48274",
    x"3F47F53",
    x"3F47C34",
    x"3F47915",
    x"3F475F7",
    x"3F472DA",
    x"3F46FBE",
    x"3F46CA2",
    x"3F46988",
    x"3F4666E",
    x"3F46354",
    x"3F4603C",
    x"3F45D24",
    x"3F45A0D",
    x"3F456F7",
    x"3F453E2",
    x"3F450CD",
    x"3F44DB9",
    x"3F44AA6",
    x"3F44794",
    x"3F44483",
    x"3F44172",
    x"3F43E62",
    x"3F43B53",
    x"3F43844",
    x"3F43537",
    x"3F4322A",
    x"3F42F1D",
    x"3F42C12",
    x"3F42907",
    x"3F425FE",
    x"3F422F4",
    x"3F41FEC",
    x"3F41CE4",
    x"3F419DE",
    x"3F416D8",
    x"3F413D2",
    x"3F410CE",
    x"3F40DCA",
    x"3F40AC7",
    x"3F407C4",
    x"3F404C3",
    x"3F401C2",
    x"3F3FEC2",
    x"3F3FBC3",
    x"3F3F8C4",
    x"3F3F5C6",
    x"3F3F2C9",
    x"3F3EFCD",
    x"3F3ECD1",
    x"3F3E9D6",
    x"3F3E6DC",
    x"3F3E3E3",
    x"3F3E0EA",
    x"3F3DDF3",
    x"3F3DAFB",
    x"3F3D805",
    x"3F3D50F",
    x"3F3D21B",
    x"3F3CF26",
    x"3F3CC33",
    x"3F3C940",
    x"3F3C64E",
    x"3F3C35D",
    x"3F3C06D",
    x"3F3BD7D",
    x"3F3BA8E",
    x"3F3B7A0",
    x"3F3B4B2",
    x"3F3B1C5",
    x"3F3AED9",
    x"3F3ABEE",
    x"3F3A903",
    x"3F3A619",
    x"3F3A330",
    x"3F3A048",
    x"3F39D60",
    x"3F39A79",
    x"3F39793",
    x"3F394AD",
    x"3F391C8",
    x"3F38EE4",
    x"3F38C01",
    x"3F3891E",
    x"3F3863C",
    x"3F3835B",
    x"3F3807B",
    x"3F37D9B",
    x"3F37ABC",
    x"3F377DE",
    x"3F37500",
    x"3F37223",
    x"3F36F47",
    x"3F36C6C",
    x"3F36991",
    x"3F366B7",
    x"3F363DD",
    x"3F36105",
    x"3F35E2D",
    x"3F35B56",
    x"3F3587F",
    x"3F355A9",
    x"3F352D4",
    x"3F35000",
    x"3F34D2C",
    x"3F34A59",
    x"3F34787",
    x"3F344B6",
    x"3F341E5",
    x"3F33F15",
    x"3F33C45",
    x"3F33977",
    x"3F336A9",
    x"3F333DB",
    x"3F3310F",
    x"3F32E43",
    x"3F32B78",
    x"3F328AD",
    x"3F325E3",
    x"3F3231A",
    x"3F32052",
    x"3F31D8A",
    x"3F31AC3",
    x"3F317FD",
    x"3F31537",
    x"3F31272",
    x"3F30FAE",
    x"3F30CEA",
    x"3F30A27",
    x"3F30765",
    x"3F304A4",
    x"3F301E3",
    x"3F2FF23",
    x"3F2FC63",
    x"3F2F9A4",
    x"3F2F6E6",
    x"3F2F429",
    x"3F2F16C",
    x"3F2EEB0",
    x"3F2EBF5",
    x"3F2E93A",
    x"3F2E680",
    x"3F2E3C7",
    x"3F2E10E",
    x"3F2DE56",
    x"3F2DB9F",
    x"3F2D8E9",
    x"3F2D633",
    x"3F2D37E",
    x"3F2D0C9",
    x"3F2CE15",
    x"3F2CB62",
    x"3F2C8AF",
    x"3F2C5FE",
    x"3F2C34C",
    x"3F2C09C",
    x"3F2BDEC",
    x"3F2BB3D",
    x"3F2B88F",
    x"3F2B5E1",
    x"3F2B334",
    x"3F2B087",
    x"3F2ADDB",
    x"3F2AB30",
    x"3F2A886",
    x"3F2A5DC",
    x"3F2A333",
    x"3F2A08A",
    x"3F29DE3",
    x"3F29B3B",
    x"3F29895",
    x"3F295EF",
    x"3F2934A",
    x"3F290A5",
    x"3F28E02",
    x"3F28B5E",
    x"3F288BC",
    x"3F2861A",
    x"3F28379",
    x"3F280D8",
    x"3F27E38",
    x"3F27B99",
    x"3F278FB",
    x"3F2765D",
    x"3F273BF",
    x"3F27123",
    x"3F26E87",
    x"3F26BEC",
    x"3F26951",
    x"3F266B7",
    x"3F2641E",
    x"3F26185",
    x"3F25EED",
    x"3F25C55",
    x"3F259BF",
    x"3F25729",
    x"3F25493",
    x"3F251FE",
    x"3F24F6A",
    x"3F24CD7",
    x"3F24A44",
    x"3F247B1",
    x"3F24520",
    x"3F2428F",
    x"3F23FFF",
    x"3F23D6F",
    x"3F23AE0",
    x"3F23851",
    x"3F235C4",
    x"3F23337",
    x"3F230AA",
    x"3F22E1E",
    x"3F22B93",
    x"3F22908",
    x"3F2267E",
    x"3F223F5",
    x"3F2216C",
    x"3F21EE4",
    x"3F21C5D",
    x"3F219D6",
    x"3F21750",
    x"3F214CB",
    x"3F21246",
    x"3F20FC1",
    x"3F20D3E",
    x"3F20ABB",
    x"3F20838",
    x"3F205B7",
    x"3F20336",
    x"3F200B5",
    x"3F1FE35",
    x"3F1FBB6",
    x"3F1F937",
    x"3F1F6B9",
    x"3F1F43C",
    x"3F1F1BF",
    x"3F1EF43",
    x"3F1ECC8",
    x"3F1EA4D",
    x"3F1E7D3",
    x"3F1E559",
    x"3F1E2E0",
    x"3F1E067",
    x"3F1DDF0",
    x"3F1DB78",
    x"3F1D902",
    x"3F1D68C",
    x"3F1D417",
    x"3F1D1A2",
    x"3F1CF2E",
    x"3F1CCBA",
    x"3F1CA47",
    x"3F1C7D5",
    x"3F1C564",
    x"3F1C2F2",
    x"3F1C082",
    x"3F1BE12",
    x"3F1BBA3",
    x"3F1B934",
    x"3F1B6C6",
    x"3F1B459",
    x"3F1B1EC",
    x"3F1AF80",
    x"3F1AD14",
    x"3F1AAAA",
    x"3F1A83F",
    x"3F1A5D5",
    x"3F1A36C",
    x"3F1A104",
    x"3F19E9C",
    x"3F19C34",
    x"3F199CE",
    x"3F19767",
    x"3F19502",
    x"3F1929D",
    x"3F19039",
    x"3F18DD5",
    x"3F18B72",
    x"3F1890F",
    x"3F186AD",
    x"3F1844C",
    x"3F181EB",
    x"3F17F8B",
    x"3F17D2B",
    x"3F17ACC",
    x"3F1786E",
    x"3F17610",
    x"3F173B3",
    x"3F17156",
    x"3F16EFA",
    x"3F16C9F",
    x"3F16A44",
    x"3F167EA",
    x"3F16590",
    x"3F16337",
    x"3F160DE",
    x"3F15E86",
    x"3F15C2F",
    x"3F159D8",
    x"3F15782",
    x"3F1552C",
    x"3F152D7",
    x"3F15083",
    x"3F14E2F",
    x"3F14BDC",
    x"3F14989",
    x"3F14737",
    x"3F144E6",
    x"3F14295",
    x"3F14044",
    x"3F13DF5",
    x"3F13BA5",
    x"3F13957",
    x"3F13709",
    x"3F134BB",
    x"3F1326E",
    x"3F13022",
    x"3F12DD6",
    x"3F12B8B",
    x"3F12941",
    x"3F126F7",
    x"3F124AD",
    x"3F12264",
    x"3F1201C",
    x"3F11DD4",
    x"3F11B8D",
    x"3F11946",
    x"3F11700",
    x"3F114BB",
    x"3F11276",
    x"3F11032",
    x"3F10DEE",
    x"3F10BAB",
    x"3F10968",
    x"3F10726",
    x"3F104E4",
    x"3F102A3",
    x"3F10063",
    x"3F0FE23",
    x"3F0FBE4",
    x"3F0F9A5",
    x"3F0F767",
    x"3F0F52A",
    x"3F0F2ED",
    x"3F0F0B0",
    x"3F0EE74",
    x"3F0EC39",
    x"3F0E9FE",
    x"3F0E7C4",
    x"3F0E58A",
    x"3F0E351",
    x"3F0E119",
    x"3F0DEE1",
    x"3F0DCA9",
    x"3F0DA72",
    x"3F0D83C",
    x"3F0D606",
    x"3F0D3D1",
    x"3F0D19C",
    x"3F0CF68",
    x"3F0CD35",
    x"3F0CB02",
    x"3F0C8CF",
    x"3F0C69D",
    x"3F0C46C",
    x"3F0C23B",
    x"3F0C00B",
    x"3F0BDDB",
    x"3F0BBAC",
    x"3F0B97D",
    x"3F0B74F",
    x"3F0B521",
    x"3F0B2F4",
    x"3F0B0C8",
    x"3F0AE9C",
    x"3F0AC71",
    x"3F0AA46",
    x"3F0A81C",
    x"3F0A5F2",
    x"3F0A3C9",
    x"3F0A1A0",
    x"3F09F78",
    x"3F09D50",
    x"3F09B29",
    x"3F09903",
    x"3F096DD",
    x"3F094B7",
    x"3F09292",
    x"3F0906E",
    x"3F08E4A",
    x"3F08C27",
    x"3F08A04",
    x"3F087E2",
    x"3F085C0",
    x"3F0839F",
    x"3F0817E",
    x"3F07F5E",
    x"3F07D3E",
    x"3F07B1F",
    x"3F07901",
    x"3F076E3",
    x"3F074C5",
    x"3F072A9",
    x"3F0708C",
    x"3F06E70",
    x"3F06C55",
    x"3F06A3A",
    x"3F06820",
    x"3F06606",
    x"3F063ED",
    x"3F061D4",
    x"3F05FBC",
    x"3F05DA4",
    x"3F05B8D",
    x"3F05976",
    x"3F05760",
    x"3F0554B",
    x"3F05336",
    x"3F05121",
    x"3F04F0D",
    x"3F04CFA",
    x"3F04AE7",
    x"3F048D4",
    x"3F046C2",
    x"3F044B1",
    x"3F042A0",
    x"3F0408F",
    x"3F03E80",
    x"3F03C70",
    x"3F03A61",
    x"3F03853",
    x"3F03645",
    x"3F03438",
    x"3F0322B",
    x"3F0301F",
    x"3F02E13",
    x"3F02C08",
    x"3F029FD",
    x"3F027F3",
    x"3F025E9",
    x"3F023E0",
    x"3F021D7",
    x"3F01FCF",
    x"3F01DC7",
    x"3F01BC0",
    x"3F019B9",
    x"3F017B3",
    x"3F015AD",
    x"3F013A8",
    x"3F011A4",
    x"3F00F9F",
    x"3F00D9C",
    x"3F00B99",
    x"3F00996",
    x"3F00794",
    x"3F00592",
    x"3F00391",
    x"3F00190",
    x"3EFFF21",
    x"3EFFB22",
    x"3EFF723",
    x"3EFF326",
    x"3EFEF2A",
    x"3EFEB2F",
    x"3EFE734",
    x"3EFE33B",
    x"3EFDF43",
    x"3EFDB4B",
    x"3EFD755",
    x"3EFD360",
    x"3EFCF6B",
    x"3EFCB78",
    x"3EFC786",
    x"3EFC394",
    x"3EFBFA4",
    x"3EFBBB4",
    x"3EFB7C6",
    x"3EFB3D9",
    x"3EFAFEC",
    x"3EFAC01",
    x"3EFA816",
    x"3EFA42D",
    x"3EFA044",
    x"3EF9C5C",
    x"3EF9876",
    x"3EF9490",
    x"3EF90AC",
    x"3EF8CC8",
    x"3EF88E5",
    x"3EF8503",
    x"3EF8123",
    x"3EF7D43",
    x"3EF7964",
    x"3EF7586",
    x"3EF71A9",
    x"3EF6DCD",
    x"3EF69F2",
    x"3EF6618",
    x"3EF623F",
    x"3EF5E67",
    x"3EF5A90",
    x"3EF56BA",
    x"3EF52E5",
    x"3EF4F10",
    x"3EF4B3D",
    x"3EF476B",
    x"3EF4399",
    x"3EF3FC9",
    x"3EF3BFA",
    x"3EF382B",
    x"3EF345D",
    x"3EF3091",
    x"3EF2CC5",
    x"3EF28FA",
    x"3EF2531",
    x"3EF2168",
    x"3EF1DA0",
    x"3EF19D9",
    x"3EF1613",
    x"3EF124E",
    x"3EF0E8A",
    x"3EF0AC7",
    x"3EF0705",
    x"3EF0343",
    x"3EEFF83",
    x"3EEFBC3",
    x"3EEF805",
    x"3EEF447",
    x"3EEF08B",
    x"3EEECCF",
    x"3EEE914",
    x"3EEE55B",
    x"3EEE1A2",
    x"3EEDDEA",
    x"3EEDA33",
    x"3EED67D",
    x"3EED2C8",
    x"3EECF13",
    x"3EECB60",
    x"3EEC7AE",
    x"3EEC3FC",
    x"3EEC04C",
    x"3EEBC9C",
    x"3EEB8ED",
    x"3EEB540",
    x"3EEB193",
    x"3EEADE7",
    x"3EEAA3C",
    x"3EEA692",
    x"3EEA2E8",
    x"3EE9F40",
    x"3EE9B99",
    x"3EE97F2",
    x"3EE944D",
    x"3EE90A8",
    x"3EE8D05",
    x"3EE8962",
    x"3EE85C0",
    x"3EE821F",
    x"3EE7E7F",
    x"3EE7AE0",
    x"3EE7741",
    x"3EE73A4",
    x"3EE7008",
    x"3EE6C6C",
    x"3EE68D1",
    x"3EE6538",
    x"3EE619F",
    x"3EE5E07",
    x"3EE5A70",
    x"3EE56DA",
    x"3EE5344",
    x"3EE4FB0",
    x"3EE4C1C",
    x"3EE488A",
    x"3EE44F8",
    x"3EE4167",
    x"3EE3DD7",
    x"3EE3A48",
    x"3EE36BA",
    x"3EE332D",
    x"3EE2FA1",
    x"3EE2C15",
    x"3EE288B",
    x"3EE2501",
    x"3EE2178",
    x"3EE1DF0",
    x"3EE1A69",
    x"3EE16E3",
    x"3EE135E",
    x"3EE0FD9",
    x"3EE0C56",
    x"3EE08D3",
    x"3EE0551",
    x"3EE01D1",
    x"3EDFE51",
    x"3EDFAD1",
    x"3EDF753",
    x"3EDF3D6",
    x"3EDF059",
    x"3EDECDE",
    x"3EDE963",
    x"3EDE5E9",
    x"3EDE270",
    x"3EDDEF8",
    x"3EDDB80",
    x"3EDD80A",
    x"3EDD494",
    x"3EDD120",
    x"3EDCDAC",
    x"3EDCA39",
    x"3EDC6C7",
    x"3EDC355",
    x"3EDBFE5",
    x"3EDBC75",
    x"3EDB907",
    x"3EDB599",
    x"3EDB22C",
    x"3EDAEC0",
    x"3EDAB55",
    x"3EDA7EA",
    x"3EDA481",
    x"3EDA118",
    x"3ED9DB0",
    x"3ED9A49",
    x"3ED96E3",
    x"3ED937E",
    x"3ED9019",
    x"3ED8CB6",
    x"3ED8953",
    x"3ED85F1",
    x"3ED8290",
    x"3ED7F30",
    x"3ED7BD0",
    x"3ED7872",
    x"3ED7514",
    x"3ED71B7",
    x"3ED6E5B",
    x"3ED6B00",
    x"3ED67A6",
    x"3ED644C",
    x"3ED60F4",
    x"3ED5D9C",
    x"3ED5A45",
    x"3ED56EF",
    x"3ED5399",
    x"3ED5045",
    x"3ED4CF1",
    x"3ED499E",
    x"3ED464C",
    x"3ED42FB",
    x"3ED3FAB",
    x"3ED3C5B",
    x"3ED390D",
    x"3ED35BF",
    x"3ED3272",
    x"3ED2F26",
    x"3ED2BDA",
    x"3ED2890",
    x"3ED2546",
    x"3ED21FD",
    x"3ED1EB5",
    x"3ED1B6E",
    x"3ED1827",
    x"3ED14E2",
    x"3ED119D",
    x"3ED0E59",
    x"3ED0B16",
    x"3ED07D3",
    x"3ED0492",
    x"3ED0151",
    x"3ECFE11",
    x"3ECFAD2",
    x"3ECF794",
    x"3ECF456",
    x"3ECF119",
    x"3ECEDDE",
    x"3ECEAA2",
    x"3ECE768",
    x"3ECE42F",
    x"3ECE0F6",
    x"3ECDDBE",
    x"3ECDA87",
    x"3ECD751",
    x"3ECD41C",
    x"3ECD0E7",
    x"3ECCDB3",
    x"3ECCA80",
    x"3ECC74E",
    x"3ECC41C",
    x"3ECC0EC",
    x"3ECBDBC",
    x"3ECBA8D",
    x"3ECB75F",
    x"3ECB431",
    x"3ECB105",
    x"3ECADD9",
    x"3ECAAAE",
    x"3ECA783",
    x"3ECA45A",
    x"3ECA131",
    x"3EC9E09",
    x"3EC9AE2",
    x"3EC97BC",
    x"3EC9496",
    x"3EC9172",
    x"3EC8E4E",
    x"3EC8B2A",
    x"3EC8808",
    x"3EC84E6",
    x"3EC81C6",
    x"3EC7EA6",
    x"3EC7B86",
    x"3EC7868",
    x"3EC754A",
    x"3EC722D",
    x"3EC6F11",
    x"3EC6BF6",
    x"3EC68DB",
    x"3EC65C1",
    x"3EC62A8",
    x"3EC5F90",
    x"3EC5C78",
    x"3EC5962",
    x"3EC564C",
    x"3EC5336",
    x"3EC5022",
    x"3EC4D0E",
    x"3EC49FC",
    x"3EC46E9",
    x"3EC43D8",
    x"3EC40C7",
    x"3EC3DB8",
    x"3EC3AA9",
    x"3EC379A",
    x"3EC348D",
    x"3EC3180",
    x"3EC2E74",
    x"3EC2B69",
    x"3EC285E",
    x"3EC2555",
    x"3EC224C",
    x"3EC1F43",
    x"3EC1C3C",
    x"3EC1935",
    x"3EC162F",
    x"3EC132A",
    x"3EC1026",
    x"3EC0D22",
    x"3EC0A1F",
    x"3EC071D",
    x"3EC041C",
    x"3EC011B",
    x"3EBFE1B",
    x"3EBFB1C",
    x"3EBF81E",
    x"3EBF520",
    x"3EBF223",
    x"3EBEF27",
    x"3EBEC2B",
    x"3EBE931",
    x"3EBE637",
    x"3EBE33E",
    x"3EBE045",
    x"3EBDD4E",
    x"3EBDA57",
    x"3EBD760",
    x"3EBD46B",
    x"3EBD176",
    x"3EBCE82",
    x"3EBCB8F",
    x"3EBC89C",
    x"3EBC5AB",
    x"3EBC2BA",
    x"3EBBFC9",
    x"3EBBCDA",
    x"3EBB9EB",
    x"3EBB6FD",
    x"3EBB40F",
    x"3EBB123",
    x"3EBAE37",
    x"3EBAB4C",
    x"3EBA861",
    x"3EBA577",
    x"3EBA28E",
    x"3EB9FA6",
    x"3EB9CBF",
    x"3EB99D8",
    x"3EB96F2",
    x"3EB940C",
    x"3EB9128",
    x"3EB8E44",
    x"3EB8B60",
    x"3EB887E",
    x"3EB859C",
    x"3EB82BB",
    x"3EB7FDB",
    x"3EB7CFB",
    x"3EB7A1C",
    x"3EB773E",
    x"3EB7461",
    x"3EB7184",
    x"3EB6EA8",
    x"3EB6BCD",
    x"3EB68F2",
    x"3EB6618",
    x"3EB633F",
    x"3EB6067",
    x"3EB5D8F",
    x"3EB5AB8",
    x"3EB57E1",
    x"3EB550C",
    x"3EB5237",
    x"3EB4F63",
    x"3EB4C8F",
    x"3EB49BC",
    x"3EB46EA",
    x"3EB4419",
    x"3EB4148",
    x"3EB3E78",
    x"3EB3BA9",
    x"3EB38DB",
    x"3EB360D",
    x"3EB3340",
    x"3EB3073",
    x"3EB2DA7",
    x"3EB2ADC",
    x"3EB2812",
    x"3EB2548",
    x"3EB227F",
    x"3EB1FB7",
    x"3EB1CEF",
    x"3EB1A28",
    x"3EB1762",
    x"3EB149D",
    x"3EB11D8",
    x"3EB0F14",
    x"3EB0C50",
    x"3EB098E",
    x"3EB06CC",
    x"3EB040A",
    x"3EB014A",
    x"3EAFE8A",
    x"3EAFBCA",
    x"3EAF90C",
    x"3EAF64E",
    x"3EAF391",
    x"3EAF0D4",
    x"3EAEE18",
    x"3EAEB5D",
    x"3EAE8A3",
    x"3EAE5E9",
    x"3EAE330",
    x"3EAE077",
    x"3EADDBF",
    x"3EADB08",
    x"3EAD852",
    x"3EAD59C",
    x"3EAD2E7",
    x"3EAD033",
    x"3EACD7F",
    x"3EACACC",
    x"3EAC81A",
    x"3EAC568",
    x"3EAC2B7",
    x"3EAC006",
    x"3EABD57",
    x"3EABAA8",
    x"3EAB7F9",
    x"3EAB54C",
    x"3EAB29F",
    x"3EAAFF2",
    x"3EAAD47",
    x"3EAAA9C",
    x"3EAA7F2",
    x"3EAA548",
    x"3EAA29F",
    x"3EA9FF7",
    x"3EA9D4F",
    x"3EA9AA8",
    x"3EA9802",
    x"3EA955C",
    x"3EA92B7",
    x"3EA9013",
    x"3EA8D6F",
    x"3EA8ACC",
    x"3EA8829",
    x"3EA8588",
    x"3EA82E7",
    x"3EA8046",
    x"3EA7DA7",
    x"3EA7B07",
    x"3EA7869",
    x"3EA75CB",
    x"3EA732E",
    x"3EA7092",
    x"3EA6DF6",
    x"3EA6B5B",
    x"3EA68C0",
    x"3EA6626",
    x"3EA638D",
    x"3EA60F5",
    x"3EA5E5D",
    x"3EA5BC5",
    x"3EA592F",
    x"3EA5699",
    x"3EA5403",
    x"3EA516F",
    x"3EA4EDB",
    x"3EA4C47",
    x"3EA49B5",
    x"3EA4722",
    x"3EA4491",
    x"3EA4200",
    x"3EA3F70",
    x"3EA3CE0",
    x"3EA3A52",
    x"3EA37C3",
    x"3EA3536",
    x"3EA32A9",
    x"3EA301C",
    x"3EA2D91",
    x"3EA2B06",
    x"3EA287B",
    x"3EA25F1",
    x"3EA2368",
    x"3EA20E0",
    x"3EA1E58",
    x"3EA1BD0",
    x"3EA194A",
    x"3EA16C4",
    x"3EA143E",
    x"3EA11BA",
    x"3EA0F36",
    x"3EA0CB2",
    x"3EA0A2F",
    x"3EA07AD",
    x"3EA052B",
    x"3EA02AA",
    x"3EA002A",
    x"3E9FDAA",
    x"3E9FB2B",
    x"3E9F8AD",
    x"3E9F62F",
    x"3E9F3B2",
    x"3E9F135",
    x"3E9EEB9",
    x"3E9EC3E",
    x"3E9E9C3",
    x"3E9E749",
    x"3E9E4CF",
    x"3E9E256",
    x"3E9DFDE",
    x"3E9DD66",
    x"3E9DAEF",
    x"3E9D879",
    x"3E9D603",
    x"3E9D38E",
    x"3E9D119",
    x"3E9CEA5",
    x"3E9CC32",
    x"3E9C9BF",
    x"3E9C74D",
    x"3E9C4DC",
    x"3E9C26B",
    x"3E9BFFA",
    x"3E9BD8B",
    x"3E9BB1C",
    x"3E9B8AD",
    x"3E9B63F",
    x"3E9B3D2",
    x"3E9B165",
    x"3E9AEF9",
    x"3E9AC8E",
    x"3E9AA23",
    x"3E9A7B9",
    x"3E9A54F",
    x"3E9A2E6",
    x"3E9A07E",
    x"3E99E16",
    x"3E99BAF",
    x"3E99948",
    x"3E996E2",
    x"3E9947D",
    x"3E99218",
    x"3E98FB4",
    x"3E98D50",
    x"3E98AED",
    x"3E9888B",
    x"3E98629",
    x"3E983C7",
    x"3E98167",
    x"3E97F07",
    x"3E97CA7",
    x"3E97A48",
    x"3E977EA",
    x"3E9758C",
    x"3E9732F",
    x"3E970D3",
    x"3E96E77",
    x"3E96C1C",
    x"3E969C1",
    x"3E96767",
    x"3E9650D",
    x"3E962B4",
    x"3E9605C",
    x"3E95E04",
    x"3E95BAD",
    x"3E95956",
    x"3E95700",
    x"3E954AB",
    x"3E95256",
    x"3E95002",
    x"3E94DAE",
    x"3E94B5B",
    x"3E94908",
    x"3E946B6",
    x"3E94465",
    x"3E94214",
    x"3E93FC4",
    x"3E93D74",
    x"3E93B25",
    x"3E938D7",
    x"3E93689",
    x"3E9343B",
    x"3E931EF",
    x"3E92FA2",
    x"3E92D57",
    x"3E92B0C",
    x"3E928C1",
    x"3E92677",
    x"3E9242E",
    x"3E921E5",
    x"3E91F9D",
    x"3E91D55",
    x"3E91B0E",
    x"3E918C8",
    x"3E91682",
    x"3E9143D",
    x"3E911F8",
    x"3E90FB4",
    x"3E90D70",
    x"3E90B2D",
    x"3E908EA",
    x"3E906A8",
    x"3E90467",
    x"3E90226",
    x"3E8FFE6",
    x"3E8FDA6",
    x"3E8FB67",
    x"3E8F929",
    x"3E8F6EB",
    x"3E8F4AD",
    x"3E8F270",
    x"3E8F034",
    x"3E8EDF8",
    x"3E8EBBD",
    x"3E8E982",
    x"3E8E748",
    x"3E8E50F",
    x"3E8E2D6",
    x"3E8E09D",
    x"3E8DE65",
    x"3E8DC2E",
    x"3E8D9F7",
    x"3E8D7C1",
    x"3E8D58B",
    x"3E8D356",
    x"3E8D122",
    x"3E8CEEE",
    x"3E8CCBA",
    x"3E8CA87",
    x"3E8C855",
    x"3E8C623",
    x"3E8C3F2",
    x"3E8C1C1",
    x"3E8BF91",
    x"3E8BD61",
    x"3E8BB32",
    x"3E8B904",
    x"3E8B6D6",
    x"3E8B4A8",
    x"3E8B27B",
    x"3E8B04F",
    x"3E8AE23",
    x"3E8ABF8",
    x"3E8A9CD",
    x"3E8A7A3",
    x"3E8A579",
    x"3E8A350",
    x"3E8A128",
    x"3E89F00",
    x"3E89CD8",
    x"3E89AB1",
    x"3E8988B",
    x"3E89665",
    x"3E89440",
    x"3E8921B",
    x"3E88FF7",
    x"3E88DD3",
    x"3E88BB0",
    x"3E8898D",
    x"3E8876B",
    x"3E88549",
    x"3E88328",
    x"3E88108",
    x"3E87EE8",
    x"3E87CC8",
    x"3E87AA9",
    x"3E8788B",
    x"3E8766D",
    x"3E87450",
    x"3E87233",
    x"3E87017",
    x"3E86DFB",
    x"3E86BE0",
    x"3E869C5",
    x"3E867AB",
    x"3E86591",
    x"3E86378",
    x"3E86160",
    x"3E85F47",
    x"3E85D30",
    x"3E85B19",
    x"3E85902",
    x"3E856EC",
    x"3E854D7",
    x"3E852C2",
    x"3E850AD",
    x"3E84E9A",
    x"3E84C86",
    x"3E84A73",
    x"3E84861",
    x"3E8464F",
    x"3E8443E",
    x"3E8422D",
    x"3E8401D",
    x"3E83E0D",
    x"3E83BFE",
    x"3E839EF",
    x"3E837E1",
    x"3E835D3",
    x"3E833C6",
    x"3E831B9",
    x"3E82FAD",
    x"3E82DA1",
    x"3E82B96",
    x"3E8298B",
    x"3E82781",
    x"3E82578",
    x"3E8236F",
    x"3E82166",
    x"3E81F5E",
    x"3E81D56",
    x"3E81B4F",
    x"3E81949",
    x"3E81743",
    x"3E8153D",
    x"3E81338",
    x"3E81133",
    x"3E80F2F",
    x"3E80D2C",
    x"3E80B29",
    x"3E80926",
    x"3E80724",
    x"3E80523",
    x"3E80322",
    x"3E80121",
    x"3E7FE43",
    x"3E7FA44",
    x"3E7F645",
    x"3E7F248",
    x"3E7EE4C",
    x"3E7EA51",
    x"3E7E657",
    x"3E7E25E",
    x"3E7DE66",
    x"3E7DA6F",
    x"3E7D679",
    x"3E7D284",
    x"3E7CE90",
    x"3E7CA9C",
    x"3E7C6AA",
    x"3E7C2B9",
    x"3E7BEC9",
    x"3E7BADA",
    x"3E7B6EB",
    x"3E7B2FE",
    x"3E7AF12",
    x"3E7AB27",
    x"3E7A73C",
    x"3E7A353",
    x"3E79F6B",
    x"3E79B83",
    x"3E7979D",
    x"3E793B8",
    x"3E78FD3",
    x"3E78BF0",
    x"3E7880D",
    x"3E7842C",
    x"3E7804B",
    x"3E77C6B",
    x"3E7788D",
    x"3E774AF",
    x"3E770D2",
    x"3E76CF7",
    x"3E7691C",
    x"3E76542",
    x"3E76169",
    x"3E75D91",
    x"3E759BB",
    x"3E755E5",
    x"3E75210",
    x"3E74E3C",
    x"3E74A68",
    x"3E74696",
    x"3E742C5",
    x"3E73EF5",
    x"3E73B26",
    x"3E73757",
    x"3E7338A",
    x"3E72FBE",
    x"3E72BF2",
    x"3E72828",
    x"3E7245E",
    x"3E72095",
    x"3E71CCE",
    x"3E71907",
    x"3E71541",
    x"3E7117C",
    x"3E70DB9",
    x"3E709F6",
    x"3E70634",
    x"3E70272",
    x"3E6FEB2",
    x"3E6FAF3",
    x"3E6F735",
    x"3E6F378",
    x"3E6EFBB",
    x"3E6EC00",
    x"3E6E845",
    x"3E6E48C",
    x"3E6E0D3",
    x"3E6DD1B",
    x"3E6D964",
    x"3E6D5AE",
    x"3E6D1F9",
    x"3E6CE45",
    x"3E6CA92",
    x"3E6C6E0",
    x"3E6C32F",
    x"3E6BF7F",
    x"3E6BBCF",
    x"3E6B821",
    x"3E6B473",
    x"3E6B0C6",
    x"3E6AD1B",
    x"3E6A970",
    x"3E6A5C6",
    x"3E6A21D",
    x"3E69E75",
    x"3E69ACE",
    x"3E69728",
    x"3E69382",
    x"3E68FDE",
    x"3E68C3A",
    x"3E68898",
    x"3E684F6",
    x"3E68155",
    x"3E67DB5",
    x"3E67A16",
    x"3E67678",
    x"3E672DB",
    x"3E66F3F",
    x"3E66BA3",
    x"3E66809",
    x"3E6646F",
    x"3E660D7",
    x"3E65D3F",
    x"3E659A8",
    x"3E65612",
    x"3E6527D",
    x"3E64EE9",
    x"3E64B56",
    x"3E647C3",
    x"3E64432",
    x"3E640A1",
    x"3E63D11",
    x"3E63983",
    x"3E635F5",
    x"3E63268",
    x"3E62EDB",
    x"3E62B50",
    x"3E627C6",
    x"3E6243C",
    x"3E620B4",
    x"3E61D2C",
    x"3E619A5",
    x"3E6161F",
    x"3E6129A",
    x"3E60F16",
    x"3E60B93",
    x"3E60810",
    x"3E6048E",
    x"3E6010E",
    x"3E5FD8E",
    x"3E5FA0F",
    x"3E5F691",
    x"3E5F314",
    x"3E5EF97",
    x"3E5EC1C",
    x"3E5E8A1",
    x"3E5E528",
    x"3E5E1AF",
    x"3E5DE37",
    x"3E5DAC0",
    x"3E5D749",
    x"3E5D3D4",
    x"3E5D05F",
    x"3E5CCEC",
    x"3E5C979",
    x"3E5C607",
    x"3E5C296",
    x"3E5BF26",
    x"3E5BBB6",
    x"3E5B848",
    x"3E5B4DA",
    x"3E5B16D",
    x"3E5AE02",
    x"3E5AA96",
    x"3E5A72C",
    x"3E5A3C3",
    x"3E5A05A",
    x"3E59CF3",
    x"3E5998C",
    x"3E59626",
    x"3E592C1",
    x"3E58F5D",
    x"3E58BF9",
    x"3E58897",
    x"3E58535",
    x"3E581D4",
    x"3E57E74",
    x"3E57B15",
    x"3E577B6",
    x"3E57459",
    x"3E570FC",
    x"3E56DA0",
    x"3E56A45",
    x"3E566EB",
    x"3E56392",
    x"3E56039",
    x"3E55CE2",
    x"3E5598B",
    x"3E55635",
    x"3E552E0",
    x"3E54F8C",
    x"3E54C38",
    x"3E548E6",
    x"3E54594",
    x"3E54243",
    x"3E53EF3",
    x"3E53BA3",
    x"3E53855",
    x"3E53507",
    x"3E531BA",
    x"3E52E6E",
    x"3E52B23",
    x"3E527D9",
    x"3E5248F",
    x"3E52146",
    x"3E51DFE",
    x"3E51AB7",
    x"3E51771",
    x"3E5142C",
    x"3E510E7",
    x"3E50DA3",
    x"3E50A60",
    x"3E5071E",
    x"3E503DD",
    x"3E5009C",
    x"3E4FD5C",
    x"3E4FA1D",
    x"3E4F6DF",
    x"3E4F3A2",
    x"3E4F065",
    x"3E4ED2A",
    x"3E4E9EF",
    x"3E4E6B5",
    x"3E4E37C",
    x"3E4E043",
    x"3E4DD0B",
    x"3E4D9D5",
    x"3E4D69E",
    x"3E4D369",
    x"3E4D035",
    x"3E4CD01",
    x"3E4C9CE",
    x"3E4C69C",
    x"3E4C36B",
    x"3E4C03A",
    x"3E4BD0B",
    x"3E4B9DC",
    x"3E4B6AE",
    x"3E4B381",
    x"3E4B054",
    x"3E4AD28",
    x"3E4A9FE",
    x"3E4A6D3",
    x"3E4A3AA",
    x"3E4A082",
    x"3E49D5A",
    x"3E49A33",
    x"3E4970D",
    x"3E493E7",
    x"3E490C3",
    x"3E48D9F",
    x"3E48A7C",
    x"3E4875A",
    x"3E48438",
    x"3E48118",
    x"3E47DF8",
    x"3E47AD9",
    x"3E477BA",
    x"3E4749D",
    x"3E47180",
    x"3E46E64",
    x"3E46B49",
    x"3E4682E",
    x"3E46515",
    x"3E461FC",
    x"3E45EE4",
    x"3E45BCC",
    x"3E458B6",
    x"3E455A0",
    x"3E4528B",
    x"3E44F77",
    x"3E44C63",
    x"3E44951",
    x"3E4463F",
    x"3E4432E",
    x"3E4401D",
    x"3E43D0D",
    x"3E439FF",
    x"3E436F0",
    x"3E433E3",
    x"3E430D7",
    x"3E42DCB",
    x"3E42AC0",
    x"3E427B5",
    x"3E424AC",
    x"3E421A3",
    x"3E41E9B",
    x"3E41B94",
    x"3E4188D",
    x"3E41587",
    x"3E41282",
    x"3E40F7E",
    x"3E40C7B",
    x"3E40978",
    x"3E40676",
    x"3E40375",
    x"3E40074",
    x"3E3FD74",
    x"3E3FA75",
    x"3E3F777",
    x"3E3F47A",
    x"3E3F17D",
    x"3E3EE81",
    x"3E3EB86",
    x"3E3E88B",
    x"3E3E591",
    x"3E3E298",
    x"3E3DFA0",
    x"3E3DCA9",
    x"3E3D9B2",
    x"3E3D6BC",
    x"3E3D3C6",
    x"3E3D0D2",
    x"3E3CDDE",
    x"3E3CAEB",
    x"3E3C7F9",
    x"3E3C507",
    x"3E3C216",
    x"3E3BF26",
    x"3E3BC36",
    x"3E3B948",
    x"3E3B65A",
    x"3E3B36D",
    x"3E3B080",
    x"3E3AD94",
    x"3E3AAA9",
    x"3E3A7BF",
    x"3E3A4D5",
    x"3E3A1ED",
    x"3E39F04",
    x"3E39C1D",
    x"3E39936",
    x"3E39650",
    x"3E3936B",
    x"3E39087",
    x"3E38DA3",
    x"3E38AC0",
    x"3E387DE",
    x"3E384FC",
    x"3E3821B",
    x"3E37F3B",
    x"3E37C5C",
    x"3E3797D",
    x"3E3769F",
    x"3E373C1",
    x"3E370E5",
    x"3E36E09",
    x"3E36B2E",
    x"3E36853",
    x"3E3657A",
    x"3E362A1",
    x"3E35FC8",
    x"3E35CF1",
    x"3E35A1A",
    x"3E35744",
    x"3E3546E",
    x"3E3519A",
    x"3E34EC6",
    x"3E34BF2",
    x"3E34920",
    x"3E3464E",
    x"3E3437C",
    x"3E340AC",
    x"3E33DDC",
    x"3E33B0D",
    x"3E3383F",
    x"3E33571",
    x"3E332A4",
    x"3E32FD7",
    x"3E32D0C",
    x"3E32A41",
    x"3E32777",
    x"3E324AD",
    x"3E321E4",
    x"3E31F1C",
    x"3E31C55",
    x"3E3198E",
    x"3E316C8",
    x"3E31403",
    x"3E3113E",
    x"3E30E7A",
    x"3E30BB7",
    x"3E308F4",
    x"3E30632",
    x"3E30371",
    x"3E300B1",
    x"3E2FDF1",
    x"3E2FB32",
    x"3E2F873",
    x"3E2F5B5",
    x"3E2F2F8",
    x"3E2F03C",
    x"3E2ED80",
    x"3E2EAC5",
    x"3E2E80B",
    x"3E2E551",
    x"3E2E298",
    x"3E2DFE0",
    x"3E2DD28",
    x"3E2DA71",
    x"3E2D7BB",
    x"3E2D505",
    x"3E2D251",
    x"3E2CF9C",
    x"3E2CCE9",
    x"3E2CA36",
    x"3E2C784",
    x"3E2C4D2",
    x"3E2C221",
    x"3E2BF71",
    x"3E2BCC1",
    x"3E2BA13",
    x"3E2B764",
    x"3E2B4B7",
    x"3E2B20A",
    x"3E2AF5E",
    x"3E2ACB2",
    x"3E2AA08",
    x"3E2A75D",
    x"3E2A4B4",
    x"3E2A20B",
    x"3E29F63",
    x"3E29CBB",
    x"3E29A14",
    x"3E2976E",
    x"3E294C9",
    x"3E29224",
    x"3E28F80",
    x"3E28CDC",
    x"3E28A39",
    x"3E28797",
    x"3E284F5",
    x"3E28255",
    x"3E27FB4",
    x"3E27D15",
    x"3E27A76",
    x"3E277D7",
    x"3E2753A",
    x"3E2729D",
    x"3E27001",
    x"3E26D65",
    x"3E26ACA",
    x"3E2682F",
    x"3E26596",
    x"3E262FD",
    x"3E26064",
    x"3E25DCC",
    x"3E25B35",
    x"3E2589F",
    x"3E25609",
    x"3E25374",
    x"3E250DF",
    x"3E24E4B",
    x"3E24BB8",
    x"3E24926",
    x"3E24694",
    x"3E24402",
    x"3E24172",
    x"3E23EE2",
    x"3E23C52",
    x"3E239C3",
    x"3E23735",
    x"3E234A8",
    x"3E2321B",
    x"3E22F8F",
    x"3E22D03",
    x"3E22A78",
    x"3E227EE",
    x"3E22564",
    x"3E222DB",
    x"3E22053",
    x"3E21DCB",
    x"3E21B44",
    x"3E218BD",
    x"3E21638",
    x"3E213B2",
    x"3E2112E",
    x"3E20EAA",
    x"3E20C26",
    x"3E209A4",
    x"3E20722",
    x"3E204A0",
    x"3E2021F",
    x"3E1FF9F",
    x"3E1FD1F",
    x"3E1FAA0",
    x"3E1F822",
    x"3E1F5A4",
    x"3E1F327",
    x"3E1F0AB",
    x"3E1EE2F",
    x"3E1EBB4",
    x"3E1E939",
    x"3E1E6BF",
    x"3E1E446",
    x"3E1E1CD",
    x"3E1DF55",
    x"3E1DCDD",
    x"3E1DA66",
    x"3E1D7F0",
    x"3E1D57A",
    x"3E1D305",
    x"3E1D091",
    x"3E1CE1D",
    x"3E1CBAA",
    x"3E1C937",
    x"3E1C6C5",
    x"3E1C454",
    x"3E1C1E3",
    x"3E1BF73",
    x"3E1BD03",
    x"3E1BA94",
    x"3E1B826",
    x"3E1B5B8",
    x"3E1B34B",
    x"3E1B0DF",
    x"3E1AE73",
    x"3E1AC07",
    x"3E1A99D",
    x"3E1A733",
    x"3E1A4C9",
    x"3E1A260",
    x"3E19FF8",
    x"3E19D90",
    x"3E19B29",
    x"3E198C3",
    x"3E1965D",
    x"3E193F7",
    x"3E19193",
    x"3E18F2F",
    x"3E18CCB",
    x"3E18A68",
    x"3E18806",
    x"3E185A4",
    x"3E18343",
    x"3E180E3",
    x"3E17E83",
    x"3E17C23",
    x"3E179C5",
    x"3E17767",
    x"3E17509",
    x"3E172AC",
    x"3E17050",
    x"3E16DF4",
    x"3E16B99",
    x"3E1693E",
    x"3E166E4",
    x"3E1648B",
    x"3E16232",
    x"3E15FD9",
    x"3E15D82",
    x"3E15B2B",
    x"3E158D4",
    x"3E1567E",
    x"3E15429",
    x"3E151D4",
    x"3E14F80",
    x"3E14D2C",
    x"3E14AD9",
    x"3E14887",
    x"3E14635",
    x"3E143E4",
    x"3E14193",
    x"3E13F43",
    x"3E13CF4",
    x"3E13AA5",
    x"3E13856",
    x"3E13609",
    x"3E133BB",
    x"3E1316F",
    x"3E12F23",
    x"3E12CD7",
    x"3E12A8C",
    x"3E12842",
    x"3E125F8",
    x"3E123AF",
    x"3E12166",
    x"3E11F1E",
    x"3E11CD7",
    x"3E11A90",
    x"3E11849",
    x"3E11604",
    x"3E113BE",
    x"3E1117A",
    x"3E10F36",
    x"3E10CF2",
    x"3E10AAF",
    x"3E1086D",
    x"3E1062B",
    x"3E103EA",
    x"3E101A9",
    x"3E0FF69",
    x"3E0FD29",
    x"3E0FAEA",
    x"3E0F8AC",
    x"3E0F66E",
    x"3E0F431",
    x"3E0F1F4",
    x"3E0EFB8",
    x"3E0ED7C",
    x"3E0EB41",
    x"3E0E906",
    x"3E0E6CC",
    x"3E0E493",
    x"3E0E25A",
    x"3E0E022",
    x"3E0DDEA",
    x"3E0DBB3",
    x"3E0D97C",
    x"3E0D746",
    x"3E0D510",
    x"3E0D2DC",
    x"3E0D0A7",
    x"3E0CE73",
    x"3E0CC40",
    x"3E0CA0D",
    x"3E0C7DB",
    x"3E0C5A9",
    x"3E0C378",
    x"3E0C147",
    x"3E0BF17",
    x"3E0BCE8",
    x"3E0BAB9",
    x"3E0B88A",
    x"3E0B65D",
    x"3E0B42F",
    x"3E0B203",
    x"3E0AFD6",
    x"3E0ADAB",
    x"3E0AB7F",
    x"3E0A955",
    x"3E0A72B",
    x"3E0A501",
    x"3E0A2D8",
    x"3E0A0B0",
    x"3E09E88",
    x"3E09C61",
    x"3E09A3A",
    x"3E09813",
    x"3E095EE",
    x"3E093C8",
    x"3E091A4",
    x"3E08F80",
    x"3E08D5C",
    x"3E08B39",
    x"3E08916",
    x"3E086F4",
    x"3E084D3",
    x"3E082B2",
    x"3E08092",
    x"3E07E72",
    x"3E07C52",
    x"3E07A34",
    x"3E07815",
    x"3E075F8",
    x"3E073DA",
    x"3E071BE",
    x"3E06FA1",
    x"3E06D86",
    x"3E06B6B",
    x"3E06950",
    x"3E06736",
    x"3E0651C",
    x"3E06303",
    x"3E060EB",
    x"3E05ED3",
    x"3E05CBC",
    x"3E05AA5",
    x"3E0588E",
    x"3E05678",
    x"3E05463",
    x"3E0524E",
    x"3E0503A",
    x"3E04E26",
    x"3E04C13",
    x"3E04A00",
    x"3E047EE",
    x"3E045DC",
    x"3E043CB",
    x"3E041BA",
    x"3E03FAA",
    x"3E03D9A",
    x"3E03B8B",
    x"3E0397D",
    x"3E0376E",
    x"3E03561",
    x"3E03354",
    x"3E03147",
    x"3E02F3B",
    x"3E02D30",
    x"3E02B25",
    x"3E0291A",
    x"3E02710",
    x"3E02506",
    x"3E022FD",
    x"3E020F5",
    x"3E01EED",
    x"3E01CE5",
    x"3E01ADF",
    x"3E018D8",
    x"3E016D2",
    x"3E014CD",
    x"3E012C8",
    x"3E010C3",
    x"3E00EBF",
    x"3E00CBC",
    x"3E00AB9",
    x"3E008B7",
    x"3E006B5",
    x"3E004B3",
    x"3E002B2",
    x"3E000B2",
    x"3DFFD64",
    x"3DFF965",
    x"3DFF568",
    x"3DFF16B",
    x"3DFED6F",
    x"3DFE974",
    x"3DFE57A",
    x"3DFE181",
    x"3DFDD89",
    x"3DFD992",
    x"3DFD59D",
    x"3DFD1A8",
    x"3DFCDB4",
    x"3DFC9C1",
    x"3DFC5CF",
    x"3DFC1DE",
    x"3DFBDEE",
    x"3DFB9FF",
    x"3DFB611",
    x"3DFB224",
    x"3DFAE38",
    x"3DFAA4D",
    x"3DFA663",
    x"3DFA27A",
    x"3DF9E91",
    x"3DF9AAA",
    x"3DF96C4",
    x"3DF92DF",
    x"3DF8EFB",
    x"3DF8B17",
    x"3DF8735",
    x"3DF8354",
    x"3DF7F73",
    x"3DF7B94",
    x"3DF77B6",
    x"3DF73D8",
    x"3DF6FFC",
    x"3DF6C20",
    x"3DF6846",
    x"3DF646C",
    x"3DF6093",
    x"3DF5CBC",
    x"3DF58E5",
    x"3DF550F",
    x"3DF513B",
    x"3DF4D67",
    x"3DF4994",
    x"3DF45C2",
    x"3DF41F1",
    x"3DF3E21",
    x"3DF3A52",
    x"3DF3684",
    x"3DF32B7",
    x"3DF2EEA",
    x"3DF2B1F",
    x"3DF2755",
    x"3DF238C",
    x"3DF1FC3",
    x"3DF1BFC",
    x"3DF1835",
    x"3DF1470",
    x"3DF10AB",
    x"3DF0CE7",
    x"3DF0924",
    x"3DF0563",
    x"3DF01A2",
    x"3DEFDE2",
    x"3DEFA23",
    x"3DEF665",
    x"3DEF2A8",
    x"3DEEEEB",
    x"3DEEB30",
    x"3DEE776",
    x"3DEE3BC",
    x"3DEE004",
    x"3DEDC4C",
    x"3DED896",
    x"3DED4E0",
    x"3DED12B",
    x"3DECD78",
    x"3DEC9C5",
    x"3DEC613",
    x"3DEC262",
    x"3DEBEB1",
    x"3DEBB02",
    x"3DEB754",
    x"3DEB3A7",
    x"3DEAFFA",
    x"3DEAC4F",
    x"3DEA8A4",
    x"3DEA4FA",
    x"3DEA152",
    x"3DE9DAA",
    x"3DE9A03",
    x"3DE965D",
    x"3DE92B7",
    x"3DE8F13",
    x"3DE8B70",
    x"3DE87CE",
    x"3DE842C",
    x"3DE808B",
    x"3DE7CEC",
    x"3DE794D",
    x"3DE75AF",
    x"3DE7212",
    x"3DE6E76",
    x"3DE6ADB",
    x"3DE6741",
    x"3DE63A7",
    x"3DE600F",
    x"3DE5C77",
    x"3DE58E1",
    x"3DE554B",
    x"3DE51B6",
    x"3DE4E22",
    x"3DE4A8F",
    x"3DE46FD",
    x"3DE436B",
    x"3DE3FDB",
    x"3DE3C4B",
    x"3DE38BD",
    x"3DE352F",
    x"3DE31A2",
    x"3DE2E16",
    x"3DE2A8B",
    x"3DE2701",
    x"3DE2378",
    x"3DE1FEF",
    x"3DE1C68",
    x"3DE18E1",
    x"3DE155B",
    x"3DE11D6",
    x"3DE0E52",
    x"3DE0ACF",
    x"3DE074D",
    x"3DE03CC",
    x"3DE004B",
    x"3DDFCCB",
    x"3DDF94D",
    x"3DDF5CF",
    x"3DDF252",
    x"3DDEED6",
    x"3DDEB5A",
    x"3DDE7E0",
    x"3DDE466",
    x"3DDE0EE",
    x"3DDDD76",
    x"3DDD9FF",
    x"3DDD689",
    x"3DDD314",
    x"3DDCF9F",
    x"3DDCC2C",
    x"3DDC8B9",
    x"3DDC548",
    x"3DDC1D7",
    x"3DDBE67",
    x"3DDBAF7",
    x"3DDB789",
    x"3DDB41C",
    x"3DDB0AF",
    x"3DDAD43",
    x"3DDA9D8",
    x"3DDA66E",
    x"3DDA305",
    x"3DD9F9D",
    x"3DD9C35",
    x"3DD98CF",
    x"3DD9569",
    x"3DD9204",
    x"3DD8EA0",
    x"3DD8B3D",
    x"3DD87DA",
    x"3DD8479",
    x"3DD8118",
    x"3DD7DB8",
    x"3DD7A59",
    x"3DD76FB",
    x"3DD739E",
    x"3DD7041",
    x"3DD6CE6",
    x"3DD698B",
    x"3DD6631",
    x"3DD62D8",
    x"3DD5F7F",
    x"3DD5C28",
    x"3DD58D1",
    x"3DD557C",
    x"3DD5227",
    x"3DD4ED3",
    x"3DD4B7F",
    x"3DD482D",
    x"3DD44DB",
    x"3DD418A",
    x"3DD3E3A",
    x"3DD3AEB",
    x"3DD379D",
    x"3DD344F",
    x"3DD3103",
    x"3DD2DB7",
    x"3DD2A6C",
    x"3DD2722",
    x"3DD23D8",
    x"3DD2090",
    x"3DD1D48",
    x"3DD1A01",
    x"3DD16BB",
    x"3DD1376",
    x"3DD1031",
    x"3DD0CEE",
    x"3DD09AB",
    x"3DD0669",
    x"3DD0328",
    x"3DCFFE7",
    x"3DCFCA8",
    x"3DCF969",
    x"3DCF62B",
    x"3DCF2EE",
    x"3DCEFB2",
    x"3DCEC76",
    x"3DCE93B",
    x"3DCE601",
    x"3DCE2C8",
    x"3DCDF90",
    x"3DCDC59",
    x"3DCD922",
    x"3DCD5EC",
    x"3DCD2B7",
    x"3DCCF83",
    x"3DCCC4F",
    x"3DCC91C",
    x"3DCC5EB",
    x"3DCC2B9",
    x"3DCBF89",
    x"3DCBC5A",
    x"3DCB92B",
    x"3DCB5FD",
    x"3DCB2D0",
    x"3DCAFA4",
    x"3DCAC78",
    x"3DCA94D",
    x"3DCA624",
    x"3DCA2FA",
    x"3DC9FD2",
    x"3DC9CAA",
    x"3DC9984",
    x"3DC965E",
    x"3DC9339",
    x"3DC9014",
    x"3DC8CF0",
    x"3DC89CE",
    x"3DC86AC",
    x"3DC838A",
    x"3DC806A",
    x"3DC7D4A",
    x"3DC7A2B",
    x"3DC770D",
    x"3DC73F0",
    x"3DC70D3",
    x"3DC6DB7",
    x"3DC6A9C",
    x"3DC6782",
    x"3DC6468",
    x"3DC6150",
    x"3DC5E38",
    x"3DC5B21",
    x"3DC580A",
    x"3DC54F5",
    x"3DC51E0",
    x"3DC4ECC",
    x"3DC4BB8",
    x"3DC48A6",
    x"3DC4594",
    x"3DC4283",
    x"3DC3F73",
    x"3DC3C63",
    x"3DC3955",
    x"3DC3647",
    x"3DC3339",
    x"3DC302D",
    x"3DC2D21",
    x"3DC2A16",
    x"3DC270C",
    x"3DC2403",
    x"3DC20FA",
    x"3DC1DF2",
    x"3DC1AEB",
    x"3DC17E5",
    x"3DC14DF",
    x"3DC11DB",
    x"3DC0ED6",
    x"3DC0BD3",
    x"3DC08D1",
    x"3DC05CF",
    x"3DC02CE",
    x"3DBFFCD",
    x"3DBFCCE",
    x"3DBF9CF",
    x"3DBF6D1",
    x"3DBF3D3",
    x"3DBF0D7",
    x"3DBEDDB",
    x"3DBEAE0",
    x"3DBE7E6",
    x"3DBE4EC",
    x"3DBE1F3",
    x"3DBDEFB",
    x"3DBDC04",
    x"3DBD90D",
    x"3DBD617",
    x"3DBD322",
    x"3DBD02E",
    x"3DBCD3A",
    x"3DBCA47",
    x"3DBC755",
    x"3DBC463",
    x"3DBC173",
    x"3DBBE83",
    x"3DBBB93",
    x"3DBB8A5",
    x"3DBB5B7",
    x"3DBB2CA",
    x"3DBAFDE",
    x"3DBACF2",
    x"3DBAA07",
    x"3DBA71D",
    x"3DBA434",
    x"3DBA14B",
    x"3DB9E63",
    x"3DB9B7C",
    x"3DB9895",
    x"3DB95AF",
    x"3DB92CA",
    x"3DB8FE6",
    x"3DB8D02",
    x"3DB8A1F",
    x"3DB873D",
    x"3DB845C",
    x"3DB817B",
    x"3DB7E9B",
    x"3DB7BBC",
    x"3DB78DD",
    x"3DB75FF",
    x"3DB7322",
    x"3DB7046",
    x"3DB6D6A",
    x"3DB6A8F",
    x"3DB67B5",
    x"3DB64DB",
    x"3DB6202",
    x"3DB5F2A",
    x"3DB5C53",
    x"3DB597C",
    x"3DB56A6",
    x"3DB53D1",
    x"3DB50FC",
    x"3DB4E28",
    x"3DB4B55",
    x"3DB4883",
    x"3DB45B1",
    x"3DB42E0",
    x"3DB400F",
    x"3DB3D40",
    x"3DB3A71",
    x"3DB37A3",
    x"3DB34D5",
    x"3DB3208",
    x"3DB2F3C",
    x"3DB2C70",
    x"3DB29A6",
    x"3DB26DC",
    x"3DB2412",
    x"3DB214A",
    x"3DB1E82",
    x"3DB1BBA",
    x"3DB18F4",
    x"3DB162E",
    x"3DB1369",
    x"3DB10A4",
    x"3DB0DE0",
    x"3DB0B1D",
    x"3DB085B",
    x"3DB0599",
    x"3DB02D8",
    x"3DB0018",
    x"3DAFD58",
    x"3DAFA99",
    x"3DAF7DB",
    x"3DAF51D",
    x"3DAF260",
    x"3DAEFA4",
    x"3DAECE8",
    x"3DAEA2D",
    x"3DAE773",
    x"3DAE4BA",
    x"3DAE201",
    x"3DADF49",
    x"3DADC91",
    x"3DAD9DA",
    x"3DAD724",
    x"3DAD46F",
    x"3DAD1BA",
    x"3DACF06",
    x"3DACC53",
    x"3DAC9A0",
    x"3DAC6EE",
    x"3DAC43C",
    x"3DAC18C",
    x"3DABEDC",
    x"3DABC2C",
    x"3DAB97D",
    x"3DAB6CF",
    x"3DAB422",
    x"3DAB175",
    x"3DAAEC9",
    x"3DAAC1E",
    x"3DAA973",
    x"3DAA6C9",
    x"3DAA420",
    x"3DAA177",
    x"3DA9ECF",
    x"3DA9C28",
    x"3DA9981",
    x"3DA96DB",
    x"3DA9436",
    x"3DA9191",
    x"3DA8EED",
    x"3DA8C49",
    x"3DA89A7",
    x"3DA8705",
    x"3DA8463",
    x"3DA81C2",
    x"3DA7F22",
    x"3DA7C83",
    x"3DA79E4",
    x"3DA7746",
    x"3DA74A8",
    x"3DA720C",
    x"3DA6F6F",
    x"3DA6CD4",
    x"3DA6A39",
    x"3DA679F",
    x"3DA6505",
    x"3DA626C",
    x"3DA5FD4",
    x"3DA5D3C",
    x"3DA5AA5",
    x"3DA580F",
    x"3DA5579",
    x"3DA52E4",
    x"3DA5050",
    x"3DA4DBC",
    x"3DA4B29",
    x"3DA4897",
    x"3DA4605",
    x"3DA4373",
    x"3DA40E3",
    x"3DA3E53",
    x"3DA3BC4",
    x"3DA3935",
    x"3DA36A7",
    x"3DA341A",
    x"3DA318D",
    x"3DA2F01",
    x"3DA2C76",
    x"3DA29EB",
    x"3DA2761",
    x"3DA24D7",
    x"3DA224E",
    x"3DA1FC6",
    x"3DA1D3E",
    x"3DA1AB7",
    x"3DA1831",
    x"3DA15AB",
    x"3DA1326",
    x"3DA10A2",
    x"3DA0E1E",
    x"3DA0B9B",
    x"3DA0918",
    x"3DA0696",
    x"3DA0415",
    x"3DA0194",
    x"3D9FF14",
    x"3D9FC95",
    x"3D9FA16",
    x"3D9F797",
    x"3D9F51A",
    x"3D9F29D",
    x"3D9F021",
    x"3D9EDA5",
    x"3D9EB2A",
    x"3D9E8AF",
    x"3D9E635",
    x"3D9E3BC",
    x"3D9E144",
    x"3D9DECC",
    x"3D9DC54",
    x"3D9D9DD",
    x"3D9D767",
    x"3D9D4F2",
    x"3D9D27D",
    x"3D9D008",
    x"3D9CD95",
    x"3D9CB22",
    x"3D9C8AF",
    x"3D9C63D",
    x"3D9C3CC",
    x"3D9C15B",
    x"3D9BEEB",
    x"3D9BC7C",
    x"3D9BA0D",
    x"3D9B79F",
    x"3D9B531",
    x"3D9B2C4",
    x"3D9B058",
    x"3D9ADEC",
    x"3D9AB81",
    x"3D9A916",
    x"3D9A6AC",
    x"3D9A443",
    x"3D9A1DA",
    x"3D99F72",
    x"3D99D0B",
    x"3D99AA4",
    x"3D9983D",
    x"3D995D7",
    x"3D99372",
    x"3D9910E",
    x"3D98EAA",
    x"3D98C46",
    x"3D989E4",
    x"3D98781",
    x"3D98520",
    x"3D982BF",
    x"3D9805F",
    x"3D97DFF",
    x"3D97BA0",
    x"3D97941",
    x"3D976E3",
    x"3D97485",
    x"3D97229",
    x"3D96FCC",
    x"3D96D71",
    x"3D96B16",
    x"3D968BB",
    x"3D96661",
    x"3D96408",
    x"3D961AF",
    x"3D95F57",
    x"3D95D00",
    x"3D95AA9",
    x"3D95852",
    x"3D955FC",
    x"3D953A7",
    x"3D95153",
    x"3D94EFF",
    x"3D94CAB",
    x"3D94A58",
    x"3D94806",
    x"3D945B4",
    x"3D94363",
    x"3D94113",
    x"3D93EC3",
    x"3D93C73",
    x"3D93A24",
    x"3D937D6",
    x"3D93588",
    x"3D9333B",
    x"3D930EF",
    x"3D92EA3",
    x"3D92C58",
    x"3D92A0D",
    x"3D927C2",
    x"3D92579",
    x"3D92330",
    x"3D920E7",
    x"3D91E9F",
    x"3D91C58",
    x"3D91A11",
    x"3D917CB",
    x"3D91585",
    x"3D91340",
    x"3D910FC",
    x"3D90EB8",
    x"3D90C74",
    x"3D90A31",
    x"3D907EF",
    x"3D905AD",
    x"3D9036C",
    x"3D9012C",
    x"3D8FEEC",
    x"3D8FCAC",
    x"3D8FA6D",
    x"3D8F82F",
    x"3D8F5F1",
    x"3D8F3B4",
    x"3D8F177",
    x"3D8EF3B",
    x"3D8ED00",
    x"3D8EAC5",
    x"3D8E88A",
    x"3D8E651",
    x"3D8E417",
    x"3D8E1DF",
    x"3D8DFA6",
    x"3D8DD6F",
    x"3D8DB38",
    x"3D8D901",
    x"3D8D6CB",
    x"3D8D496",
    x"3D8D261",
    x"3D8D02C",
    x"3D8CDF9",
    x"3D8CBC6",
    x"3D8C993",
    x"3D8C761",
    x"3D8C52F",
    x"3D8C2FE",
    x"3D8C0CE",
    x"3D8BE9E",
    x"3D8BC6E",
    x"3D8BA40",
    x"3D8B811",
    x"3D8B5E3",
    x"3D8B3B6",
    x"3D8B18A",
    x"3D8AF5D",
    x"3D8AD32",
    x"3D8AB07",
    x"3D8A8DC",
    x"3D8A6B2",
    x"3D8A489",
    x"3D8A260",
    x"3D8A038",
    x"3D89E10",
    x"3D89BE9",
    x"3D899C2",
    x"3D8979C",
    x"3D89576",
    x"3D89351",
    x"3D8912D",
    x"3D88F09",
    x"3D88CE5",
    x"3D88AC2",
    x"3D888A0",
    x"3D8867E",
    x"3D8845D",
    x"3D8823C",
    x"3D8801B",
    x"3D87DFC",
    x"3D87BDC",
    x"3D879BE",
    x"3D877A0",
    x"3D87582",
    x"3D87365",
    x"3D87148",
    x"3D86F2C",
    x"3D86D11",
    x"3D86AF6",
    x"3D868DB",
    x"3D866C1",
    x"3D864A8",
    x"3D8628F",
    x"3D86076",
    x"3D85E5F",
    x"3D85C47",
    x"3D85A30",
    x"3D8581A",
    x"3D85604",
    x"3D853EF",
    x"3D851DA",
    x"3D84FC6",
    x"3D84DB3",
    x"3D84B9F",
    x"3D8498D",
    x"3D8477B",
    x"3D84569",
    x"3D84358",
    x"3D84147",
    x"3D83F37",
    x"3D83D28",
    x"3D83B19",
    x"3D8390A",
    x"3D836FC",
    x"3D834EF",
    x"3D832E2",
    x"3D830D5",
    x"3D82EC9",
    x"3D82CBE",
    x"3D82AB3",
    x"3D828A9",
    x"3D8269F",
    x"3D82495",
    x"3D8228C",
    x"3D82084",
    x"3D81E7C",
    x"3D81C75",
    x"3D81A6E",
    x"3D81867",
    x"3D81662",
    x"3D8145C",
    x"3D81257",
    x"3D81053",
    x"3D80E4F",
    x"3D80C4C",
    x"3D80A49",
    x"3D80847",
    x"3D80645",
    x"3D80444",
    x"3D80243",
    x"3D80043",
    x"3D7FC86",
    x"3D7F887",
    x"3D7F48A",
    x"3D7F08D",
    x"3D7EC91",
    x"3D7E897",
    x"3D7E49D",
    x"3D7E0A4",
    x"3D7DCAD",
    x"3D7D8B6",
    x"3D7D4C0",
    x"3D7D0CC",
    x"3D7CCD8",
    x"3D7C8E5",
    x"3D7C4F4",
    x"3D7C103",
    x"3D7BD13",
    x"3D7B924",
    x"3D7B536",
    x"3D7B14A",
    x"3D7AD5E",
    x"3D7A973",
    x"3D7A589",
    x"3D7A1A0",
    x"3D79DB8",
    x"3D799D1",
    x"3D795EB",
    x"3D79206",
    x"3D78E22",
    x"3D78A3F",
    x"3D7865D",
    x"3D7827C",
    x"3D77E9C",
    x"3D77ABD",
    x"3D776DF",
    x"3D77301",
    x"3D76F25",
    x"3D76B4A",
    x"3D7676F",
    x"3D76396",
    x"3D75FBE",
    x"3D75BE6",
    x"3D75810",
    x"3D7543A",
    x"3D75066",
    x"3D74C92",
    x"3D748BF",
    x"3D744EE",
    x"3D7411D",
    x"3D73D4D",
    x"3D7397E",
    x"3D735B0",
    x"3D731E3",
    x"3D72E17",
    x"3D72A4C",
    x"3D72682",
    x"3D722B9",
    x"3D71EF1",
    x"3D71B2A",
    x"3D71763",
    x"3D7139E",
    x"3D70FD9",
    x"3D70C16",
    x"3D70853",
    x"3D70492",
    x"3D700D1",
    x"3D6FD11",
    x"3D6F953",
    x"3D6F595",
    x"3D6F1D8",
    x"3D6EE1C",
    x"3D6EA61",
    x"3D6E6A7",
    x"3D6E2ED",
    x"3D6DF35",
    x"3D6DB7E",
    x"3D6D7C7",
    x"3D6D412",
    x"3D6D05D",
    x"3D6CCAA",
    x"3D6C8F7",
    x"3D6C545",
    x"3D6C194",
    x"3D6BDE4",
    x"3D6BA35",
    x"3D6B687",
    x"3D6B2DA",
    x"3D6AF2E",
    x"3D6AB83",
    x"3D6A7D8",
    x"3D6A42F",
    x"3D6A086",
    x"3D69CDE",
    x"3D69938",
    x"3D69592",
    x"3D691ED",
    x"3D68E49",
    x"3D68AA6",
    x"3D68704",
    x"3D68362",
    x"3D67FC2",
    x"3D67C22",
    x"3D67884",
    x"3D674E6",
    x"3D67149",
    x"3D66DAD",
    x"3D66A12",
    x"3D66678",
    x"3D662DF",
    x"3D65F47",
    x"3D65BB0",
    x"3D65819",
    x"3D65484",
    x"3D650EF",
    x"3D64D5B",
    x"3D649C8",
    x"3D64636",
    x"3D642A5",
    x"3D63F15",
    x"3D63B86",
    x"3D637F7",
    x"3D6346A",
    x"3D630DD",
    x"3D62D51",
    x"3D629C6",
    x"3D6263C",
    x"3D622B3",
    x"3D61F2B",
    x"3D61BA4",
    x"3D6181D",
    x"3D61497",
    x"3D61113",
    x"3D60D8F",
    x"3D60A0C",
    x"3D6068A",
    x"3D60309",
    x"3D5FF88",
    x"3D5FC09",
    x"3D5F88A",
    x"3D5F50D",
    x"3D5F190",
    x"3D5EE14",
    x"3D5EA99",
    x"3D5E71F",
    x"3D5E3A5",
    x"3D5E02D",
    x"3D5DCB5",
    x"3D5D93E",
    x"3D5D5C9",
    x"3D5D253",
    x"3D5CEDF",
    x"3D5CB6C",
    x"3D5C7FA",
    x"3D5C488",
    x"3D5C117",
    x"3D5BDA8",
    x"3D5BA39",
    x"3D5B6CA",
    x"3D5B35D",
    x"3D5AFF1",
    x"3D5AC85",
    x"3D5A91A",
    x"3D5A5B1",
    x"3D5A248",
    x"3D59EDF",
    x"3D59B78",
    x"3D59812",
    x"3D594AC",
    x"3D59147",
    x"3D58DE4",
    x"3D58A80",
    x"3D5871E",
    x"3D583BD",
    x"3D5805C",
    x"3D57CFD",
    x"3D5799E",
    x"3D57640",
    x"3D572E3",
    x"3D56F86",
    x"3D56C2B",
    x"3D568D0",
    x"3D56577",
    x"3D5621E",
    x"3D55EC6",
    x"3D55B6E",
    x"3D55818",
    x"3D554C2",
    x"3D5516D",
    x"3D54E19",
    x"3D54AC6",
    x"3D54774",
    x"3D54423",
    x"3D540D2",
    x"3D53D82",
    x"3D53A33",
    x"3D536E5",
    x"3D53398",
    x"3D5304B",
    x"3D52D00",
    x"3D529B5",
    x"3D5266B",
    x"3D52322",
    x"3D51FD9",
    x"3D51C92",
    x"3D5194B",
    x"3D51605",
    x"3D512C0",
    x"3D50F7C",
    x"3D50C38",
    x"3D508F6",
    x"3D505B4",
    x"3D50273",
    x"3D4FF33",
    x"3D4FBF3",
    x"3D4F8B5",
    x"3D4F577",
    x"3D4F23A",
    x"3D4EEFE",
    x"3D4EBC2",
    x"3D4E888",
    x"3D4E54E",
    x"3D4E215",
    x"3D4DEDD",
    x"3D4DBA6",
    x"3D4D86F",
    x"3D4D539",
    x"3D4D205",
    x"3D4CED0",
    x"3D4CB9D",
    x"3D4C86B",
    x"3D4C539",
    x"3D4C208",
    x"3D4BED8",
    x"3D4BBA9",
    x"3D4B87A",
    x"3D4B54C",
    x"3D4B21F",
    x"3D4AEF3",
    x"3D4ABC8",
    x"3D4A89D",
    x"3D4A574",
    x"3D4A24B",
    x"3D49F23",
    x"3D49BFB",
    x"3D498D5",
    x"3D495AF",
    x"3D4928A",
    x"3D48F65",
    x"3D48C42",
    x"3D4891F",
    x"3D485FD",
    x"3D482DC",
    x"3D47FBC",
    x"3D47C9C",
    x"3D4797E",
    x"3D47660",
    x"3D47342",
    x"3D47026",
    x"3D46D0A",
    x"3D469F0",
    x"3D466D5",
    x"3D463BC",
    x"3D460A4",
    x"3D45D8C",
    x"3D45A75",
    x"3D4575F",
    x"3D45449",
    x"3D45134",
    x"3D44E21",
    x"3D44B0D",
    x"3D447FB",
    x"3D444E9",
    x"3D441D9",
    x"3D43EC8",
    x"3D43BB9",
    x"3D438AB",
    x"3D4359D",
    x"3D43290",
    x"3D42F84",
    x"3D42C78",
    x"3D4296D",
    x"3D42663",
    x"3D4235A",
    x"3D42052",
    x"3D41D4A",
    x"3D41A43",
    x"3D4173D",
    x"3D41437",
    x"3D41133",
    x"3D40E2F",
    x"3D40B2C",
    x"3D40829",
    x"3D40528",
    x"3D40227",
    x"3D3FF26",
    x"3D3FC27",
    x"3D3F928",
    x"3D3F62A",
    x"3D3F32D",
    x"3D3F031",
    x"3D3ED35",
    x"3D3EA3A",
    x"3D3E740",
    x"3D3E447",
    x"3D3E14E",
    x"3D3DE56",
    x"3D3DB5F",
    x"3D3D868",
    x"3D3D573",
    x"3D3D27E",
    x"3D3CF89",
    x"3D3CC96",
    x"3D3C9A3",
    x"3D3C6B1",
    x"3D3C3C0",
    x"3D3C0CF",
    x"3D3BDDF",
    x"3D3BAF0",
    x"3D3B802",
    x"3D3B514",
    x"3D3B227",
    x"3D3AF3B",
    x"3D3AC50",
    x"3D3A965",
    x"3D3A67B",
    x"3D3A392",
    x"3D3A0A9",
    x"3D39DC1",
    x"3D39ADA",
    x"3D397F4",
    x"3D3950E",
    x"3D39229",
    x"3D38F45",
    x"3D38C62",
    x"3D3897F",
    x"3D3869D",
    x"3D383BC",
    x"3D380DB",
    x"3D37DFB",
    x"3D37B1C",
    x"3D3783E",
    x"3D37560",
    x"3D37283",
    x"3D36FA7",
    x"3D36CCB",
    x"3D369F0",
    x"3D36716",
    x"3D3643D",
    x"3D36164",
    x"3D35E8C",
    x"3D35BB5",
    x"3D358DE",
    x"3D35608",
    x"3D35333",
    x"3D3505F",
    x"3D34D8B",
    x"3D34AB8",
    x"3D347E6",
    x"3D34514",
    x"3D34243",
    x"3D33F73",
    x"3D33CA3",
    x"3D339D5",
    x"3D33707",
    x"3D33439",
    x"3D3316C",
    x"3D32EA0",
    x"3D32BD5",
    x"3D3290A",
    x"3D32641",
    x"3D32377",
    x"3D320AF",
    x"3D31DE7",
    x"3D31B20",
    x"3D31859",
    x"3D31594",
    x"3D312CF",
    x"3D3100A",
    x"3D30D47",
    x"3D30A84",
    x"3D307C1",
    x"3D30500",
    x"3D3023F",
    x"3D2FF7F",
    x"3D2FCBF",
    x"3D2FA00",
    x"3D2F742",
    x"3D2F485",
    x"3D2F1C8",
    x"3D2EF0C",
    x"3D2EC50",
    x"3D2E996",
    x"3D2E6DC",
    x"3D2E422",
    x"3D2E169",
    x"3D2DEB1",
    x"3D2DBFA",
    x"3D2D943",
    x"3D2D68E",
    x"3D2D3D8",
    x"3D2D124",
    x"3D2CE70",
    x"3D2CBBC",
    x"3D2C90A",
    x"3D2C658",
    x"3D2C3A7",
    x"3D2C0F6",
    x"3D2BE46",
    x"3D2BB97",
    x"3D2B8E8",
    x"3D2B63A",
    x"3D2B38D",
    x"3D2B0E1",
    x"3D2AE35",
    x"3D2AB8A",
    x"3D2A8DF",
    x"3D2A635",
    x"3D2A38C",
    x"3D2A0E3",
    x"3D29E3B",
    x"3D29B94",
    x"3D298EE",
    x"3D29648",
    x"3D293A3",
    x"3D290FE",
    x"3D28E5A",
    x"3D28BB7",
    x"3D28914",
    x"3D28672",
    x"3D283D1",
    x"3D28130",
    x"3D27E90",
    x"3D27BF1",
    x"3D27952",
    x"3D276B4",
    x"3D27417",
    x"3D2717A",
    x"3D26EDE",
    x"3D26C43",
    x"3D269A8",
    x"3D2670E",
    x"3D26475",
    x"3D261DC",
    x"3D25F44",
    x"3D25CAC",
    x"3D25A15",
    x"3D2577F",
    x"3D254EA",
    x"3D25255",
    x"3D24FC0",
    x"3D24D2D",
    x"3D24A9A",
    x"3D24808",
    x"3D24576",
    x"3D242E5",
    x"3D24054",
    x"3D23DC5",
    x"3D23B35",
    x"3D238A7",
    x"3D23619",
    x"3D2338C",
    x"3D230FF",
    x"3D22E73",
    x"3D22BE8",
    x"3D2295E",
    x"3D226D3",
    x"3D2244A",
    x"3D221C1",
    x"3D21F39",
    x"3D21CB2",
    x"3D21A2B",
    x"3D217A5",
    x"3D2151F",
    x"3D2129A",
    x"3D21016",
    x"3D20D92",
    x"3D20B0F",
    x"3D2088D",
    x"3D2060B",
    x"3D20389",
    x"3D20109",
    x"3D1FE89",
    x"3D1FC0A",
    x"3D1F98B",
    x"3D1F70D",
    x"3D1F48F",
    x"3D1F213",
    x"3D1EF96",
    x"3D1ED1B",
    x"3D1EAA0",
    x"3D1E825",
    x"3D1E5AC",
    x"3D1E333",
    x"3D1E0BA",
    x"3D1DE42",
    x"3D1DBCB",
    x"3D1D954",
    x"3D1D6DE",
    x"3D1D469",
    x"3D1D1F4",
    x"3D1CF80",
    x"3D1CD0C",
    x"3D1CA99",
    x"3D1C827",
    x"3D1C5B5",
    x"3D1C344",
    x"3D1C0D4",
    x"3D1BE64",
    x"3D1BBF5",
    x"3D1B986",
    x"3D1B718",
    x"3D1B4AA",
    x"3D1B23D",
    x"3D1AFD1",
    x"3D1AD66",
    x"3D1AAFA",
    x"3D1A890",
    x"3D1A626",
    x"3D1A3BD",
    x"3D1A154",
    x"3D19EEC",
    x"3D19C85",
    x"3D19A1E",
    x"3D197B8",
    x"3D19552",
    x"3D192ED",
    x"3D19089",
    x"3D18E25",
    x"3D18BC2",
    x"3D1895F",
    x"3D186FD",
    x"3D1849C",
    x"3D1823B",
    x"3D17FDA",
    x"3D17D7B",
    x"3D17B1C",
    x"3D178BD",
    x"3D1765F",
    x"3D17402",
    x"3D171A5",
    x"3D16F49",
    x"3D16CEE",
    x"3D16A93",
    x"3D16838",
    x"3D165DF",
    x"3D16385",
    x"3D1612D",
    x"3D15ED5",
    x"3D15C7D",
    x"3D15A27",
    x"3D157D0",
    x"3D1557B",
    x"3D15326",
    x"3D150D1",
    x"3D14E7D",
    x"3D14C2A",
    x"3D149D7",
    x"3D14785",
    x"3D14533",
    x"3D142E2",
    x"3D14092",
    x"3D13E42",
    x"3D13BF3",
    x"3D139A4",
    x"3D13756",
    x"3D13508",
    x"3D132BB",
    x"3D1306F",
    x"3D12E23",
    x"3D12BD8",
    x"3D1298D",
    x"3D12743",
    x"3D124FA",
    x"3D122B1",
    x"3D12068",
    x"3D11E20",
    x"3D11BD9",
    x"3D11993",
    x"3D1174C",
    x"3D11507",
    x"3D112C2",
    x"3D1107E",
    x"3D10E3A",
    x"3D10BF6",
    x"3D109B4",
    x"3D10772",
    x"3D10530",
    x"3D102EF",
    x"3D100AF",
    x"3D0FE6F",
    x"3D0FC2F",
    x"3D0F9F1",
    x"3D0F7B2",
    x"3D0F575",
    x"3D0F338",
    x"3D0F0FB",
    x"3D0EEBF",
    x"3D0EC84",
    x"3D0EA49",
    x"3D0E80F",
    x"3D0E5D5",
    x"3D0E39C",
    x"3D0E163",
    x"3D0DF2B",
    x"3D0DCF3",
    x"3D0DABC",
    x"3D0D886",
    x"3D0D650",
    x"3D0D41B",
    x"3D0D1E6",
    x"3D0CFB2",
    x"3D0CD7E",
    x"3D0CB4B",
    x"3D0C919",
    x"3D0C6E7",
    x"3D0C4B5",
    x"3D0C284",
    x"3D0C054",
    x"3D0BE24",
    x"3D0BBF5",
    x"3D0B9C6",
    x"3D0B798",
    x"3D0B56A",
    x"3D0B33D",
    x"3D0B111",
    x"3D0AEE5",
    x"3D0ACB9",
    x"3D0AA8E",
    x"3D0A864",
    x"3D0A63A",
    x"3D0A411",
    x"3D0A1E8",
    x"3D09FC0",
    x"3D09D98",
    x"3D09B71",
    x"3D0994B",
    x"3D09724",
    x"3D094FF",
    x"3D092DA",
    x"3D090B6",
    x"3D08E92",
    x"3D08C6E",
    x"3D08A4B",
    x"3D08829",
    x"3D08607",
    x"3D083E6",
    x"3D081C5",
    x"3D07FA5",
    x"3D07D86",
    x"3D07B66",
    x"3D07948",
    x"3D0772A",
    x"3D0750C",
    x"3D072EF",
    x"3D070D3",
    x"3D06EB7",
    x"3D06C9B",
    x"3D06A81",
    x"3D06866",
    x"3D0664C",
    x"3D06433",
    x"3D0621A",
    x"3D06002",
    x"3D05DEA",
    x"3D05BD3",
    x"3D059BC",
    x"3D057A6",
    x"3D05591",
    x"3D0537B",
    x"3D05167",
    x"3D04F53",
    x"3D04D3F",
    x"3D04B2C",
    x"3D0491A",
    x"3D04708",
    x"3D044F6",
    x"3D042E5",
    x"3D040D5",
    x"3D03EC5",
    x"3D03CB5",
    x"3D03AA6",
    x"3D03898",
    x"3D0368A",
    x"3D0347D",
    x"3D03270",
    x"3D03063",
    x"3D02E58",
    x"3D02C4C",
    x"3D02A41",
    x"3D02837",
    x"3D0262D",
    x"3D02424",
    x"3D0221B",
    x"3D02013",
    x"3D01E0B",
    x"3D01C04",
    x"3D019FD",
    x"3D017F7",
    x"3D015F1",
    x"3D013EC",
    x"3D011E7",
    x"3D00FE3",
    x"3D00DDF",
    x"3D00BDC",
    x"3D009D9",
    x"3D007D7",
    x"3D005D5",
    x"3D003D4",
    x"3D001D3",
    x"3CFFFA7",
    x"3CFFBA8",
    x"3CFF7A9",
    x"3CFF3AC",
    x"3CFEFAF",
    x"3CFEBB4",
    x"3CFE7BA",
    x"3CFE3C0",
    x"3CFDFC8",
    x"3CFDBD0",
    x"3CFD7DA",
    x"3CFD3E4",
    x"3CFCFF0",
    x"3CFCBFC",
    x"3CFC80A",
    x"3CFC418",
    x"3CFC028",
    x"3CFBC38",
    x"3CFB84A",
    x"3CFB45C",
    x"3CFB06F",
    x"3CFAC84",
    x"3CFA899",
    x"3CFA4B0",
    x"3CFA0C7",
    x"3CF9CDF",
    x"3CF98F8",
    x"3CF9513",
    x"3CF912E",
    x"3CF8D4A",
    x"3CF8967",
    x"3CF8585",
    x"3CF81A4",
    x"3CF7DC5",
    x"3CF79E6",
    x"3CF7608",
    x"3CF722B",
    x"3CF6E4E",
    x"3CF6A73",
    x"3CF6699",
    x"3CF62C0",
    x"3CF5EE8",
    x"3CF5B11",
    x"3CF573A",
    x"3CF5365",
    x"3CF4F91",
    x"3CF4BBD",
    x"3CF47EB",
    x"3CF4419",
    x"3CF4049",
    x"3CF3C79",
    x"3CF38AB",
    x"3CF34DD",
    x"3CF3110",
    x"3CF2D44",
    x"3CF2979",
    x"3CF25B0",
    x"3CF21E7",
    x"3CF1E1F",
    x"3CF1A58",
    x"3CF1691",
    x"3CF12CC",
    x"3CF0F08",
    x"3CF0B45",
    x"3CF0782",
    x"3CF03C1",
    x"3CF0001",
    x"3CEFC41",
    x"3CEF882",
    x"3CEF4C5",
    x"3CEF108",
    x"3CEED4C",
    x"3CEE991",
    x"3CEE5D7",
    x"3CEE21E",
    x"3CEDE66",
    x"3CEDAAF",
    x"3CED6F9",
    x"3CED344",
    x"3CECF8F",
    x"3CECBDC",
    x"3CEC829",
    x"3CEC478",
    x"3CEC0C7",
    x"3CEBD17",
    x"3CEB969",
    x"3CEB5BB",
    x"3CEB20E",
    x"3CEAE62",
    x"3CEAAB7",
    x"3CEA70C",
    x"3CEA363",
    x"3CE9FBB",
    x"3CE9C13",
    x"3CE986D",
    x"3CE94C7",
    x"3CE9122",
    x"3CE8D7E",
    x"3CE89DC",
    x"3CE8639",
    x"3CE8298",
    x"3CE7EF8",
    x"3CE7B59",
    x"3CE77BB",
    x"3CE741D",
    x"3CE7080",
    x"3CE6CE5",
    x"3CE694A",
    x"3CE65B0",
    x"3CE6217",
    x"3CE5E7F",
    x"3CE5AE8",
    x"3CE5752",
    x"3CE53BC",
    x"3CE5028",
    x"3CE4C94",
    x"3CE4901",
    x"3CE4570",
    x"3CE41DF",
    x"3CE3E4F",
    x"3CE3AC0",
    x"3CE3731",
    x"3CE33A4",
    x"3CE3018",
    x"3CE2C8C",
    x"3CE2901",
    x"3CE2577",
    x"3CE21EF",
    x"3CE1E66",
    x"3CE1ADF",
    x"3CE1759",
    x"3CE13D4",
    x"3CE104F",
    x"3CE0CCC",
    x"3CE0949",
    x"3CE05C7",
    x"3CE0246",
    x"3CDFEC6",
    x"3CDFB46",
    x"3CDF7C8",
    x"3CDF44B",
    x"3CDF0CE",
    x"3CDED52",
    x"3CDE9D7",
    x"3CDE65D",
    x"3CDE2E4",
    x"3CDDF6C",
    x"3CDDBF4",
    x"3CDD87E",
    x"3CDD508",
    x"3CDD193",
    x"3CDCE1F",
    x"3CDCAAC",
    x"3CDC73A",
    x"3CDC3C9",
    x"3CDC058",
    x"3CDBCE8",
    x"3CDB97A",
    x"3CDB60C",
    x"3CDB29F",
    x"3CDAF32",
    x"3CDABC7",
    x"3CDA85D",
    x"3CDA4F3",
    x"3CDA18A",
    x"3CD9E22",
    x"3CD9ABB",
    x"3CD9755",
    x"3CD93EF",
    x"3CD908B",
    x"3CD8D27",
    x"3CD89C4",
    x"3CD8662",
    x"3CD8301",
    x"3CD7FA1",
    x"3CD7C41",
    x"3CD78E3",
    x"3CD7585",
    x"3CD7228",
    x"3CD6ECC",
    x"3CD6B70",
    x"3CD6816",
    x"3CD64BC",
    x"3CD6164",
    x"3CD5E0C",
    x"3CD5AB5",
    x"3CD575E",
    x"3CD5409",
    x"3CD50B4",
    x"3CD4D60",
    x"3CD4A0E",
    x"3CD46BB",
    x"3CD436A",
    x"3CD401A",
    x"3CD3CCA",
    x"3CD397B",
    x"3CD362D",
    x"3CD32E0",
    x"3CD2F94",
    x"3CD2C48",
    x"3CD28FE",
    x"3CD25B4",
    x"3CD226B",
    x"3CD1F23",
    x"3CD1BDB",
    x"3CD1895",
    x"3CD154F",
    x"3CD120A",
    x"3CD0EC6",
    x"3CD0B83",
    x"3CD0840",
    x"3CD04FF",
    x"3CD01BE",
    x"3CCFE7E",
    x"3CCFB3F",
    x"3CCF800",
    x"3CCF4C3",
    x"3CCF186",
    x"3CCEE4A",
    x"3CCEB0F",
    x"3CCE7D4",
    x"3CCE49B",
    x"3CCE162",
    x"3CCDE2A",
    x"3CCDAF3",
    x"3CCD7BD",
    x"3CCD487",
    x"3CCD152",
    x"3CCCE1E",
    x"3CCCAEB",
    x"3CCC7B9",
    x"3CCC487",
    x"3CCC157",
    x"3CCBE27",
    x"3CCBAF8",
    x"3CCB7C9",
    x"3CCB49C",
    x"3CCB16F",
    x"3CCAE43",
    x"3CCAB18",
    x"3CCA7ED",
    x"3CCA4C4",
    x"3CCA19B",
    x"3CC9E73",
    x"3CC9B4C",
    x"3CC9825",
    x"3CC9500",
    x"3CC91DB",
    x"3CC8EB7",
    x"3CC8B94",
    x"3CC8871",
    x"3CC854F",
    x"3CC822E",
    x"3CC7F0E",
    x"3CC7BEF",
    x"3CC78D0",
    x"3CC75B2",
    x"3CC7295",
    x"3CC6F79",
    x"3CC6C5E",
    x"3CC6943",
    x"3CC6629",
    x"3CC6310",
    x"3CC5FF7",
    x"3CC5CE0",
    x"3CC59C9",
    x"3CC56B3",
    x"3CC539E",
    x"3CC5089",
    x"3CC4D75",
    x"3CC4A62",
    x"3CC4750",
    x"3CC443F",
    x"3CC412E",
    x"3CC3E1E",
    x"3CC3B0F",
    x"3CC3801",
    x"3CC34F3",
    x"3CC31E6",
    x"3CC2EDA",
    x"3CC2BCF",
    x"3CC28C4",
    x"3CC25BA",
    x"3CC22B1",
    x"3CC1FA9",
    x"3CC1CA1",
    x"3CC199B",
    x"3CC1695",
    x"3CC138F",
    x"3CC108B",
    x"3CC0D87",
    x"3CC0A84",
    x"3CC0782",
    x"3CC0480",
    x"3CC0180",
    x"3CBFE80",
    x"3CBFB80",
    x"3CBF882",
    x"3CBF584",
    x"3CBF287",
    x"3CBEF8B",
    x"3CBEC8F",
    x"3CBE995",
    x"3CBE69B",
    x"3CBE3A1",
    x"3CBE0A9",
    x"3CBDDB1",
    x"3CBDABA",
    x"3CBD7C4",
    x"3CBD4CE",
    x"3CBD1D9",
    x"3CBCEE5",
    x"3CBCBF2",
    x"3CBC8FF",
    x"3CBC60D",
    x"3CBC31C",
    x"3CBC02C",
    x"3CBBD3C",
    x"3CBBA4D",
    x"3CBB75F",
    x"3CBB471",
    x"3CBB185",
    x"3CBAE99",
    x"3CBABAD",
    x"3CBA8C3",
    x"3CBA5D9",
    x"3CBA2F0",
    x"3CBA007",
    x"3CB9D20",
    x"3CB9A39",
    x"3CB9753",
    x"3CB946D",
    x"3CB9189",
    x"3CB8EA4",
    x"3CB8BC1",
    x"3CB88DF",
    x"3CB85FD",
    x"3CB831C",
    x"3CB803B",
    x"3CB7D5B",
    x"3CB7A7D",
    x"3CB779E",
    x"3CB74C1",
    x"3CB71E4",
    x"3CB6F08",
    x"3CB6C2C",
    x"3CB6952",
    x"3CB6678",
    x"3CB639E",
    x"3CB60C6",
    x"3CB5DEE",
    x"3CB5B17",
    x"3CB5840",
    x"3CB556B",
    x"3CB5296",
    x"3CB4FC1",
    x"3CB4CEE",
    x"3CB4A1B",
    x"3CB4749",
    x"3CB4477",
    x"3CB41A7",
    x"3CB3ED7",
    x"3CB3C07",
    x"3CB3939",
    x"3CB366B",
    x"3CB339D",
    x"3CB30D1",
    x"3CB2E05",
    x"3CB2B3A",
    x"3CB286F",
    x"3CB25A6",
    x"3CB22DC",
    x"3CB2014",
    x"3CB1D4C",
    x"3CB1A85",
    x"3CB17BF",
    x"3CB14FA",
    x"3CB1235",
    x"3CB0F70",
    x"3CB0CAD",
    x"3CB09EA",
    x"3CB0728",
    x"3CB0467",
    x"3CB01A6",
    x"3CAFEE6",
    x"3CAFC26",
    x"3CAF968",
    x"3CAF6AA",
    x"3CAF3EC",
    x"3CAF130",
    x"3CAEE74",
    x"3CAEBB8",
    x"3CAE8FE",
    x"3CAE644",
    x"3CAE38B",
    x"3CAE0D2",
    x"3CADE1A",
    x"3CADB63",
    x"3CAD8AD",
    x"3CAD5F7",
    x"3CAD342",
    x"3CAD08D",
    x"3CACDD9",
    x"3CACB26",
    x"3CAC874",
    x"3CAC5C2",
    x"3CAC311",
    x"3CAC060",
    x"3CABDB1",
    x"3CABB02",
    x"3CAB853",
    x"3CAB5A5",
    x"3CAB2F8",
    x"3CAB04C",
    x"3CAADA0",
    x"3CAAAF5",
    x"3CAA84B",
    x"3CAA5A1",
    x"3CAA2F8",
    x"3CAA050",
    x"3CA9DA8",
    x"3CA9B01",
    x"3CA985A",
    x"3CA95B5",
    x"3CA930F",
    x"3CA906B",
    x"3CA8DC7",
    x"3CA8B24",
    x"3CA8882",
    x"3CA85E0",
    x"3CA833F",
    x"3CA809E",
    x"3CA7DFE",
    x"3CA7B5F",
    x"3CA78C1",
    x"3CA7623",
    x"3CA7386",
    x"3CA70E9",
    x"3CA6E4D",
    x"3CA6BB2",
    x"3CA6917",
    x"3CA667D",
    x"3CA63E4",
    x"3CA614B",
    x"3CA5EB3",
    x"3CA5C1C",
    x"3CA5985",
    x"3CA56EF",
    x"3CA545A",
    x"3CA51C5",
    x"3CA4F31",
    x"3CA4C9E",
    x"3CA4A0B",
    x"3CA4779",
    x"3CA44E7",
    x"3CA4256",
    x"3CA3FC6",
    x"3CA3D36",
    x"3CA3AA7",
    x"3CA3819",
    x"3CA358B",
    x"3CA32FE",
    x"3CA3072",
    x"3CA2DE6",
    x"3CA2B5B",
    x"3CA28D0",
    x"3CA2646",
    x"3CA23BD",
    x"3CA2134",
    x"3CA1EAC",
    x"3CA1C25",
    x"3CA199E",
    x"3CA1718",
    x"3CA1493",
    x"3CA120E",
    x"3CA0F8A",
    x"3CA0D06",
    x"3CA0A83",
    x"3CA0801",
    x"3CA057F",
    x"3CA02FE",
    x"3CA007E",
    x"3C9FDFE",
    x"3C9FB7F",
    x"3C9F900",
    x"3C9F682",
    x"3C9F405",
    x"3C9F188",
    x"3C9EF0C",
    x"3C9EC91",
    x"3C9EA16",
    x"3C9E79C",
    x"3C9E522",
    x"3C9E2A9",
    x"3C9E031",
    x"3C9DDB9",
    x"3C9DB42",
    x"3C9D8CB",
    x"3C9D656",
    x"3C9D3E0",
    x"3C9D16C",
    x"3C9CEF8",
    x"3C9CC84",
    x"3C9CA11",
    x"3C9C79F",
    x"3C9C52D",
    x"3C9C2BC",
    x"3C9C04C",
    x"3C9BDDC",
    x"3C9BB6D",
    x"3C9B8FF",
    x"3C9B691",
    x"3C9B423",
    x"3C9B1B7",
    x"3C9AF4A",
    x"3C9ACDF",
    x"3C9AA74",
    x"3C9A80A",
    x"3C9A5A0",
    x"3C9A337",
    x"3C9A0CE",
    x"3C99E67",
    x"3C99BFF",
    x"3C99999",
    x"3C99732",
    x"3C994CD",
    x"3C99268",
    x"3C99004",
    x"3C98DA0",
    x"3C98B3D",
    x"3C988DA",
    x"3C98678",
    x"3C98417",
    x"3C981B6",
    x"3C97F56",
    x"3C97CF7",
    x"3C97A98",
    x"3C97839",
    x"3C975DC",
    x"3C9737F",
    x"3C97122",
    x"3C96EC6",
    x"3C96C6B",
    x"3C96A10",
    x"3C967B6",
    x"3C9655C",
    x"3C96303",
    x"3C960AA",
    x"3C95E53",
    x"3C95BFB",
    x"3C959A5",
    x"3C9574E",
    x"3C954F9",
    x"3C952A4",
    x"3C95050",
    x"3C94DFC",
    x"3C94BA9",
    x"3C94956",
    x"3C94704",
    x"3C944B2",
    x"3C94262",
    x"3C94011",
    x"3C93DC2",
    x"3C93B72",
    x"3C93924",
    x"3C936D6",
    x"3C93488",
    x"3C9323C",
    x"3C92FEF",
    x"3C92DA4",
    x"3C92B58",
    x"3C9290E",
    x"3C926C4",
    x"3C9247A",
    x"3C92232",
    x"3C91FE9",
    x"3C91DA2",
    x"3C91B5B",
    x"3C91914",
    x"3C916CE",
    x"3C91489",
    x"3C91244",
    x"3C90FFF",
    x"3C90DBC",
    x"3C90B79",
    x"3C90936",
    x"3C906F4",
    x"3C904B3",
    x"3C90272",
    x"3C90031",
    x"3C8FDF2",
    x"3C8FBB2",
    x"3C8F974",
    x"3C8F736",
    x"3C8F4F8",
    x"3C8F2BB",
    x"3C8F07F",
    x"3C8EE43",
    x"3C8EC08",
    x"3C8E9CD",
    x"3C8E793",
    x"3C8E559",
    x"3C8E320",
    x"3C8E0E8",
    x"3C8DEB0",
    x"3C8DC78",
    x"3C8DA41",
    x"3C8D80B",
    x"3C8D5D5",
    x"3C8D3A0",
    x"3C8D16C",
    x"3C8CF37",
    x"3C8CD04",
    x"3C8CAD1",
    x"3C8C89E",
    x"3C8C66D",
    x"3C8C43B",
    x"3C8C20A",
    x"3C8BFDA",
    x"3C8BDAB",
    x"3C8BB7B",
    x"3C8B94D",
    x"3C8B71F",
    x"3C8B4F1",
    x"3C8B2C4",
    x"3C8B098",
    x"3C8AE6C",
    x"3C8AC41",
    x"3C8AA16",
    x"3C8A7EC",
    x"3C8A5C2",
    x"3C8A399",
    x"3C8A170",
    x"3C89F48",
    x"3C89D20",
    x"3C89AF9",
    x"3C898D3",
    x"3C896AD",
    x"3C89488",
    x"3C89263",
    x"3C8903E",
    x"3C88E1B",
    x"3C88BF7",
    x"3C889D5",
    x"3C887B2",
    x"3C88591",
    x"3C88370",
    x"3C8814F",
    x"3C87F2F",
    x"3C87D10",
    x"3C87AF1",
    x"3C878D2",
    x"3C876B4",
    x"3C87497",
    x"3C8727A",
    x"3C8705D",
    x"3C86E42",
    x"3C86C26",
    x"3C86A0C",
    x"3C867F1",
    x"3C865D8",
    x"3C863BE",
    x"3C861A6",
    x"3C85F8E",
    x"3C85D76",
    x"3C85B5F",
    x"3C85948",
    x"3C85732",
    x"3C8551D",
    x"3C85308",
    x"3C850F3",
    x"3C84EDF",
    x"3C84CCC",
    x"3C84AB9",
    x"3C848A6",
    x"3C84694",
    x"3C84483",
    x"3C84272",
    x"3C84062",
    x"3C83E52",
    x"3C83C43",
    x"3C83A34",
    x"3C83826",
    x"3C83618",
    x"3C8340A",
    x"3C831FE",
    x"3C82FF1",
    x"3C82DE6",
    x"3C82BDB",
    x"3C829D0",
    x"3C827C6",
    x"3C825BC",
    x"3C823B3",
    x"3C821AA",
    x"3C81FA2",
    x"3C81D9A",
    x"3C81B93",
    x"3C8198C",
    x"3C81786",
    x"3C81581",
    x"3C8137C",
    x"3C81177",
    x"3C80F73",
    x"3C80D6F",
    x"3C80B6C",
    x"3C8096A",
    x"3C80767",
    x"3C80566",
    x"3C80365",
    x"3C80164",
    x"3C7FEC9",
    x"3C7FAC9",
    x"3C7F6CB",
    x"3C7F2CE",
    x"3C7EED2",
    x"3C7EAD7",
    x"3C7E6DC",
    x"3C7E2E3",
    x"3C7DEEB",
    x"3C7DAF4",
    x"3C7D6FD",
    x"3C7D308",
    x"3C7CF14",
    x"3C7CB21",
    x"3C7C72E",
    x"3C7C33D",
    x"3C7BF4D",
    x"3C7BB5D",
    x"3C7B76F",
    x"3C7B382",
    x"3C7AF95",
    x"3C7ABAA",
    x"3C7A7BF",
    x"3C7A3D6",
    x"3C79FEE",
    x"3C79C06",
    x"3C79820",
    x"3C7943A",
    x"3C79055",
    x"3C78C72",
    x"3C7888F",
    x"3C784AE",
    x"3C780CD",
    x"3C77CED",
    x"3C7790E",
    x"3C77531",
    x"3C77154",
    x"3C76D78",
    x"3C7699D",
    x"3C765C3",
    x"3C761EA",
    x"3C75E12",
    x"3C75A3B",
    x"3C75665",
    x"3C75290",
    x"3C74EBC",
    x"3C74AE9",
    x"3C74716",
    x"3C74345",
    x"3C73F75",
    x"3C73BA5",
    x"3C737D7",
    x"3C73409",
    x"3C7303D",
    x"3C72C71",
    x"3C728A7",
    x"3C724DD",
    x"3C72114",
    x"3C71D4C",
    x"3C71986",
    x"3C715C0",
    x"3C711FB",
    x"3C70E37",
    x"3C70A74",
    x"3C706B1",
    x"3C702F0",
    x"3C6FF30",
    x"3C6FB71",
    x"3C6F7B2",
    x"3C6F3F5",
    x"3C6F038",
    x"3C6EC7D",
    x"3C6E8C2",
    x"3C6E508",
    x"3C6E14F",
    x"3C6DD98",
    x"3C6D9E1",
    x"3C6D62B",
    x"3C6D276",
    x"3C6CEC1",
    x"3C6CB0E",
    x"3C6C75C",
    x"3C6C3AB",
    x"3C6BFFA",
    x"3C6BC4B",
    x"3C6B89C",
    x"3C6B4EE",
    x"3C6B141",
    x"3C6AD96",
    x"3C6A9EB",
    x"3C6A641",
    x"3C6A298",
    x"3C69EEF",
    x"3C69B48",
    x"3C697A2",
    x"3C693FC",
    x"3C69058",
    x"3C68CB4",
    x"3C68911",
    x"3C68570",
    x"3C681CF",
    x"3C67E2F",
    x"3C67A90",
    x"3C676F1",
    x"3C67354",
    x"3C66FB8",
    x"3C66C1C",
    x"3C66882",
    x"3C664E8",
    x"3C6614F",
    x"3C65DB7",
    x"3C65A20",
    x"3C6568A",
    x"3C652F5",
    x"3C64F61",
    x"3C64BCD",
    x"3C6483B",
    x"3C644A9",
    x"3C64119",
    x"3C63D89",
    x"3C639FA",
    x"3C6366C",
    x"3C632DF",
    x"3C62F52",
    x"3C62BC7",
    x"3C6283C",
    x"3C624B3",
    x"3C6212A",
    x"3C61DA2",
    x"3C61A1B",
    x"3C61695",
    x"3C61310",
    x"3C60F8C",
    x"3C60C08",
    x"3C60886",
    x"3C60504",
    x"3C60183",
    x"3C5FE03",
    x"3C5FA84",
    x"3C5F706",
    x"3C5F389",
    x"3C5F00C",
    x"3C5EC91",
    x"3C5E916",
    x"3C5E59C",
    x"3C5E223",
    x"3C5DEAB",
    x"3C5DB34",
    x"3C5D7BD",
    x"3C5D448",
    x"3C5D0D3",
    x"3C5CD5F",
    x"3C5C9EC",
    x"3C5C67A",
    x"3C5C309",
    x"3C5BF99",
    x"3C5BC29",
    x"3C5B8BB",
    x"3C5B54D",
    x"3C5B1E0",
    x"3C5AE74",
    x"3C5AB09",
    x"3C5A79F",
    x"3C5A435",
    x"3C5A0CD",
    x"3C59D65",
    x"3C599FE",
    x"3C59698",
    x"3C59333",
    x"3C58FCE",
    x"3C58C6B",
    x"3C58908",
    x"3C585A6",
    x"3C58245",
    x"3C57EE5",
    x"3C57B86",
    x"3C57827",
    x"3C574CA",
    x"3C5716D",
    x"3C56E11",
    x"3C56AB6",
    x"3C5675C",
    x"3C56402",
    x"3C560A9",
    x"3C55D52",
    x"3C559FB",
    x"3C556A5",
    x"3C55350",
    x"3C54FFB",
    x"3C54CA8",
    x"3C54955",
    x"3C54603",
    x"3C542B2",
    x"3C53F62",
    x"3C53C12",
    x"3C538C3",
    x"3C53576",
    x"3C53229",
    x"3C52EDD",
    x"3C52B91",
    x"3C52847",
    x"3C524FD",
    x"3C521B4",
    x"3C51E6C",
    x"3C51B25",
    x"3C517DF",
    x"3C51499",
    x"3C51154",
    x"3C50E11",
    x"3C50ACD",
    x"3C5078B",
    x"3C5044A",
    x"3C50109",
    x"3C4FDC9",
    x"3C4FA8A",
    x"3C4F74C",
    x"3C4F40E",
    x"3C4F0D2",
    x"3C4ED96",
    x"3C4EA5B",
    x"3C4E721",
    x"3C4E3E7",
    x"3C4E0AF",
    x"3C4DD77",
    x"3C4DA40",
    x"3C4D70A",
    x"3C4D3D5",
    x"3C4D0A0",
    x"3C4CD6C",
    x"3C4CA39",
    x"3C4C707",
    x"3C4C3D6",
    x"3C4C0A5",
    x"3C4BD76",
    x"3C4BA47",
    x"3C4B718",
    x"3C4B3EB",
    x"3C4B0BE",
    x"3C4AD93",
    x"3C4AA68",
    x"3C4A73D",
    x"3C4A414",
    x"3C4A0EB",
    x"3C49DC4",
    x"3C49A9D",
    x"3C49776",
    x"3C49451",
    x"3C4912C",
    x"3C48E08",
    x"3C48AE5",
    x"3C487C3",
    x"3C484A1",
    x"3C48180",
    x"3C47E60",
    x"3C47B41",
    x"3C47823",
    x"3C47505",
    x"3C471E8",
    x"3C46ECC",
    x"3C46BB1",
    x"3C46896",
    x"3C4657D",
    x"3C46264",
    x"3C45F4B",
    x"3C45C34",
    x"3C4591D",
    x"3C45607",
    x"3C452F2",
    x"3C44FDE",
    x"3C44CCA",
    x"3C449B8",
    x"3C446A5",
    x"3C44394",
    x"3C44084",
    x"3C43D74",
    x"3C43A65",
    x"3C43757",
    x"3C43449",
    x"3C4313D",
    x"3C42E31",
    x"3C42B26",
    x"3C4281B",
    x"3C42511",
    x"3C42209",
    x"3C41F00",
    x"3C41BF9",
    x"3C418F2",
    x"3C415ED",
    x"3C412E7",
    x"3C40FE3",
    x"3C40CE0",
    x"3C409DD",
    x"3C406DB",
    x"3C403D9",
    x"3C400D9",
    x"3C3FDD9",
    x"3C3FADA",
    x"3C3F7DB",
    x"3C3F4DE",
    x"3C3F1E1",
    x"3C3EEE5",
    x"3C3EBEA",
    x"3C3E8EF",
    x"3C3E5F5",
    x"3C3E2FC",
    x"3C3E004",
    x"3C3DD0C",
    x"3C3DA15",
    x"3C3D71F",
    x"3C3D429",
    x"3C3D135",
    x"3C3CE41",
    x"3C3CB4E",
    x"3C3C85B",
    x"3C3C56A",
    x"3C3C279",
    x"3C3BF88",
    x"3C3BC99",
    x"3C3B9AA",
    x"3C3B6BC",
    x"3C3B3CF",
    x"3C3B0E2",
    x"3C3ADF6",
    x"3C3AB0B",
    x"3C3A821",
    x"3C3A537",
    x"3C3A24E",
    x"3C39F66",
    x"3C39C7E",
    x"3C39998",
    x"3C396B2",
    x"3C393CC",
    x"3C390E8",
    x"3C38E04",
    x"3C38B21",
    x"3C3883E",
    x"3C3855D",
    x"3C3827C",
    x"3C37F9B",
    x"3C37CBC",
    x"3C379DD",
    x"3C376FF",
    x"3C37421",
    x"3C37145",
    x"3C36E69",
    x"3C36B8E",
    x"3C368B3",
    x"3C365D9",
    x"3C36300",
    x"3C36028",
    x"3C35D50",
    x"3C35A79",
    x"3C357A3",
    x"3C354CD",
    x"3C351F8",
    x"3C34F24",
    x"3C34C51",
    x"3C3497E",
    x"3C346AC",
    x"3C343DB",
    x"3C3410A",
    x"3C33E3A",
    x"3C33B6B",
    x"3C3389C",
    x"3C335CF",
    x"3C33302",
    x"3C33035",
    x"3C32D69",
    x"3C32A9E",
    x"3C327D4",
    x"3C3250B",
    x"3C32242",
    x"3C31F79",
    x"3C31CB2",
    x"3C319EB",
    x"3C31725",
    x"3C3145F",
    x"3C3119B",
    x"3C30ED7",
    x"3C30C13",
    x"3C30951",
    x"3C3068F",
    x"3C303CD",
    x"3C3010D",
    x"3C2FE4D",
    x"3C2FB8E",
    x"3C2F8CF",
    x"3C2F611",
    x"3C2F354",
    x"3C2F098",
    x"3C2EDDC",
    x"3C2EB21",
    x"3C2E866",
    x"3C2E5AC",
    x"3C2E2F3",
    x"3C2E03B",
    x"3C2DD83",
    x"3C2DACC",
    x"3C2D816",
    x"3C2D560",
    x"3C2D2AB",
    x"3C2CFF7",
    x"3C2CD43",
    x"3C2CA90",
    x"3C2C7DE",
    x"3C2C52C",
    x"3C2C27B",
    x"3C2BFCB",
    x"3C2BD1B",
    x"3C2BA6C",
    x"3C2B7BE",
    x"3C2B511",
    x"3C2B264",
    x"3C2AFB7",
    x"3C2AD0C",
    x"3C2AA61",
    x"3C2A7B7",
    x"3C2A50D",
    x"3C2A264",
    x"3C29FBC",
    x"3C29D14",
    x"3C29A6D",
    x"3C297C7",
    x"3C29521",
    x"3C2927C",
    x"3C28FD8",
    x"3C28D34",
    x"3C28A92",
    x"3C287EF",
    x"3C2854E",
    x"3C282AD",
    x"3C2800C",
    x"3C27D6D",
    x"3C27ACD",
    x"3C2782F",
    x"3C27591",
    x"3C272F4",
    x"3C27058",
    x"3C26DBC",
    x"3C26B21",
    x"3C26887",
    x"3C265ED",
    x"3C26354",
    x"3C260BB",
    x"3C25E23",
    x"3C25B8C",
    x"3C258F5",
    x"3C25660",
    x"3C253CA",
    x"3C25136",
    x"3C24EA2",
    x"3C24C0E",
    x"3C2497C",
    x"3C246EA",
    x"3C24458",
    x"3C241C7",
    x"3C23F37",
    x"3C23CA8",
    x"3C23A19",
    x"3C2378B",
    x"3C234FD",
    x"3C23270",
    x"3C22FE4",
    x"3C22D58",
    x"3C22ACD",
    x"3C22843",
    x"3C225B9",
    x"3C22330",
    x"3C220A8",
    x"3C21E20",
    x"3C21B99",
    x"3C21912",
    x"3C2168C",
    x"3C21407",
    x"3C21182",
    x"3C20EFE",
    x"3C20C7A",
    x"3C209F8",
    x"3C20776",
    x"3C204F4",
    x"3C20273",
    x"3C1FFF3",
    x"3C1FD73",
    x"3C1FAF4",
    x"3C1F876",
    x"3C1F5F8",
    x"3C1F37B",
    x"3C1F0FE",
    x"3C1EE82",
    x"3C1EC07",
    x"3C1E98C",
    x"3C1E712",
    x"3C1E499",
    x"3C1E220",
    x"3C1DFA7",
    x"3C1DD30",
    x"3C1DAB9",
    x"3C1D843",
    x"3C1D5CD",
    x"3C1D358",
    x"3C1D0E3",
    x"3C1CE6F",
    x"3C1CBFC",
    x"3C1C989",
    x"3C1C717",
    x"3C1C4A6",
    x"3C1C235",
    x"3C1BFC5",
    x"3C1BD55",
    x"3C1BAE6",
    x"3C1B877",
    x"3C1B60A",
    x"3C1B39C",
    x"3C1B130",
    x"3C1AEC4",
    x"3C1AC58",
    x"3C1A9EE",
    x"3C1A783",
    x"3C1A51A",
    x"3C1A2B1",
    x"3C1A049",
    x"3C19DE1",
    x"3C19B7A",
    x"3C19913",
    x"3C196AD",
    x"3C19448",
    x"3C191E3",
    x"3C18F7F",
    x"3C18D1B",
    x"3C18AB8",
    x"3C18856",
    x"3C185F4",
    x"3C18393",
    x"3C18132",
    x"3C17ED2",
    x"3C17C73",
    x"3C17A14",
    x"3C177B6",
    x"3C17558",
    x"3C172FB",
    x"3C1709F",
    x"3C16E43",
    x"3C16BE8",
    x"3C1698D",
    x"3C16733",
    x"3C164D9",
    x"3C16280",
    x"3C16028",
    x"3C15DD0",
    x"3C15B79",
    x"3C15923",
    x"3C156CD",
    x"3C15477",
    x"3C15222",
    x"3C14FCE",
    x"3C14D7A",
    x"3C14B27",
    x"3C148D5",
    x"3C14683",
    x"3C14432",
    x"3C141E1",
    x"3C13F91",
    x"3C13D41",
    x"3C13AF2",
    x"3C138A4",
    x"3C13656",
    x"3C13408",
    x"3C131BC",
    x"3C12F6F",
    x"3C12D24",
    x"3C12AD9",
    x"3C1288E",
    x"3C12645",
    x"3C123FB",
    x"3C121B3",
    x"3C11F6B",
    x"3C11D23",
    x"3C11ADC",
    x"3C11896",
    x"3C11650",
    x"3C1140A",
    x"3C111C6",
    x"3C10F81",
    x"3C10D3E",
    x"3C10AFB",
    x"3C108B8",
    x"3C10676",
    x"3C10435",
    x"3C101F4",
    x"3C0FFB4",
    x"3C0FD75",
    x"3C0FB35",
    x"3C0F8F7",
    x"3C0F6B9",
    x"3C0F47C",
    x"3C0F23F",
    x"3C0F002",
    x"3C0EDC7",
    x"3C0EB8C",
    x"3C0E951",
    x"3C0E717",
    x"3C0E4DD",
    x"3C0E2A4",
    x"3C0E06C",
    x"3C0DE34",
    x"3C0DBFD",
    x"3C0D9C6",
    x"3C0D790",
    x"3C0D55A",
    x"3C0D325",
    x"3C0D0F1",
    x"3C0CEBD",
    x"3C0CC8A",
    x"3C0CA57",
    x"3C0C824",
    x"3C0C5F3",
    x"3C0C3C1",
    x"3C0C191",
    x"3C0BF61",
    x"3C0BD31",
    x"3C0BB02",
    x"3C0B8D4",
    x"3C0B6A6",
    x"3C0B478",
    x"3C0B24B",
    x"3C0B01F",
    x"3C0ADF3",
    x"3C0ABC8",
    x"3C0A99D",
    x"3C0A773",
    x"3C0A54A",
    x"3C0A321",
    x"3C0A0F8",
    x"3C09ED0",
    x"3C09CA9",
    x"3C09A82",
    x"3C0985B",
    x"3C09636",
    x"3C09410",
    x"3C091EC",
    x"3C08FC7",
    x"3C08DA4",
    x"3C08B81",
    x"3C0895E",
    x"3C0873C",
    x"3C0851A",
    x"3C082F9",
    x"3C080D9",
    x"3C07EB9",
    x"3C07C99",
    x"3C07A7B",
    x"3C0785C",
    x"3C0763E",
    x"3C07421",
    x"3C07204",
    x"3C06FE8",
    x"3C06DCC",
    x"3C06BB1",
    x"3C06997",
    x"3C0677C",
    x"3C06563",
    x"3C0634A",
    x"3C06131",
    x"3C05F19",
    x"3C05D02",
    x"3C05AEB",
    x"3C058D4",
    x"3C056BE",
    x"3C054A9",
    x"3C05294",
    x"3C0507F",
    x"3C04E6C",
    x"3C04C58",
    x"3C04A45",
    x"3C04833",
    x"3C04621",
    x"3C04410",
    x"3C041FF",
    x"3C03FEF",
    x"3C03DDF",
    x"3C03BD0",
    x"3C039C1",
    x"3C037B3",
    x"3C035A6",
    x"3C03398",
    x"3C0318C",
    x"3C02F80",
    x"3C02D74",
    x"3C02B69",
    x"3C0295E",
    x"3C02754",
    x"3C0254B",
    x"3C02342",
    x"3C02139",
    x"3C01F31",
    x"3C01D29",
    x"3C01B22",
    x"3C0191C",
    x"3C01716",
    x"3C01510",
    x"3C0130B",
    x"3C01107",
    x"3C00F03",
    x"3C00CFF",
    x"3C00AFC",
    x"3C008FA",
    x"3C006F8",
    x"3C004F6",
    x"3C002F5",
    x"3C000F5",
    x"3BFFDEA",
    x"3BFF9EB",
    x"3BFF5ED",
    x"3BFF1F0",
    x"3BFEDF4",
    x"3BFE9F9",
    x"3BFE5FF",
    x"3BFE206",
    x"3BFDE0E",
    x"3BFDA17",
    x"3BFD621",
    x"3BFD22C",
    x"3BFCE38",
    x"3BFCA45",
    x"3BFC653",
    x"3BFC262",
    x"3BFBE72",
    x"3BFBA83",
    x"3BFB695",
    x"3BFB2A7",
    x"3BFAEBB",
    x"3BFAAD0",
    x"3BFA6E6",
    x"3BFA2FD",
    x"3BF9F14",
    x"3BF9B2D",
    x"3BF9747",
    x"3BF9361",
    x"3BF8F7D",
    x"3BF8B9A",
    x"3BF87B7",
    x"3BF83D6",
    x"3BF7FF5",
    x"3BF7C16",
    x"3BF7837",
    x"3BF745A",
    x"3BF707D",
    x"3BF6CA1",
    x"3BF68C7",
    x"3BF64ED",
    x"3BF6114",
    x"3BF5D3C",
    x"3BF5966",
    x"3BF5590",
    x"3BF51BB",
    x"3BF4DE7",
    x"3BF4A14",
    x"3BF4642",
    x"3BF4271",
    x"3BF3EA1",
    x"3BF3AD1",
    x"3BF3703",
    x"3BF3336",
    x"3BF2F6A",
    x"3BF2B9E",
    x"3BF27D4",
    x"3BF240A",
    x"3BF2042",
    x"3BF1C7A",
    x"3BF18B4",
    x"3BF14EE",
    x"3BF1129",
    x"3BF0D65",
    x"3BF09A2",
    x"3BF05E0",
    x"3BF021F",
    x"3BEFE5F",
    x"3BEFAA0",
    x"3BEF6E2",
    x"3BEF325",
    x"3BEEF69",
    x"3BEEBAD",
    x"3BEE7F3",
    x"3BEE439",
    x"3BEE081",
    x"3BEDCC9",
    x"3BED912",
    x"3BED55C",
    x"3BED1A7",
    x"3BECDF4",
    x"3BECA41",
    x"3BEC68E",
    x"3BEC2DD",
    x"3BEBF2D",
    x"3BEBB7E",
    x"3BEB7CF",
    x"3BEB422",
    x"3BEB075",
    x"3BEACCA",
    x"3BEA91F",
    x"3BEA575",
    x"3BEA1CC",
    x"3BE9E24",
    x"3BE9A7D",
    x"3BE96D7",
    x"3BE9332",
    x"3BE8F8D",
    x"3BE8BEA",
    x"3BE8847",
    x"3BE84A6",
    x"3BE8105",
    x"3BE7D65",
    x"3BE79C6",
    x"3BE7628",
    x"3BE728B",
    x"3BE6EEF",
    x"3BE6B54",
    x"3BE67B9",
    x"3BE6420",
    x"3BE6087",
    x"3BE5CF0",
    x"3BE5959",
    x"3BE55C3",
    x"3BE522E",
    x"3BE4E9A",
    x"3BE4B07",
    x"3BE4774",
    x"3BE43E3",
    x"3BE4052",
    x"3BE3CC3",
    x"3BE3934",
    x"3BE35A6",
    x"3BE3219",
    x"3BE2E8D",
    x"3BE2B02",
    x"3BE2778",
    x"3BE23EE",
    x"3BE2066",
    x"3BE1CDE",
    x"3BE1957",
    x"3BE15D1",
    x"3BE124C",
    x"3BE0EC8",
    x"3BE0B45",
    x"3BE07C2",
    x"3BE0441",
    x"3BE00C0",
    x"3BDFD41",
    x"3BDF9C2",
    x"3BDF644",
    x"3BDF2C7",
    x"3BDEF4A",
    x"3BDEBCF",
    x"3BDE854",
    x"3BDE4DB",
    x"3BDE162",
    x"3BDDDEA",
    x"3BDDA73",
    x"3BDD6FD",
    x"3BDD388",
    x"3BDD013",
    x"3BDCC9F",
    x"3BDC92D",
    x"3BDC5BB",
    x"3BDC24A",
    x"3BDBEDA",
    x"3BDBB6A",
    x"3BDB7FC",
    x"3BDB48E",
    x"3BDB122",
    x"3BDADB6",
    x"3BDAA4B",
    x"3BDA6E1",
    x"3BDA377",
    x"3BDA00F",
    x"3BD9CA7",
    x"3BD9941",
    x"3BD95DB",
    x"3BD9276",
    x"3BD8F12",
    x"3BD8BAE",
    x"3BD884C",
    x"3BD84EA",
    x"3BD8189",
    x"3BD7E29",
    x"3BD7ACA",
    x"3BD776C",
    x"3BD740E",
    x"3BD70B2",
    x"3BD6D56",
    x"3BD69FB",
    x"3BD66A1",
    x"3BD6348",
    x"3BD5FEF",
    x"3BD5C98",
    x"3BD5941",
    x"3BD55EB",
    x"3BD5296",
    x"3BD4F42",
    x"3BD4BEF",
    x"3BD489C",
    x"3BD454A",
    x"3BD41F9",
    x"3BD3EA9",
    x"3BD3B5A",
    x"3BD380C",
    x"3BD34BE",
    x"3BD3171",
    x"3BD2E25",
    x"3BD2ADA",
    x"3BD2790",
    x"3BD2446",
    x"3BD20FE",
    x"3BD1DB6",
    x"3BD1A6F",
    x"3BD1729",
    x"3BD13E3",
    x"3BD109F",
    x"3BD0D5B",
    x"3BD0A18",
    x"3BD06D6",
    x"3BD0395",
    x"3BD0054",
    x"3BCFD14",
    x"3BCF9D6",
    x"3BCF698",
    x"3BCF35A",
    x"3BCF01E",
    x"3BCECE2",
    x"3BCE9A7",
    x"3BCE66D",
    x"3BCE334",
    x"3BCDFFC",
    x"3BCDCC4",
    x"3BCD98D",
    x"3BCD657",
    x"3BCD322",
    x"3BCCFEE",
    x"3BCCCBA",
    x"3BCC988",
    x"3BCC656",
    x"3BCC324",
    x"3BCBFF4",
    x"3BCBCC4",
    x"3BCB996",
    x"3BCB668",
    x"3BCB33A",
    x"3BCB00E",
    x"3BCACE2",
    x"3BCA9B8",
    x"3BCA68D",
    x"3BCA364",
    x"3BCA03C",
    x"3BC9D14",
    x"3BC99ED",
    x"3BC96C7",
    x"3BC93A2",
    x"3BC907D",
    x"3BC8D5A",
    x"3BC8A37",
    x"3BC8715",
    x"3BC83F3",
    x"3BC80D3",
    x"3BC7DB3",
    x"3BC7A94",
    x"3BC7775",
    x"3BC7458",
    x"3BC713B",
    x"3BC6E1F",
    x"3BC6B04",
    x"3BC67EA",
    x"3BC64D0",
    x"3BC61B7",
    x"3BC5E9F",
    x"3BC5B88",
    x"3BC5872",
    x"3BC555C",
    x"3BC5247",
    x"3BC4F33",
    x"3BC4C1F",
    x"3BC490D",
    x"3BC45FB",
    x"3BC42EA",
    x"3BC3FD9",
    x"3BC3CCA",
    x"3BC39BB",
    x"3BC36AD",
    x"3BC33A0",
    x"3BC3093",
    x"3BC2D87",
    x"3BC2A7C",
    x"3BC2772",
    x"3BC2469",
    x"3BC2160",
    x"3BC1E58",
    x"3BC1B51",
    x"3BC184A",
    x"3BC1545",
    x"3BC1240",
    x"3BC0F3B",
    x"3BC0C38",
    x"3BC0935",
    x"3BC0633",
    x"3BC0332",
    x"3BC0032",
    x"3BBFD32",
    x"3BBFA33",
    x"3BBF735",
    x"3BBF438",
    x"3BBF13B",
    x"3BBEE3F",
    x"3BBEB44",
    x"3BBE849",
    x"3BBE550",
    x"3BBE257",
    x"3BBDF5E",
    x"3BBDC67",
    x"3BBD970",
    x"3BBD67A",
    x"3BBD385",
    x"3BBD091",
    x"3BBCD9D",
    x"3BBCAAA",
    x"3BBC7B7",
    x"3BBC4C6",
    x"3BBC1D5",
    x"3BBBEE5",
    x"3BBBBF6",
    x"3BBB907",
    x"3BBB619",
    x"3BBB32C",
    x"3BBB03F",
    x"3BBAD54",
    x"3BBAA69",
    x"3BBA77F",
    x"3BBA495",
    x"3BBA1AC",
    x"3BB9EC4",
    x"3BB9BDD",
    x"3BB98F6",
    x"3BB9610",
    x"3BB932B",
    x"3BB9047",
    x"3BB8D63",
    x"3BB8A80",
    x"3BB879E",
    x"3BB84BC",
    x"3BB81DB",
    x"3BB7EFB",
    x"3BB7C1C",
    x"3BB793D",
    x"3BB765F",
    x"3BB7382",
    x"3BB70A6",
    x"3BB6DCA",
    x"3BB6AEF",
    x"3BB6814",
    x"3BB653B",
    x"3BB6262",
    x"3BB5F89",
    x"3BB5CB2",
    x"3BB59DB",
    x"3BB5705",
    x"3BB5430",
    x"3BB515B",
    x"3BB4E87",
    x"3BB4BB4",
    x"3BB48E1",
    x"3BB460F",
    x"3BB433E",
    x"3BB406E",
    x"3BB3D9E",
    x"3BB3ACF",
    x"3BB3800",
    x"3BB3533",
    x"3BB3266",
    x"3BB2F9A",
    x"3BB2CCE",
    x"3BB2A03",
    x"3BB2739",
    x"3BB2470",
    x"3BB21A7",
    x"3BB1EDF",
    x"3BB1C17",
    x"3BB1951",
    x"3BB168B",
    x"3BB13C5",
    x"3BB1101",
    x"3BB0E3D",
    x"3BB0B7A",
    x"3BB08B7",
    x"3BB05F5",
    x"3BB0334",
    x"3BB0074",
    x"3BAFDB4",
    x"3BAFAF5",
    x"3BAF837",
    x"3BAF579",
    x"3BAF2BC",
    x"3BAEFFF",
    x"3BAED44",
    x"3BAEA89",
    x"3BAE7CF",
    x"3BAE515",
    x"3BAE25C",
    x"3BADFA4",
    x"3BADCEC",
    x"3BADA35",
    x"3BAD77F",
    x"3BAD4CA",
    x"3BAD215",
    x"3BACF60",
    x"3BACCAD",
    x"3BAC9FA",
    x"3BAC748",
    x"3BAC496",
    x"3BAC1E6",
    x"3BABF36",
    x"3BABC86",
    x"3BAB9D7",
    x"3BAB729",
    x"3BAB47C",
    x"3BAB1CF",
    x"3BAAF23",
    x"3BAAC77",
    x"3BAA9CD",
    x"3BAA722",
    x"3BAA479",
    x"3BAA1D0",
    x"3BA9F28",
    x"3BA9C81",
    x"3BA99DA",
    x"3BA9734",
    x"3BA948E",
    x"3BA91E9",
    x"3BA8F45",
    x"3BA8CA2",
    x"3BA89FF",
    x"3BA875D",
    x"3BA84BB",
    x"3BA821A",
    x"3BA7F7A",
    x"3BA7CDB",
    x"3BA7A3C",
    x"3BA779E",
    x"3BA7500",
    x"3BA7263",
    x"3BA6FC7",
    x"3BA6D2B",
    x"3BA6A90",
    x"3BA67F6",
    x"3BA655C",
    x"3BA62C3",
    x"3BA602B",
    x"3BA5D93",
    x"3BA5AFC",
    x"3BA5866",
    x"3BA55D0",
    x"3BA533B",
    x"3BA50A6",
    x"3BA4E12",
    x"3BA4B7F",
    x"3BA48ED",
    x"3BA465B",
    x"3BA43C9",
    x"3BA4139",
    x"3BA3EA9",
    x"3BA3C19",
    x"3BA398B",
    x"3BA36FD",
    x"3BA346F",
    x"3BA31E3",
    x"3BA2F56",
    x"3BA2CCB",
    x"3BA2A40",
    x"3BA27B6",
    x"3BA252C",
    x"3BA22A3",
    x"3BA201B",
    x"3BA1D93",
    x"3BA1B0C",
    x"3BA1886",
    x"3BA1600",
    x"3BA137B",
    x"3BA10F6",
    x"3BA0E72",
    x"3BA0BEF",
    x"3BA096C",
    x"3BA06EA",
    x"3BA0469",
    x"3BA01E8",
    x"3B9FF68",
    x"3B9FCE8",
    x"3B9FA69",
    x"3B9F7EB",
    x"3B9F56D",
    x"3B9F2F0",
    x"3B9F074",
    x"3B9EDF8",
    x"3B9EB7D",
    x"3B9E902",
    x"3B9E688",
    x"3B9E40F",
    x"3B9E196",
    x"3B9DF1E",
    x"3B9DCA7",
    x"3B9DA30",
    x"3B9D7BA",
    x"3B9D544",
    x"3B9D2CF",
    x"3B9D05B",
    x"3B9CDE7",
    x"3B9CB74",
    x"3B9C901",
    x"3B9C68F",
    x"3B9C41E",
    x"3B9C1AD",
    x"3B9BF3D",
    x"3B9BCCD",
    x"3B9BA5F",
    x"3B9B7F0",
    x"3B9B583",
    x"3B9B316",
    x"3B9B0A9",
    x"3B9AE3D",
    x"3B9ABD2",
    x"3B9A967",
    x"3B9A6FD",
    x"3B9A494",
    x"3B9A22B",
    x"3B99FC3",
    x"3B99D5B",
    x"3B99AF4",
    x"3B9988E",
    x"3B99628",
    x"3B993C2",
    x"3B9915E",
    x"3B98EFA",
    x"3B98C96",
    x"3B98A34",
    x"3B987D1",
    x"3B98570",
    x"3B9830F",
    x"3B980AE",
    x"3B97E4E",
    x"3B97BEF",
    x"3B97990",
    x"3B97732",
    x"3B974D5",
    x"3B97278",
    x"3B9701B",
    x"3B96DC0",
    x"3B96B65",
    x"3B9690A",
    x"3B966B0",
    x"3B96457",
    x"3B961FE",
    x"3B95FA6",
    x"3B95D4E",
    x"3B95AF7",
    x"3B958A1",
    x"3B9564B",
    x"3B953F5",
    x"3B951A1",
    x"3B94F4D",
    x"3B94CF9",
    x"3B94AA6",
    x"3B94854",
    x"3B94602",
    x"3B943B1",
    x"3B94160",
    x"3B93F10",
    x"3B93CC1",
    x"3B93A72",
    x"3B93823",
    x"3B935D6",
    x"3B93388",
    x"3B9313C",
    x"3B92EF0",
    x"3B92CA4",
    x"3B92A59",
    x"3B9280F",
    x"3B925C5",
    x"3B9237C",
    x"3B92134",
    x"3B91EEC",
    x"3B91CA4",
    x"3B91A5D",
    x"3B91817",
    x"3B915D1",
    x"3B9138C",
    x"3B91148",
    x"3B90F03",
    x"3B90CC0",
    x"3B90A7D",
    x"3B9083B",
    x"3B905F9",
    x"3B903B8",
    x"3B90177",
    x"3B8FF37",
    x"3B8FCF8",
    x"3B8FAB9",
    x"3B8F87A",
    x"3B8F63C",
    x"3B8F3FF",
    x"3B8F1C2",
    x"3B8EF86",
    x"3B8ED4B",
    x"3B8EB10",
    x"3B8E8D5",
    x"3B8E69B",
    x"3B8E462",
    x"3B8E229",
    x"3B8DFF1",
    x"3B8DDB9",
    x"3B8DB82",
    x"3B8D94B",
    x"3B8D715",
    x"3B8D4E0",
    x"3B8D2AB",
    x"3B8D076",
    x"3B8CE42",
    x"3B8CC0F",
    x"3B8C9DC",
    x"3B8C7AA",
    x"3B8C579",
    x"3B8C348",
    x"3B8C117",
    x"3B8BEE7",
    x"3B8BCB8",
    x"3B8BA89",
    x"3B8B85A",
    x"3B8B62C",
    x"3B8B3FF",
    x"3B8B1D2",
    x"3B8AFA6",
    x"3B8AD7B",
    x"3B8AB4F",
    x"3B8A925",
    x"3B8A6FB",
    x"3B8A4D1",
    x"3B8A2A9",
    x"3B8A080",
    x"3B89E58",
    x"3B89C31",
    x"3B89A0A",
    x"3B897E4",
    x"3B895BE",
    x"3B89399",
    x"3B89174",
    x"3B88F50",
    x"3B88D2D",
    x"3B88B0A",
    x"3B888E7",
    x"3B886C5",
    x"3B884A4",
    x"3B88283",
    x"3B88063",
    x"3B87E43",
    x"3B87C23",
    x"3B87A05",
    x"3B877E6",
    x"3B875C9",
    x"3B873AC",
    x"3B8718F",
    x"3B86F73",
    x"3B86D57",
    x"3B86B3C",
    x"3B86922",
    x"3B86708",
    x"3B864EE",
    x"3B862D5",
    x"3B860BD",
    x"3B85EA5",
    x"3B85C8D",
    x"3B85A76",
    x"3B85860",
    x"3B8564A",
    x"3B85435",
    x"3B85220",
    x"3B8500C",
    x"3B84DF8",
    x"3B84BE5",
    x"3B849D2",
    x"3B847C0",
    x"3B845AE",
    x"3B8439D",
    x"3B8418C",
    x"3B83F7C",
    x"3B83D6D",
    x"3B83B5E",
    x"3B8394F",
    x"3B83741",
    x"3B83533",
    x"3B83326",
    x"3B8311A",
    x"3B82F0E",
    x"3B82D02",
    x"3B82AF7",
    x"3B828ED",
    x"3B826E3",
    x"3B824D9",
    x"3B822D0",
    x"3B820C8",
    x"3B81EC0",
    x"3B81CB9",
    x"3B81AB2",
    x"3B818AB",
    x"3B816A5",
    x"3B814A0",
    x"3B8129B",
    x"3B81097",
    x"3B80E93",
    x"3B80C8F",
    x"3B80A8C",
    x"3B8088A",
    x"3B80688",
    x"3B80487",
    x"3B80286",
    x"3B80086",
    x"3B7FD0C",
    x"3B7F90D",
    x"3B7F50F",
    x"3B7F112",
    x"3B7ED17",
    x"3B7E91C",
    x"3B7E522",
    x"3B7E129",
    x"3B7DD32",
    x"3B7D93B",
    x"3B7D545",
    x"3B7D150",
    x"3B7CD5C",
    x"3B7C969",
    x"3B7C578",
    x"3B7C187",
    x"3B7BD97",
    x"3B7B9A8",
    x"3B7B5BA",
    x"3B7B1CD",
    x"3B7ADE1",
    x"3B7A9F6",
    x"3B7A60C",
    x"3B7A223",
    x"3B79E3B",
    x"3B79A54",
    x"3B7966E",
    x"3B79289",
    x"3B78EA5",
    x"3B78AC1",
    x"3B786DF",
    x"3B782FE",
    x"3B77F1E",
    x"3B77B3E",
    x"3B77760",
    x"3B77383",
    x"3B76FA6",
    x"3B76BCB",
    x"3B767F0",
    x"3B76417",
    x"3B7603E",
    x"3B75C67",
    x"3B75890",
    x"3B754BB",
    x"3B750E6",
    x"3B74D12",
    x"3B7493F",
    x"3B7456D",
    x"3B7419D",
    x"3B73DCD",
    x"3B739FE",
    x"3B73630",
    x"3B73263",
    x"3B72E96",
    x"3B72ACB",
    x"3B72701",
    x"3B72338",
    x"3B71F6F",
    x"3B71BA8",
    x"3B717E2",
    x"3B7141C",
    x"3B71058",
    x"3B70C94",
    x"3B708D1",
    x"3B70510",
    x"3B7014F",
    x"3B6FD8F",
    x"3B6F9D0",
    x"3B6F612",
    x"3B6F255",
    x"3B6EE99",
    x"3B6EADE",
    x"3B6E723",
    x"3B6E36A",
    x"3B6DFB2",
    x"3B6DBFA",
    x"3B6D844",
    x"3B6D48E",
    x"3B6D0D9",
    x"3B6CD26",
    x"3B6C973",
    x"3B6C5C1",
    x"3B6C210",
    x"3B6BE60",
    x"3B6BAB1",
    x"3B6B703",
    x"3B6B355",
    x"3B6AFA9",
    x"3B6ABFD",
    x"3B6A853",
    x"3B6A4A9",
    x"3B6A101",
    x"3B69D59",
    x"3B699B2",
    x"3B6960C",
    x"3B69267",
    x"3B68EC3",
    x"3B68B1F",
    x"3B6877D",
    x"3B683DC",
    x"3B6803B",
    x"3B67C9C",
    x"3B678FD",
    x"3B6755F",
    x"3B671C2",
    x"3B66E26",
    x"3B66A8B",
    x"3B666F1",
    x"3B66358",
    x"3B65FBF",
    x"3B65C28",
    x"3B65891",
    x"3B654FC",
    x"3B65167",
    x"3B64DD3",
    x"3B64A40",
    x"3B646AE",
    x"3B6431C",
    x"3B63F8C",
    x"3B63BFD",
    x"3B6386E",
    x"3B634E0",
    x"3B63154",
    x"3B62DC8",
    x"3B62A3D",
    x"3B626B3",
    x"3B62329",
    x"3B61FA1",
    x"3B61C1A",
    x"3B61893",
    x"3B6150D",
    x"3B61189",
    x"3B60E05",
    x"3B60A82",
    x"3B606FF",
    x"3B6037E",
    x"3B5FFFE",
    x"3B5FC7E",
    x"3B5F8FF",
    x"3B5F582",
    x"3B5F205",
    x"3B5EE89",
    x"3B5EB0D",
    x"3B5E793",
    x"3B5E41A",
    x"3B5E0A1",
    x"3B5DD29",
    x"3B5D9B2",
    x"3B5D63C",
    x"3B5D2C7",
    x"3B5CF53",
    x"3B5CBE0",
    x"3B5C86D",
    x"3B5C4FB",
    x"3B5C18B",
    x"3B5BE1B",
    x"3B5BAAC",
    x"3B5B73D",
    x"3B5B3D0",
    x"3B5B063",
    x"3B5ACF8",
    x"3B5A98D",
    x"3B5A623",
    x"3B5A2BA",
    x"3B59F52",
    x"3B59BEA",
    x"3B59884",
    x"3B5951E",
    x"3B591B9",
    x"3B58E55",
    x"3B58AF2",
    x"3B58790",
    x"3B5842E",
    x"3B580CD",
    x"3B57D6E",
    x"3B57A0F",
    x"3B576B1",
    x"3B57353",
    x"3B56FF7",
    x"3B56C9B",
    x"3B56941",
    x"3B565E7",
    x"3B5628E",
    x"3B55F36",
    x"3B55BDE",
    x"3B55888",
    x"3B55532",
    x"3B551DD",
    x"3B54E89",
    x"3B54B36",
    x"3B547E3",
    x"3B54492",
    x"3B54141",
    x"3B53DF1",
    x"3B53AA2",
    x"3B53754",
    x"3B53406",
    x"3B530BA",
    x"3B52D6E",
    x"3B52A23",
    x"3B526D9",
    x"3B52390",
    x"3B52047",
    x"3B51D00",
    x"3B519B9",
    x"3B51673",
    x"3B5132D",
    x"3B50FE9",
    x"3B50CA6",
    x"3B50963",
    x"3B50621",
    x"3B502E0",
    x"3B4FF9F",
    x"3B4FC60",
    x"3B4F921",
    x"3B4F5E3",
    x"3B4F2A6",
    x"3B4EF6A",
    x"3B4EC2F",
    x"3B4E8F4",
    x"3B4E5BA",
    x"3B4E281",
    x"3B4DF49",
    x"3B4DC11",
    x"3B4D8DB",
    x"3B4D5A5",
    x"3B4D270",
    x"3B4CF3C",
    x"3B4CC08",
    x"3B4C8D6",
    x"3B4C5A4",
    x"3B4C273",
    x"3B4BF43",
    x"3B4BC13",
    x"3B4B8E5",
    x"3B4B5B7",
    x"3B4B28A",
    x"3B4AF5E",
    x"3B4AC32",
    x"3B4A907",
    x"3B4A5DE",
    x"3B4A2B5",
    x"3B49F8C",
    x"3B49C65",
    x"3B4993E",
    x"3B49618",
    x"3B492F3",
    x"3B48FCF",
    x"3B48CAB",
    x"3B48988",
    x"3B48666",
    x"3B48345",
    x"3B48025",
    x"3B47D05",
    x"3B479E6",
    x"3B476C8",
    x"3B473AB",
    x"3B4708E",
    x"3B46D72",
    x"3B46A58",
    x"3B4673D",
    x"3B46424",
    x"3B4610B",
    x"3B45DF3",
    x"3B45ADC",
    x"3B457C6",
    x"3B454B0",
    x"3B4519C",
    x"3B44E88",
    x"3B44B74",
    x"3B44862",
    x"3B44550",
    x"3B4423F",
    x"3B43F2F",
    x"3B43C20",
    x"3B43911",
    x"3B43603",
    x"3B432F6",
    x"3B42FEA",
    x"3B42CDE",
    x"3B429D3",
    x"3B426C9",
    x"3B423C0",
    x"3B420B7",
    x"3B41DAF",
    x"3B41AA8",
    x"3B417A2",
    x"3B4149D",
    x"3B41198",
    x"3B40E94",
    x"3B40B90",
    x"3B4088E",
    x"3B4058C",
    x"3B4028B",
    x"3B3FF8B",
    x"3B3FC8B",
    x"3B3F98D",
    x"3B3F68F",
    x"3B3F391",
    x"3B3F095",
    x"3B3ED99",
    x"3B3EA9E",
    x"3B3E7A4",
    x"3B3E4AA",
    x"3B3E1B1",
    x"3B3DEB9",
    x"3B3DBC2",
    x"3B3D8CB",
    x"3B3D5D6",
    x"3B3D2E1",
    x"3B3CFEC",
    x"3B3CCF9",
    x"3B3CA06",
    x"3B3C714",
    x"3B3C422",
    x"3B3C132",
    x"3B3BE42",
    x"3B3BB52",
    x"3B3B864",
    x"3B3B576",
    x"3B3B289",
    x"3B3AF9D",
    x"3B3ACB1",
    x"3B3A9C7",
    x"3B3A6DD",
    x"3B3A3F3",
    x"3B3A10B",
    x"3B39E23",
    x"3B39B3B",
    x"3B39855",
    x"3B3956F",
    x"3B3928A",
    x"3B38FA6",
    x"3B38CC2",
    x"3B389E0",
    x"3B386FE",
    x"3B3841C",
    x"3B3813B",
    x"3B37E5C",
    x"3B37B7C",
    x"3B3789E",
    x"3B375C0",
    x"3B372E3",
    x"3B37007",
    x"3B36D2B",
    x"3B36A50",
    x"3B36776",
    x"3B3649C",
    x"3B361C3",
    x"3B35EEB",
    x"3B35C14",
    x"3B3593D",
    x"3B35667",
    x"3B35392",
    x"3B350BE",
    x"3B34DEA",
    x"3B34B17",
    x"3B34844",
    x"3B34572",
    x"3B342A1",
    x"3B33FD1",
    x"3B33D02",
    x"3B33A33",
    x"3B33764",
    x"3B33497",
    x"3B331CA",
    x"3B32EFE",
    x"3B32C33",
    x"3B32968",
    x"3B3269E",
    x"3B323D5",
    x"3B3210C",
    x"3B31E44",
    x"3B31B7D",
    x"3B318B6",
    x"3B315F1",
    x"3B3132B",
    x"3B31067",
    x"3B30DA3",
    x"3B30AE0",
    x"3B3081E",
    x"3B3055C",
    x"3B3029B",
    x"3B2FFDB",
    x"3B2FD1B",
    x"3B2FA5C",
    x"3B2F79E",
    x"3B2F4E0",
    x"3B2F224",
    x"3B2EF67",
    x"3B2ECAC",
    x"3B2E9F1",
    x"3B2E737",
    x"3B2E47D",
    x"3B2E1C5",
    x"3B2DF0D",
    x"3B2DC55",
    x"3B2D99E",
    x"3B2D6E8",
    x"3B2D433",
    x"3B2D17E",
    x"3B2CECA",
    x"3B2CC17",
    x"3B2C964",
    x"3B2C6B2",
    x"3B2C401",
    x"3B2C150",
    x"3B2BEA0",
    x"3B2BBF1",
    x"3B2B942",
    x"3B2B694",
    x"3B2B3E7",
    x"3B2B13A",
    x"3B2AE8E",
    x"3B2ABE3",
    x"3B2A938",
    x"3B2A68E",
    x"3B2A3E5",
    x"3B2A13C",
    x"3B29E94",
    x"3B29BED",
    x"3B29946",
    x"3B296A0",
    x"3B293FB",
    x"3B29156",
    x"3B28EB2",
    x"3B28C0F",
    x"3B2896C",
    x"3B286CA",
    x"3B28429",
    x"3B28188",
    x"3B27EE8",
    x"3B27C49",
    x"3B279AA",
    x"3B2770C",
    x"3B2746F",
    x"3B271D2",
    x"3B26F36",
    x"3B26C9A",
    x"3B269FF",
    x"3B26765",
    x"3B264CC",
    x"3B26233",
    x"3B25F9B",
    x"3B25D03",
    x"3B25A6C",
    x"3B257D6",
    x"3B25540",
    x"3B252AB",
    x"3B25017",
    x"3B24D83",
    x"3B24AF0",
    x"3B2485E",
    x"3B245CC",
    x"3B2433B",
    x"3B240AA",
    x"3B23E1A",
    x"3B23B8B",
    x"3B238FD",
    x"3B2366F",
    x"3B233E1",
    x"3B23155",
    x"3B22EC9",
    x"3B22C3D",
    x"3B229B3",
    x"3B22729",
    x"3B2249F",
    x"3B22216",
    x"3B21F8E",
    x"3B21D06",
    x"3B21A7F",
    x"3B217F9",
    x"3B21573",
    x"3B212EE",
    x"3B2106A",
    x"3B20DE6",
    x"3B20B63",
    x"3B208E1",
    x"3B2065F",
    x"3B203DD",
    x"3B2015D",
    x"3B1FEDD",
    x"3B1FC5D",
    x"3B1F9DE",
    x"3B1F760",
    x"3B1F4E3",
    x"3B1F266",
    x"3B1EFEA",
    x"3B1ED6E",
    x"3B1EAF3",
    x"3B1E878",
    x"3B1E5FF",
    x"3B1E385",
    x"3B1E10D",
    x"3B1DE95",
    x"3B1DC1E",
    x"3B1D9A7",
    x"3B1D731",
    x"3B1D4BB",
    x"3B1D246",
    x"3B1CFD2",
    x"3B1CD5E",
    x"3B1CAEB",
    x"3B1C879",
    x"3B1C607",
    x"3B1C396",
    x"3B1C125",
    x"3B1BEB5",
    x"3B1BC46",
    x"3B1B9D7",
    x"3B1B769",
    x"3B1B4FC",
    x"3B1B28F",
    x"3B1B022",
    x"3B1ADB7",
    x"3B1AB4B",
    x"3B1A8E1",
    x"3B1A677",
    x"3B1A40E",
    x"3B1A1A5",
    x"3B19F3D",
    x"3B19CD5",
    x"3B19A6E",
    x"3B19808",
    x"3B195A2",
    x"3B1933D",
    x"3B190D9",
    x"3B18E75",
    x"3B18C12",
    x"3B189AF",
    x"3B1874D",
    x"3B184EB",
    x"3B1828A",
    x"3B1802A",
    x"3B17DCA",
    x"3B17B6B",
    x"3B1790C",
    x"3B176AF",
    x"3B17451",
    x"3B171F4",
    x"3B16F98",
    x"3B16D3D",
    x"3B16AE2",
    x"3B16887",
    x"3B1662D",
    x"3B163D4",
    x"3B1617B",
    x"3B15F23",
    x"3B15CCC",
    x"3B15A75",
    x"3B1581F",
    x"3B155C9",
    x"3B15374",
    x"3B1511F",
    x"3B14ECB",
    x"3B14C78",
    x"3B14A25",
    x"3B147D3",
    x"3B14581",
    x"3B14330",
    x"3B140DF",
    x"3B13E8F",
    x"3B13C40",
    x"3B139F1",
    x"3B137A3",
    x"3B13555",
    x"3B13308",
    x"3B130BC",
    x"3B12E70",
    x"3B12C25",
    x"3B129DA",
    x"3B12790",
    x"3B12546",
    x"3B122FD",
    x"3B120B5",
    x"3B11E6D",
    x"3B11C26",
    x"3B119DF",
    x"3B11799",
    x"3B11553",
    x"3B1130E",
    x"3B110C9",
    x"3B10E86",
    x"3B10C42",
    x"3B109FF",
    x"3B107BD",
    x"3B1057C",
    x"3B1033A",
    x"3B100FA",
    x"3B0FEBA",
    x"3B0FC7B",
    x"3B0FA3C",
    x"3B0F7FD",
    x"3B0F5C0",
    x"3B0F383",
    x"3B0F146",
    x"3B0EF0A",
    x"3B0ECCE",
    x"3B0EA94",
    x"3B0E859",
    x"3B0E61F",
    x"3B0E3E6",
    x"3B0E1AD",
    x"3B0DF75",
    x"3B0DD3E",
    x"3B0DB07",
    x"3B0D8D0",
    x"3B0D69A",
    x"3B0D465",
    x"3B0D230",
    x"3B0CFFC",
    x"3B0CDC8",
    x"3B0CB95",
    x"3B0C962",
    x"3B0C730",
    x"3B0C4FF",
    x"3B0C2CE",
    x"3B0C09D",
    x"3B0BE6D",
    x"3B0BC3E",
    x"3B0BA0F",
    x"3B0B7E1",
    x"3B0B5B3",
    x"3B0B386",
    x"3B0B15A",
    x"3B0AF2D",
    x"3B0AD02",
    x"3B0AAD7",
    x"3B0A8AD",
    x"3B0A683",
    x"3B0A459",
    x"3B0A230",
    x"3B0A008",
    x"3B09DE0",
    x"3B09BB9",
    x"3B09993",
    x"3B0976C",
    x"3B09547",
    x"3B09322",
    x"3B090FD",
    x"3B08ED9",
    x"3B08CB6",
    x"3B08A93",
    x"3B08871",
    x"3B0864F",
    x"3B0842D",
    x"3B0820D",
    x"3B07FEC",
    x"3B07DCD",
    x"3B07BAD",
    x"3B0798F",
    x"3B07771",
    x"3B07553",
    x"3B07336",
    x"3B0711A",
    x"3B06EFD",
    x"3B06CE2",
    x"3B06AC7",
    x"3B068AD",
    x"3B06693",
    x"3B06479",
    x"3B06260",
    x"3B06048",
    x"3B05E30",
    x"3B05C19",
    x"3B05A02",
    x"3B057EC",
    x"3B055D6",
    x"3B053C1",
    x"3B051AC",
    x"3B04F98",
    x"3B04D85",
    x"3B04B72",
    x"3B0495F",
    x"3B0474D",
    x"3B0453B",
    x"3B0432A",
    x"3B0411A",
    x"3B03F0A",
    x"3B03CFA",
    x"3B03AEB",
    x"3B038DD",
    x"3B036CF",
    x"3B034C1",
    x"3B032B4",
    x"3B030A8",
    x"3B02E9C",
    x"3B02C91",
    x"3B02A86",
    x"3B0287B",
    x"3B02672",
    x"3B02468",
    x"3B0225F",
    x"3B02057",
    x"3B01E4F",
    x"3B01C48",
    x"3B01A41",
    x"3B0183B",
    x"3B01635",
    x"3B01430",
    x"3B0122B",
    x"3B01026",
    x"3B00E23",
    x"3B00C1F",
    x"3B00A1D",
    x"3B0081A",
    x"3B00619",
    x"3B00417",
    x"3B00217",
    x"3B00016",
    x"3AFFC2D",
    x"3AFF82F",
    x"3AFF431",
    x"3AFF035",
    x"3AFEC39",
    x"3AFE83F",
    x"3AFE445",
    x"3AFE04D",
    x"3AFDC55",
    x"3AFD85E",
    x"3AFD469",
    x"3AFD074",
    x"3AFCC81",
    x"3AFC88E",
    x"3AFC49C",
    x"3AFC0AC",
    x"3AFBCBC",
    x"3AFB8CD",
    x"3AFB4E0",
    x"3AFB0F3",
    x"3AFAD07",
    x"3AFA91C",
    x"3AFA533",
    x"3AFA14A",
    x"3AF9D62",
    x"3AF997B",
    x"3AF9595",
    x"3AF91B0",
    x"3AF8DCC",
    x"3AF89E9",
    x"3AF8607",
    x"3AF8226",
    x"3AF7E46",
    x"3AF7A67",
    x"3AF7689",
    x"3AF72AC",
    x"3AF6ED0",
    x"3AF6AF5",
    x"3AF671A",
    x"3AF6341",
    x"3AF5F69",
    x"3AF5B91",
    x"3AF57BB",
    x"3AF53E5",
    x"3AF5011",
    x"3AF4C3D",
    x"3AF486B",
    x"3AF4499",
    x"3AF40C8",
    x"3AF3CF9",
    x"3AF392A",
    x"3AF355C",
    x"3AF318F",
    x"3AF2DC3",
    x"3AF29F8",
    x"3AF262E",
    x"3AF2265",
    x"3AF1E9D",
    x"3AF1AD6",
    x"3AF1710",
    x"3AF134A",
    x"3AF0F86",
    x"3AF0BC3",
    x"3AF0800",
    x"3AF043F",
    x"3AF007E",
    x"3AEFCBE",
    x"3AEF900",
    x"3AEF542",
    x"3AEF185",
    x"3AEEDC9",
    x"3AEEA0E",
    x"3AEE654",
    x"3AEE29B",
    x"3AEDEE3",
    x"3AEDB2C",
    x"3AED775",
    x"3AED3C0",
    x"3AED00B",
    x"3AECC58",
    x"3AEC8A5",
    x"3AEC4F4",
    x"3AEC143",
    x"3AEBD93",
    x"3AEB9E4",
    x"3AEB636",
    x"3AEB289",
    x"3AEAEDD",
    x"3AEAB31",
    x"3AEA787",
    x"3AEA3DE",
    x"3AEA035",
    x"3AE9C8E",
    x"3AE98E7",
    x"3AE9541",
    x"3AE919C",
    x"3AE8DF8",
    x"3AE8A55",
    x"3AE86B3",
    x"3AE8312",
    x"3AE7F72",
    x"3AE7BD2",
    x"3AE7834",
    x"3AE7496",
    x"3AE70F9",
    x"3AE6D5E",
    x"3AE69C3",
    x"3AE6629",
    x"3AE6290",
    x"3AE5EF7",
    x"3AE5B60",
    x"3AE57CA",
    x"3AE5434",
    x"3AE50A0",
    x"3AE4D0C",
    x"3AE4979",
    x"3AE45E7",
    x"3AE4256",
    x"3AE3EC6",
    x"3AE3B37",
    x"3AE37A8",
    x"3AE341B",
    x"3AE308E",
    x"3AE2D03",
    x"3AE2978",
    x"3AE25EE",
    x"3AE2265",
    x"3AE1EDD",
    x"3AE1B55",
    x"3AE17CF",
    x"3AE144A",
    x"3AE10C5",
    x"3AE0D41",
    x"3AE09BE",
    x"3AE063C",
    x"3AE02BB",
    x"3ADFF3B",
    x"3ADFBBC",
    x"3ADF83D",
    x"3ADF4BF",
    x"3ADF143",
    x"3ADEDC7",
    x"3ADEA4C",
    x"3ADE6D2",
    x"3ADE358",
    x"3ADDFE0",
    x"3ADDC68",
    x"3ADD8F2",
    x"3ADD57C",
    x"3ADD207",
    x"3ADCE93",
    x"3ADCB20",
    x"3ADC7AD",
    x"3ADC43C",
    x"3ADC0CB",
    x"3ADBD5C",
    x"3ADB9ED",
    x"3ADB67F",
    x"3ADB311",
    x"3ADAFA5",
    x"3ADAC3A",
    x"3ADA8CF",
    x"3ADA565",
    x"3ADA1FC",
    x"3AD9E94",
    x"3AD9B2D",
    x"3AD97C7",
    x"3AD9461",
    x"3AD90FC",
    x"3AD8D99",
    x"3AD8A36",
    x"3AD86D3",
    x"3AD8372",
    x"3AD8012",
    x"3AD7CB2",
    x"3AD7953",
    x"3AD75F5",
    x"3AD7298",
    x"3AD6F3C",
    x"3AD6BE1",
    x"3AD6886",
    x"3AD652C",
    x"3AD61D4",
    x"3AD5E7C",
    x"3AD5B24",
    x"3AD57CE",
    x"3AD5478",
    x"3AD5124",
    x"3AD4DD0",
    x"3AD4A7D",
    x"3AD472B",
    x"3AD43D9",
    x"3AD4089",
    x"3AD3D39",
    x"3AD39EA",
    x"3AD369C",
    x"3AD334F",
    x"3AD3002",
    x"3AD2CB7",
    x"3AD296C",
    x"3AD2622",
    x"3AD22D9",
    x"3AD1F91",
    x"3AD1C49",
    x"3AD1903",
    x"3AD15BD",
    x"3AD1278",
    x"3AD0F33",
    x"3AD0BF0",
    x"3AD08AD",
    x"3AD056C",
    x"3AD022B",
    x"3ACFEEB",
    x"3ACFBAB",
    x"3ACF86D",
    x"3ACF52F",
    x"3ACF1F2",
    x"3ACEEB6",
    x"3ACEB7B",
    x"3ACE840",
    x"3ACE507",
    x"3ACE1CE",
    x"3ACDE96",
    x"3ACDB5F",
    x"3ACD828",
    x"3ACD4F2",
    x"3ACD1BE",
    x"3ACCE8A",
    x"3ACCB56",
    x"3ACC824",
    x"3ACC4F2",
    x"3ACC1C1",
    x"3ACBE91",
    x"3ACBB62",
    x"3ACB834",
    x"3ACB506",
    x"3ACB1D9",
    x"3ACAEAD",
    x"3ACAB82",
    x"3ACA857",
    x"3ACA52E",
    x"3ACA205",
    x"3AC9EDD",
    x"3AC9BB5",
    x"3AC988F",
    x"3AC9569",
    x"3AC9244",
    x"3AC8F20",
    x"3AC8BFD",
    x"3AC88DA",
    x"3AC85B8",
    x"3AC8297",
    x"3AC7F77",
    x"3AC7C57",
    x"3AC7939",
    x"3AC761B",
    x"3AC72FE",
    x"3AC6FE1",
    x"3AC6CC6",
    x"3AC69AB",
    x"3AC6691",
    x"3AC6378",
    x"3AC605F",
    x"3AC5D47",
    x"3AC5A30",
    x"3AC571A",
    x"3AC5405",
    x"3AC50F0",
    x"3AC4DDC",
    x"3AC4AC9",
    x"3AC47B7",
    x"3AC44A6",
    x"3AC4195",
    x"3AC3E85",
    x"3AC3B75",
    x"3AC3867",
    x"3AC3559",
    x"3AC324C",
    x"3AC2F40",
    x"3AC2C35",
    x"3AC292A",
    x"3AC2620",
    x"3AC2317",
    x"3AC200F",
    x"3AC1D07",
    x"3AC1A00",
    x"3AC16FA",
    x"3AC13F5",
    x"3AC10F0",
    x"3AC0DEC",
    x"3AC0AE9",
    x"3AC07E7",
    x"3AC04E5",
    x"3AC01E4",
    x"3ABFEE4",
    x"3ABFBE5",
    x"3ABF8E6",
    x"3ABF5E8",
    x"3ABF2EB",
    x"3ABEFEF",
    x"3ABECF3",
    x"3ABE9F8",
    x"3ABE6FE",
    x"3ABE405",
    x"3ABE10C",
    x"3ABDE14",
    x"3ABDB1D",
    x"3ABD827",
    x"3ABD531",
    x"3ABD23C",
    x"3ABCF48",
    x"3ABCC55",
    x"3ABC962",
    x"3ABC670",
    x"3ABC37F",
    x"3ABC08E",
    x"3ABBD9E",
    x"3ABBAAF",
    x"3ABB7C1",
    x"3ABB4D3",
    x"3ABB1E7",
    x"3ABAEFA",
    x"3ABAC0F",
    x"3ABA924",
    x"3ABA63A",
    x"3ABA351",
    x"3ABA069",
    x"3AB9D81",
    x"3AB9A9A",
    x"3AB97B4",
    x"3AB94CE",
    x"3AB91E9",
    x"3AB8F05",
    x"3AB8C22",
    x"3AB893F",
    x"3AB865D",
    x"3AB837C",
    x"3AB809C",
    x"3AB7DBC",
    x"3AB7ADD",
    x"3AB77FE",
    x"3AB7521",
    x"3AB7244",
    x"3AB6F68",
    x"3AB6C8C",
    x"3AB69B1",
    x"3AB66D7",
    x"3AB63FE",
    x"3AB6125",
    x"3AB5E4D",
    x"3AB5B76",
    x"3AB58A0",
    x"3AB55CA",
    x"3AB52F5",
    x"3AB5020",
    x"3AB4D4D",
    x"3AB4A7A",
    x"3AB47A7",
    x"3AB44D6",
    x"3AB4205",
    x"3AB3F35",
    x"3AB3C65",
    x"3AB3997",
    x"3AB36C8",
    x"3AB33FB",
    x"3AB312F",
    x"3AB2E63",
    x"3AB2B97",
    x"3AB28CD",
    x"3AB2603",
    x"3AB233A",
    x"3AB2071",
    x"3AB1DAA",
    x"3AB1AE2",
    x"3AB181C",
    x"3AB1556",
    x"3AB1291",
    x"3AB0FCD",
    x"3AB0D0A",
    x"3AB0A47",
    x"3AB0784",
    x"3AB04C3",
    x"3AB0202",
    x"3AAFF42",
    x"3AAFC82",
    x"3AAF9C4",
    x"3AAF705",
    x"3AAF448",
    x"3AAF18B",
    x"3AAEECF",
    x"3AAEC14",
    x"3AAE959",
    x"3AAE69F",
    x"3AAE3E6",
    x"3AAE12D",
    x"3AADE75",
    x"3AADBBE",
    x"3AAD907",
    x"3AAD652",
    x"3AAD39C",
    x"3AAD0E8",
    x"3AACE34",
    x"3AACB81",
    x"3AAC8CE",
    x"3AAC61C",
    x"3AAC36B",
    x"3AAC0BB",
    x"3AABE0B",
    x"3AABB5C",
    x"3AAB8AD",
    x"3AAB5FF",
    x"3AAB352",
    x"3AAB0A6",
    x"3AAADFA",
    x"3AAAB4F",
    x"3AAA8A4",
    x"3AAA5FA",
    x"3AAA351",
    x"3AAA0A9",
    x"3AA9E01",
    x"3AA9B5A",
    x"3AA98B3",
    x"3AA960D",
    x"3AA9368",
    x"3AA90C3",
    x"3AA8E20",
    x"3AA8B7C",
    x"3AA88DA",
    x"3AA8638",
    x"3AA8397",
    x"3AA80F6",
    x"3AA7E56",
    x"3AA7BB7",
    x"3AA7918",
    x"3AA767A",
    x"3AA73DD",
    x"3AA7141",
    x"3AA6EA5",
    x"3AA6C09",
    x"3AA696F",
    x"3AA66D5",
    x"3AA643B",
    x"3AA61A2",
    x"3AA5F0A",
    x"3AA5C73",
    x"3AA59DC",
    x"3AA5746",
    x"3AA54B0",
    x"3AA521C",
    x"3AA4F87",
    x"3AA4CF4",
    x"3AA4A61",
    x"3AA47CF",
    x"3AA453D",
    x"3AA42AC",
    x"3AA401C",
    x"3AA3D8C",
    x"3AA3AFD",
    x"3AA386E",
    x"3AA35E1",
    x"3AA3354",
    x"3AA30C7",
    x"3AA2E3B",
    x"3AA2BB0",
    x"3AA2925",
    x"3AA269B",
    x"3AA2412",
    x"3AA2189",
    x"3AA1F01",
    x"3AA1C7A",
    x"3AA19F3",
    x"3AA176D",
    x"3AA14E7",
    x"3AA1262",
    x"3AA0FDE",
    x"3AA0D5A",
    x"3AA0AD7",
    x"3AA0855",
    x"3AA05D3",
    x"3AA0352",
    x"3AA00D2",
    x"3A9FE52",
    x"3A9FBD2",
    x"3A9F954",
    x"3A9F6D6",
    x"3A9F458",
    x"3A9F1DC",
    x"3A9EF5F",
    x"3A9ECE4",
    x"3A9EA69",
    x"3A9E7EF",
    x"3A9E575",
    x"3A9E2FC",
    x"3A9E084",
    x"3A9DE0C",
    x"3A9DB94",
    x"3A9D91E",
    x"3A9D6A8",
    x"3A9D433",
    x"3A9D1BE",
    x"3A9CF4A",
    x"3A9CCD6",
    x"3A9CA63",
    x"3A9C7F1",
    x"3A9C57F",
    x"3A9C30E",
    x"3A9C09E",
    x"3A9BE2E",
    x"3A9BBBF",
    x"3A9B950",
    x"3A9B6E2",
    x"3A9B475",
    x"3A9B208",
    x"3A9AF9C",
    x"3A9AD30",
    x"3A9AAC5",
    x"3A9A85B",
    x"3A9A5F1",
    x"3A9A388",
    x"3A9A11F",
    x"3A99EB7",
    x"3A99C50",
    x"3A999E9",
    x"3A99783",
    x"3A9951D",
    x"3A992B8",
    x"3A99054",
    x"3A98DF0",
    x"3A98B8D",
    x"3A9892A",
    x"3A986C8",
    x"3A98467",
    x"3A98206",
    x"3A97FA6",
    x"3A97D46",
    x"3A97AE7",
    x"3A97889",
    x"3A9762B",
    x"3A973CE",
    x"3A97171",
    x"3A96F15",
    x"3A96CB9",
    x"3A96A5F",
    x"3A96804",
    x"3A965AB",
    x"3A96351",
    x"3A960F9",
    x"3A95EA1",
    x"3A95C4A",
    x"3A959F3",
    x"3A9579D",
    x"3A95547",
    x"3A952F2",
    x"3A9509E",
    x"3A94E4A",
    x"3A94BF6",
    x"3A949A4",
    x"3A94752",
    x"3A94500",
    x"3A942AF",
    x"3A9405F",
    x"3A93E0F",
    x"3A93BC0",
    x"3A93971",
    x"3A93723",
    x"3A934D5",
    x"3A93289",
    x"3A9303C",
    x"3A92DF0",
    x"3A92BA5",
    x"3A9295B",
    x"3A92711",
    x"3A924C7",
    x"3A9227E",
    x"3A92036",
    x"3A91DEE",
    x"3A91BA7",
    x"3A91960",
    x"3A9171A",
    x"3A914D5",
    x"3A91290",
    x"3A9104B",
    x"3A90E08",
    x"3A90BC4",
    x"3A90982",
    x"3A90740",
    x"3A904FE",
    x"3A902BD",
    x"3A9007D",
    x"3A8FE3D",
    x"3A8FBFE",
    x"3A8F9BF",
    x"3A8F781",
    x"3A8F543",
    x"3A8F306",
    x"3A8F0CA",
    x"3A8EE8E",
    x"3A8EC52",
    x"3A8EA18",
    x"3A8E7DD",
    x"3A8E5A4",
    x"3A8E36A",
    x"3A8E132",
    x"3A8DEFA",
    x"3A8DCC2",
    x"3A8DA8B",
    x"3A8D855",
    x"3A8D61F",
    x"3A8D3EA",
    x"3A8D1B5",
    x"3A8CF81",
    x"3A8CD4E",
    x"3A8CB1B",
    x"3A8C8E8",
    x"3A8C6B6",
    x"3A8C485",
    x"3A8C254",
    x"3A8C024",
    x"3A8BDF4",
    x"3A8BBC5",
    x"3A8B996",
    x"3A8B768",
    x"3A8B53A",
    x"3A8B30D",
    x"3A8B0E1",
    x"3A8AEB5",
    x"3A8AC89",
    x"3A8AA5E",
    x"3A8A834",
    x"3A8A60A",
    x"3A8A3E1",
    x"3A8A1B8",
    x"3A89F90",
    x"3A89D69",
    x"3A89B42",
    x"3A8991B",
    x"3A896F5",
    x"3A894CF",
    x"3A892AB",
    x"3A89086",
    x"3A88E62",
    x"3A88C3F",
    x"3A88A1C",
    x"3A887FA",
    x"3A885D8",
    x"3A883B7",
    x"3A88196",
    x"3A87F76",
    x"3A87D57",
    x"3A87B38",
    x"3A87919",
    x"3A876FB",
    x"3A874DD",
    x"3A872C1",
    x"3A870A4",
    x"3A86E88",
    x"3A86C6D",
    x"3A86A52",
    x"3A86838",
    x"3A8661E",
    x"3A86405",
    x"3A861EC",
    x"3A85FD4",
    x"3A85DBC",
    x"3A85BA5",
    x"3A8598E",
    x"3A85778",
    x"3A85562",
    x"3A8534D",
    x"3A85139",
    x"3A84F25",
    x"3A84D11",
    x"3A84AFE",
    x"3A848EC",
    x"3A846DA",
    x"3A844C8",
    x"3A842B7",
    x"3A840A7",
    x"3A83E97",
    x"3A83C88",
    x"3A83A79",
    x"3A8386A",
    x"3A8365D",
    x"3A8344F",
    x"3A83242",
    x"3A83036",
    x"3A82E2A",
    x"3A82C1F",
    x"3A82A14",
    x"3A8280A",
    x"3A82600",
    x"3A823F7",
    x"3A821EE",
    x"3A81FE6",
    x"3A81DDE",
    x"3A81BD7",
    x"3A819D0",
    x"3A817CA",
    x"3A815C4",
    x"3A813BF",
    x"3A811BB",
    x"3A80FB6",
    x"3A80DB3",
    x"3A80BB0",
    x"3A809AD",
    x"3A807AB",
    x"3A805A9",
    x"3A803A8",
    x"3A801A7",
    x"3A7FF4F",
    x"3A7FB4F",
    x"3A7F751",
    x"3A7F354",
    x"3A7EF57",
    x"3A7EB5C",
    x"3A7E762",
    x"3A7E368",
    x"3A7DF70",
    x"3A7DB78",
    x"3A7D782",
    x"3A7D38D",
    x"3A7CF98",
    x"3A7CBA5",
    x"3A7C7B2",
    x"3A7C3C1",
    x"3A7BFD1",
    x"3A7BBE1",
    x"3A7B7F3",
    x"3A7B405",
    x"3A7B019",
    x"3A7AC2D",
    x"3A7A843",
    x"3A7A459",
    x"3A7A070",
    x"3A79C89",
    x"3A798A2",
    x"3A794BC",
    x"3A790D8",
    x"3A78CF4",
    x"3A78911",
    x"3A7852F",
    x"3A7814F",
    x"3A77D6F",
    x"3A77990",
    x"3A775B2",
    x"3A771D5",
    x"3A76DF9",
    x"3A76A1E",
    x"3A76644",
    x"3A7626B",
    x"3A75E93",
    x"3A75ABC",
    x"3A756E5",
    x"3A75310",
    x"3A74F3C",
    x"3A74B69",
    x"3A74796",
    x"3A743C5",
    x"3A73FF4",
    x"3A73C25",
    x"3A73856",
    x"3A73489",
    x"3A730BC",
    x"3A72CF0",
    x"3A72926",
    x"3A7255C",
    x"3A72193",
    x"3A71DCB",
    x"3A71A04",
    x"3A7163E",
    x"3A71279",
    x"3A70EB5",
    x"3A70AF2",
    x"3A7072F",
    x"3A7036E",
    x"3A6FFAE",
    x"3A6FBEE",
    x"3A6F830",
    x"3A6F472",
    x"3A6F0B5",
    x"3A6ECFA",
    x"3A6E93F",
    x"3A6E585",
    x"3A6E1CC",
    x"3A6DE14",
    x"3A6DA5D",
    x"3A6D6A7",
    x"3A6D2F2",
    x"3A6CF3D",
    x"3A6CB8A",
    x"3A6C7D8",
    x"3A6C426",
    x"3A6C076",
    x"3A6BCC6",
    x"3A6B917",
    x"3A6B569",
    x"3A6B1BD",
    x"3A6AE11",
    x"3A6AA65",
    x"3A6A6BB",
    x"3A6A312",
    x"3A69F6A",
    x"3A69BC2",
    x"3A6981C",
    x"3A69476",
    x"3A690D2",
    x"3A68D2E",
    x"3A6898B",
    x"3A685E9",
    x"3A68248",
    x"3A67EA8",
    x"3A67B09",
    x"3A6776A",
    x"3A673CD",
    x"3A67031",
    x"3A66C95",
    x"3A668FA",
    x"3A66561",
    x"3A661C8",
    x"3A65E30",
    x"3A65A99",
    x"3A65702",
    x"3A6536D",
    x"3A64FD9",
    x"3A64C45",
    x"3A648B2",
    x"3A64521",
    x"3A64190",
    x"3A63E00",
    x"3A63A71",
    x"3A636E3",
    x"3A63355",
    x"3A62FC9",
    x"3A62C3E",
    x"3A628B3",
    x"3A62529",
    x"3A621A0",
    x"3A61E18",
    x"3A61A91",
    x"3A6170B",
    x"3A61386",
    x"3A61001",
    x"3A60C7E",
    x"3A608FB",
    x"3A60579",
    x"3A601F8",
    x"3A5FE78",
    x"3A5FAF9",
    x"3A5F77B",
    x"3A5F3FD",
    x"3A5F081",
    x"3A5ED05",
    x"3A5E98A",
    x"3A5E610",
    x"3A5E297",
    x"3A5DF1F",
    x"3A5DBA8",
    x"3A5D831",
    x"3A5D4BC",
    x"3A5D147",
    x"3A5CDD3",
    x"3A5CA60",
    x"3A5C6EE",
    x"3A5C37C",
    x"3A5C00C",
    x"3A5BC9C",
    x"3A5B92E",
    x"3A5B5C0",
    x"3A5B253",
    x"3A5AEE7",
    x"3A5AB7B",
    x"3A5A811",
    x"3A5A4A7",
    x"3A5A13F",
    x"3A59DD7",
    x"3A59A70",
    x"3A5970A",
    x"3A593A4",
    x"3A59040",
    x"3A58CDC",
    x"3A58979",
    x"3A58617",
    x"3A582B6",
    x"3A57F56",
    x"3A57BF7",
    x"3A57898",
    x"3A5753A",
    x"3A571DD",
    x"3A56E81",
    x"3A56B26",
    x"3A567CC",
    x"3A56472",
    x"3A5611A",
    x"3A55DC2",
    x"3A55A6B",
    x"3A55714",
    x"3A553BF",
    x"3A5506B",
    x"3A54D17",
    x"3A549C4",
    x"3A54672",
    x"3A54321",
    x"3A53FD0",
    x"3A53C81",
    x"3A53932",
    x"3A535E4",
    x"3A53297",
    x"3A52F4B",
    x"3A52C00",
    x"3A528B5",
    x"3A5256B",
    x"3A52222",
    x"3A51EDA",
    x"3A51B93",
    x"3A5184C",
    x"3A51507",
    x"3A511C2",
    x"3A50E7E",
    x"3A50B3B",
    x"3A507F8",
    x"3A504B7",
    x"3A50176",
    x"3A4FE36",
    x"3A4FAF7",
    x"3A4F7B8",
    x"3A4F47B",
    x"3A4F13E",
    x"3A4EE02",
    x"3A4EAC7",
    x"3A4E78D",
    x"3A4E453",
    x"3A4E11B",
    x"3A4DDE3",
    x"3A4DAAC",
    x"3A4D776",
    x"3A4D440",
    x"3A4D10B",
    x"3A4CDD8",
    x"3A4CAA4",
    x"3A4C772",
    x"3A4C441",
    x"3A4C110",
    x"3A4BDE0",
    x"3A4BAB1",
    x"3A4B783",
    x"3A4B455",
    x"3A4B129",
    x"3A4ADFD",
    x"3A4AAD2",
    x"3A4A7A7",
    x"3A4A47E",
    x"3A4A155",
    x"3A49E2D",
    x"3A49B06",
    x"3A497E0",
    x"3A494BA",
    x"3A49195",
    x"3A48E71",
    x"3A48B4E",
    x"3A4882C",
    x"3A4850A",
    x"3A481E9",
    x"3A47EC9",
    x"3A47BAA",
    x"3A4788B",
    x"3A4756D",
    x"3A47251",
    x"3A46F34",
    x"3A46C19",
    x"3A468FE",
    x"3A465E4",
    x"3A462CB",
    x"3A45FB3",
    x"3A45C9B",
    x"3A45985",
    x"3A4566F",
    x"3A45359",
    x"3A45045",
    x"3A44D31",
    x"3A44A1E",
    x"3A4470C",
    x"3A443FB",
    x"3A440EA",
    x"3A43DDA",
    x"3A43ACB",
    x"3A437BD",
    x"3A434B0",
    x"3A431A3",
    x"3A42E97",
    x"3A42B8B",
    x"3A42881",
    x"3A42577",
    x"3A4226E",
    x"3A41F66",
    x"3A41C5E",
    x"3A41958",
    x"3A41652",
    x"3A4134D",
    x"3A41048",
    x"3A40D44",
    x"3A40A42",
    x"3A4073F",
    x"3A4043E",
    x"3A4013D",
    x"3A3FE3D",
    x"3A3FB3E",
    x"3A3F840",
    x"3A3F542",
    x"3A3F245",
    x"3A3EF49",
    x"3A3EC4D",
    x"3A3E953",
    x"3A3E659",
    x"3A3E360",
    x"3A3E067",
    x"3A3DD6F",
    x"3A3DA78",
    x"3A3D782",
    x"3A3D48D",
    x"3A3D198",
    x"3A3CEA4",
    x"3A3CBB0",
    x"3A3C8BE",
    x"3A3C5CC",
    x"3A3C2DB",
    x"3A3BFEB",
    x"3A3BCFB",
    x"3A3BA0C",
    x"3A3B71E",
    x"3A3B431",
    x"3A3B144",
    x"3A3AE58",
    x"3A3AB6D",
    x"3A3A882",
    x"3A3A599",
    x"3A3A2AF",
    x"3A39FC7",
    x"3A39CE0",
    x"3A399F9",
    x"3A39713",
    x"3A3942D",
    x"3A39149",
    x"3A38E65",
    x"3A38B81",
    x"3A3889F",
    x"3A385BD",
    x"3A382DC",
    x"3A37FFC",
    x"3A37D1C",
    x"3A37A3D",
    x"3A3775F",
    x"3A37481",
    x"3A371A5",
    x"3A36EC9",
    x"3A36BED",
    x"3A36913",
    x"3A36639",
    x"3A3635F",
    x"3A36087",
    x"3A35DAF",
    x"3A35AD8",
    x"3A35802",
    x"3A3552C",
    x"3A35257",
    x"3A34F83",
    x"3A34CAF",
    x"3A349DD",
    x"3A3470A",
    x"3A34439",
    x"3A34168",
    x"3A33E98",
    x"3A33BC9",
    x"3A338FA",
    x"3A3362D",
    x"3A3335F",
    x"3A33093",
    x"3A32DC7",
    x"3A32AFC",
    x"3A32832",
    x"3A32568",
    x"3A3229F",
    x"3A31FD7",
    x"3A31D0F",
    x"3A31A48",
    x"3A31782",
    x"3A314BC",
    x"3A311F7",
    x"3A30F33",
    x"3A30C70",
    x"3A309AD",
    x"3A306EB",
    x"3A3042A",
    x"3A30169",
    x"3A2FEA9",
    x"3A2FBEA",
    x"3A2F92B",
    x"3A2F66D",
    x"3A2F3B0",
    x"3A2F0F3",
    x"3A2EE37",
    x"3A2EB7C",
    x"3A2E8C2",
    x"3A2E608",
    x"3A2E34F",
    x"3A2E096",
    x"3A2DDDE",
    x"3A2DB27",
    x"3A2D871",
    x"3A2D5BB",
    x"3A2D306",
    x"3A2D051",
    x"3A2CD9E",
    x"3A2CAEB",
    x"3A2C838",
    x"3A2C586",
    x"3A2C2D5",
    x"3A2C025",
    x"3A2BD75",
    x"3A2BAC6",
    x"3A2B818",
    x"3A2B56A",
    x"3A2B2BD",
    x"3A2B011",
    x"3A2AD65",
    x"3A2AABA",
    x"3A2A810",
    x"3A2A566",
    x"3A2A2BD",
    x"3A2A015",
    x"3A29D6D",
    x"3A29AC6",
    x"3A29820",
    x"3A2957A",
    x"3A292D5",
    x"3A29031",
    x"3A28D8D",
    x"3A28AEA",
    x"3A28847",
    x"3A285A6",
    x"3A28305",
    x"3A28064",
    x"3A27DC4",
    x"3A27B25",
    x"3A27887",
    x"3A275E9",
    x"3A2734C",
    x"3A270AF",
    x"3A26E14",
    x"3A26B78",
    x"3A268DE",
    x"3A26644",
    x"3A263AB",
    x"3A26112",
    x"3A25E7A",
    x"3A25BE3",
    x"3A2594C",
    x"3A256B6",
    x"3A25421",
    x"3A2518C",
    x"3A24EF8",
    x"3A24C65",
    x"3A249D2",
    x"3A24740",
    x"3A244AE",
    x"3A2421D",
    x"3A23F8D",
    x"3A23CFE",
    x"3A23A6F",
    x"3A237E0",
    x"3A23553",
    x"3A232C6",
    x"3A23039",
    x"3A22DAE",
    x"3A22B22",
    x"3A22898",
    x"3A2260E",
    x"3A22385",
    x"3A220FC",
    x"3A21E74",
    x"3A21BED",
    x"3A21967",
    x"3A216E0",
    x"3A2145B",
    x"3A211D6",
    x"3A20F52",
    x"3A20CCF",
    x"3A20A4C",
    x"3A207C9",
    x"3A20548",
    x"3A202C7",
    x"3A20046",
    x"3A1FDC7",
    x"3A1FB48",
    x"3A1F8C9",
    x"3A1F64B",
    x"3A1F3CE",
    x"3A1F151",
    x"3A1EED5",
    x"3A1EC5A",
    x"3A1E9DF",
    x"3A1E765",
    x"3A1E4EB",
    x"3A1E272",
    x"3A1DFFA",
    x"3A1DD82",
    x"3A1DB0B",
    x"3A1D895",
    x"3A1D61F",
    x"3A1D3AA",
    x"3A1D135",
    x"3A1CEC1",
    x"3A1CC4E",
    x"3A1C9DB",
    x"3A1C769",
    x"3A1C4F7",
    x"3A1C286",
    x"3A1C016",
    x"3A1BDA6",
    x"3A1BB37",
    x"3A1B8C9",
    x"3A1B65B",
    x"3A1B3EE",
    x"3A1B181",
    x"3A1AF15",
    x"3A1ACA9",
    x"3A1AA3F",
    x"3A1A7D4",
    x"3A1A56B",
    x"3A1A302",
    x"3A1A099",
    x"3A19E31",
    x"3A19BCA",
    x"3A19963",
    x"3A196FD",
    x"3A19498",
    x"3A19233",
    x"3A18FCF",
    x"3A18D6B",
    x"3A18B08",
    x"3A188A6",
    x"3A18644",
    x"3A183E3",
    x"3A18182",
    x"3A17F22",
    x"3A17CC2",
    x"3A17A63",
    x"3A17805",
    x"3A175A7",
    x"3A1734A",
    x"3A170EE",
    x"3A16E92",
    x"3A16C36",
    x"3A169DC",
    x"3A16782",
    x"3A16528",
    x"3A162CF",
    x"3A16077",
    x"3A15E1F",
    x"3A15BC7",
    x"3A15971",
    x"3A1571B",
    x"3A154C5",
    x"3A15270",
    x"3A1501C",
    x"3A14DC8",
    x"3A14B75",
    x"3A14923",
    x"3A146D1",
    x"3A1447F",
    x"3A1422E",
    x"3A13FDE",
    x"3A13D8E",
    x"3A13B3F",
    x"3A138F1",
    x"3A136A3",
    x"3A13455",
    x"3A13209",
    x"3A12FBC",
    x"3A12D71",
    x"3A12B26",
    x"3A128DB",
    x"3A12691",
    x"3A12448",
    x"3A121FF",
    x"3A11FB7",
    x"3A11D6F",
    x"3A11B28",
    x"3A118E2",
    x"3A1169C",
    x"3A11456",
    x"3A11212",
    x"3A10FCD",
    x"3A10D8A",
    x"3A10B47",
    x"3A10904",
    x"3A106C2",
    x"3A10481",
    x"3A10240",
    x"3A10000",
    x"3A0FDC0",
    x"3A0FB81",
    x"3A0F942",
    x"3A0F704",
    x"3A0F4C7",
    x"3A0F28A",
    x"3A0F04D",
    x"3A0EE11",
    x"3A0EBD6",
    x"3A0E99C",
    x"3A0E761",
    x"3A0E528",
    x"3A0E2EF",
    x"3A0E0B6",
    x"3A0DE7F",
    x"3A0DC47",
    x"3A0DA10",
    x"3A0D7DA",
    x"3A0D5A4",
    x"3A0D36F",
    x"3A0D13B",
    x"3A0CF07",
    x"3A0CCD3",
    x"3A0CAA0",
    x"3A0C86E",
    x"3A0C63C",
    x"3A0C40B",
    x"3A0C1DA",
    x"3A0BFAA",
    x"3A0BD7A",
    x"3A0BB4B",
    x"3A0B91D",
    x"3A0B6EF",
    x"3A0B4C1",
    x"3A0B294",
    x"3A0B068",
    x"3A0AE3C",
    x"3A0AC11",
    x"3A0A9E6",
    x"3A0A7BC",
    x"3A0A592",
    x"3A0A369",
    x"3A0A140",
    x"3A09F18",
    x"3A09CF1",
    x"3A09ACA",
    x"3A098A3",
    x"3A0967E",
    x"3A09458",
    x"3A09233",
    x"3A0900F",
    x"3A08DEB",
    x"3A08BC8",
    x"3A089A5",
    x"3A08783",
    x"3A08562",
    x"3A08341",
    x"3A08120",
    x"3A07F00",
    x"3A07CE1",
    x"3A07AC2",
    x"3A078A3",
    x"3A07685",
    x"3A07468",
    x"3A0724B",
    x"3A0702F",
    x"3A06E13",
    x"3A06BF8",
    x"3A069DD",
    x"3A067C3",
    x"3A065A9",
    x"3A06390",
    x"3A06177",
    x"3A05F5F",
    x"3A05D48",
    x"3A05B31",
    x"3A0591A",
    x"3A05704",
    x"3A054EF",
    x"3A052DA",
    x"3A050C5",
    x"3A04EB1",
    x"3A04C9E",
    x"3A04A8B",
    x"3A04878",
    x"3A04667",
    x"3A04455",
    x"3A04244",
    x"3A04034",
    x"3A03E24",
    x"3A03C15",
    x"3A03A06",
    x"3A037F8",
    x"3A035EA",
    x"3A033DD",
    x"3A031D0",
    x"3A02FC4",
    x"3A02DB9",
    x"3A02BAD",
    x"3A029A3",
    x"3A02799",
    x"3A0258F",
    x"3A02386",
    x"3A0217D",
    x"3A01F75",
    x"3A01D6D",
    x"3A01B66",
    x"3A01960",
    x"3A0175A",
    x"3A01554",
    x"3A0134F",
    x"3A0114A",
    x"3A00F46",
    x"3A00D43",
    x"3A00B40",
    x"3A0093D",
    x"3A0073B",
    x"3A00539",
    x"3A00338",
    x"3A00138",
    x"39FFE70",
    x"39FFA71",
    x"39FF673",
    x"39FF276",
    x"39FEE7A",
    x"39FEA7F",
    x"39FE684",
    x"39FE28B",
    x"39FDE93",
    x"39FDA9C",
    x"39FD6A6",
    x"39FD2B1",
    x"39FCEBC",
    x"39FCAC9",
    x"39FC6D7",
    x"39FC2E6",
    x"39FBEF6",
    x"39FBB06",
    x"39FB718",
    x"39FB32B",
    x"39FAF3F",
    x"39FAB53",
    x"39FA769",
    x"39FA37F",
    x"39F9F97",
    x"39F9BB0",
    x"39F97C9",
    x"39F93E4",
    x"39F8FFF",
    x"39F8C1C",
    x"39F8839",
    x"39F8458",
    x"39F8077",
    x"39F7C97",
    x"39F78B9",
    x"39F74DB",
    x"39F70FE",
    x"39F6D23",
    x"39F6948",
    x"39F656E",
    x"39F6195",
    x"39F5DBD",
    x"39F59E6",
    x"39F5610",
    x"39F523B",
    x"39F4E67",
    x"39F4A94",
    x"39F46C2",
    x"39F42F1",
    x"39F3F20",
    x"39F3B51",
    x"39F3783",
    x"39F33B5",
    x"39F2FE9",
    x"39F2C1D",
    x"39F2853",
    x"39F2489",
    x"39F20C0",
    x"39F1CF9",
    x"39F1932",
    x"39F156C",
    x"39F11A7",
    x"39F0DE3",
    x"39F0A20",
    x"39F065E",
    x"39F029D",
    x"39EFEDD",
    x"39EFB1E",
    x"39EF75F",
    x"39EF3A2",
    x"39EEFE6",
    x"39EEC2A",
    x"39EE870",
    x"39EE4B6",
    x"39EE0FD",
    x"39EDD45",
    x"39ED98F",
    x"39ED5D9",
    x"39ED224",
    x"39ECE70",
    x"39ECABC",
    x"39EC70A",
    x"39EC359",
    x"39EBFA8",
    x"39EBBF9",
    x"39EB84A",
    x"39EB49D",
    x"39EB0F0",
    x"39EAD44",
    x"39EA99A",
    x"39EA5F0",
    x"39EA247",
    x"39E9E9E",
    x"39E9AF7",
    x"39E9751",
    x"39E93AC",
    x"39E9007",
    x"39E8C64",
    x"39E88C1",
    x"39E851F",
    x"39E817E",
    x"39E7DDE",
    x"39E7A3F",
    x"39E76A1",
    x"39E7304",
    x"39E6F68",
    x"39E6BCC",
    x"39E6832",
    x"39E6498",
    x"39E6100",
    x"39E5D68",
    x"39E59D1",
    x"39E563B",
    x"39E52A6",
    x"39E4F12",
    x"39E4B7E",
    x"39E47EC",
    x"39E445A",
    x"39E40CA",
    x"39E3D3A",
    x"39E39AB",
    x"39E361D",
    x"39E3290",
    x"39E2F04",
    x"39E2B78",
    x"39E27EE",
    x"39E2465",
    x"39E20DC",
    x"39E1D54",
    x"39E19CD",
    x"39E1647",
    x"39E12C2",
    x"39E0F3E",
    x"39E0BBA",
    x"39E0838",
    x"39E04B6",
    x"39E0136",
    x"39DFDB6",
    x"39DFA37",
    x"39DF6B9",
    x"39DF33B",
    x"39DEFBF",
    x"39DEC43",
    x"39DE8C9",
    x"39DE54F",
    x"39DE1D6",
    x"39DDE5E",
    x"39DDAE7",
    x"39DD771",
    x"39DD3FB",
    x"39DD087",
    x"39DCD13",
    x"39DC9A0",
    x"39DC62E",
    x"39DC2BD",
    x"39DBF4D",
    x"39DBBDD",
    x"39DB86F",
    x"39DB501",
    x"39DB194",
    x"39DAE28",
    x"39DAABD",
    x"39DA753",
    x"39DA3EA",
    x"39DA081",
    x"39D9D19",
    x"39D99B3",
    x"39D964D",
    x"39D92E7",
    x"39D8F83",
    x"39D8C20",
    x"39D88BD",
    x"39D855B",
    x"39D81FA",
    x"39D7E9A",
    x"39D7B3B",
    x"39D77DD",
    x"39D747F",
    x"39D7122",
    x"39D6DC7",
    x"39D6A6C",
    x"39D6711",
    x"39D63B8",
    x"39D605F",
    x"39D5D08",
    x"39D59B1",
    x"39D565B",
    x"39D5306",
    x"39D4FB1",
    x"39D4C5E",
    x"39D490B",
    x"39D45B9",
    x"39D4268",
    x"39D3F18",
    x"39D3BC9",
    x"39D387A",
    x"39D352D",
    x"39D31E0",
    x"39D2E94",
    x"39D2B48",
    x"39D27FE",
    x"39D24B4",
    x"39D216C",
    x"39D1E24",
    x"39D1ADD",
    x"39D1796",
    x"39D1451",
    x"39D110C",
    x"39D0DC8",
    x"39D0A85",
    x"39D0743",
    x"39D0402",
    x"39D00C1",
    x"39CFD81",
    x"39CFA42",
    x"39CF704",
    x"39CF3C7",
    x"39CF08A",
    x"39CED4F",
    x"39CEA14",
    x"39CE6D9",
    x"39CE3A0",
    x"39CE068",
    x"39CDD30",
    x"39CD9F9",
    x"39CD6C3",
    x"39CD38E",
    x"39CD059",
    x"39CCD25",
    x"39CC9F3",
    x"39CC6C1",
    x"39CC38F",
    x"39CC05F",
    x"39CBD2F",
    x"39CBA00",
    x"39CB6D2",
    x"39CB3A5",
    x"39CB078",
    x"39CAD4C",
    x"39CAA22",
    x"39CA6F7",
    x"39CA3CE",
    x"39CA0A6",
    x"39C9D7E",
    x"39C9A57",
    x"39C9731",
    x"39C940B",
    x"39C90E7",
    x"39C8DC3",
    x"39C8AA0",
    x"39C877D",
    x"39C845C",
    x"39C813B",
    x"39C7E1B",
    x"39C7AFC",
    x"39C77DE",
    x"39C74C0",
    x"39C71A3",
    x"39C6E87",
    x"39C6B6C",
    x"39C6852",
    x"39C6538",
    x"39C621F",
    x"39C5F07",
    x"39C5BF0",
    x"39C58D9",
    x"39C55C3",
    x"39C52AE",
    x"39C4F9A",
    x"39C4C86",
    x"39C4974",
    x"39C4662",
    x"39C4350",
    x"39C4040",
    x"39C3D30",
    x"39C3A21",
    x"39C3713",
    x"39C3406",
    x"39C30F9",
    x"39C2DED",
    x"39C2AE2",
    x"39C27D8",
    x"39C24CE",
    x"39C21C5",
    x"39C1EBD",
    x"39C1BB6",
    x"39C18B0",
    x"39C15AA",
    x"39C12A5",
    x"39C0FA0",
    x"39C0C9D",
    x"39C099A",
    x"39C0698",
    x"39C0397",
    x"39C0096",
    x"39BFD97",
    x"39BFA97",
    x"39BF799",
    x"39BF49C",
    x"39BF19F",
    x"39BEEA3",
    x"39BEBA8",
    x"39BE8AD",
    x"39BE5B3",
    x"39BE2BA",
    x"39BDFC2",
    x"39BDCCA",
    x"39BD9D3",
    x"39BD6DD",
    x"39BD3E8",
    x"39BD0F3",
    x"39BCE00",
    x"39BCB0C",
    x"39BC81A",
    x"39BC528",
    x"39BC237",
    x"39BBF47",
    x"39BBC58",
    x"39BB969",
    x"39BB67B",
    x"39BB38E",
    x"39BB0A1",
    x"39BADB6",
    x"39BAACB",
    x"39BA7E0",
    x"39BA4F7",
    x"39BA20E",
    x"39B9F26",
    x"39B9C3E",
    x"39B9957",
    x"39B9671",
    x"39B938C",
    x"39B90A8",
    x"39B8DC4",
    x"39B8AE1",
    x"39B87FE",
    x"39B851D",
    x"39B823C",
    x"39B7F5C",
    x"39B7C7C",
    x"39B799D",
    x"39B76BF",
    x"39B73E2",
    x"39B7105",
    x"39B6E2A",
    x"39B6B4E",
    x"39B6874",
    x"39B659A",
    x"39B62C1",
    x"39B5FE9",
    x"39B5D11",
    x"39B5A3A",
    x"39B5764",
    x"39B548F",
    x"39B51BA",
    x"39B4EE6",
    x"39B4C12",
    x"39B4940",
    x"39B466E",
    x"39B439C",
    x"39B40CC",
    x"39B3DFC",
    x"39B3B2D",
    x"39B385E",
    x"39B3591",
    x"39B32C4",
    x"39B2FF7",
    x"39B2D2C",
    x"39B2A61",
    x"39B2796",
    x"39B24CD",
    x"39B2204",
    x"39B1F3C",
    x"39B1C74",
    x"39B19AE",
    x"39B16E8",
    x"39B1422",
    x"39B115E",
    x"39B0E9A",
    x"39B0BD6",
    x"39B0914",
    x"39B0652",
    x"39B0390",
    x"39B00D0",
    x"39AFE10",
    x"39AFB51",
    x"39AF892",
    x"39AF5D5",
    x"39AF317",
    x"39AF05B",
    x"39AED9F",
    x"39AEAE4",
    x"39AE82A",
    x"39AE570",
    x"39AE2B7",
    x"39ADFFF",
    x"39ADD47",
    x"39ADA90",
    x"39AD7DA",
    x"39AD524",
    x"39AD26F",
    x"39ACFBB",
    x"39ACD07",
    x"39ACA54",
    x"39AC7A2",
    x"39AC4F1",
    x"39AC240",
    x"39ABF90",
    x"39ABCE0",
    x"39ABA31",
    x"39AB783",
    x"39AB4D5",
    x"39AB228",
    x"39AAF7C",
    x"39AACD1",
    x"39AAA26",
    x"39AA77C",
    x"39AA4D2",
    x"39AA229",
    x"39A9F81",
    x"39A9CD9",
    x"39A9A33",
    x"39A978C",
    x"39A94E7",
    x"39A9242",
    x"39A8F9E",
    x"39A8CFA",
    x"39A8A57",
    x"39A87B5",
    x"39A8513",
    x"39A8272",
    x"39A7FD2",
    x"39A7D32",
    x"39A7A94",
    x"39A77F5",
    x"39A7558",
    x"39A72BB",
    x"39A701E",
    x"39A6D82",
    x"39A6AE7",
    x"39A684D",
    x"39A65B3",
    x"39A631A",
    x"39A6082",
    x"39A5DEA",
    x"39A5B53",
    x"39A58BC",
    x"39A5626",
    x"39A5391",
    x"39A50FD",
    x"39A4E69",
    x"39A4BD5",
    x"39A4943",
    x"39A46B1",
    x"39A441F",
    x"39A418F",
    x"39A3EFF",
    x"39A3C6F",
    x"39A39E0",
    x"39A3752",
    x"39A34C5",
    x"39A3238",
    x"39A2FAC",
    x"39A2D20",
    x"39A2A95",
    x"39A280B",
    x"39A2581",
    x"39A22F8",
    x"39A2070",
    x"39A1DE8",
    x"39A1B61",
    x"39A18DA",
    x"39A1654",
    x"39A13CF",
    x"39A114A",
    x"39A0EC6",
    x"39A0C43",
    x"39A09C0",
    x"39A073E",
    x"39A04BD",
    x"39A023C",
    x"399FFBB",
    x"399FD3C",
    x"399FABD",
    x"399F83E",
    x"399F5C1",
    x"399F344",
    x"399F0C7",
    x"399EE4B",
    x"399EBD0",
    x"399E955",
    x"399E6DB",
    x"399E462",
    x"399E1E9",
    x"399DF71",
    x"399DCF9",
    x"399DA82",
    x"399D80C",
    x"399D596",
    x"399D321",
    x"399D0AD",
    x"399CE39",
    x"399CBC6",
    x"399C953",
    x"399C6E1",
    x"399C470",
    x"399C1FF",
    x"399BF8F",
    x"399BD1F",
    x"399BAB0",
    x"399B842",
    x"399B5D4",
    x"399B367",
    x"399B0FA",
    x"399AE8E",
    x"399AC23",
    x"399A9B8",
    x"399A74E",
    x"399A4E5",
    x"399A27C",
    x"399A013",
    x"3999DAC",
    x"3999B44",
    x"39998DE",
    x"3999678",
    x"3999413",
    x"39991AE",
    x"3998F4A",
    x"3998CE6",
    x"3998A83",
    x"3998821",
    x"39985BF",
    x"399835E",
    x"39980FE",
    x"3997E9E",
    x"3997C3E",
    x"39979E0",
    x"3997781",
    x"3997524",
    x"39972C7",
    x"399706A",
    x"3996E0F",
    x"3996BB3",
    x"3996959",
    x"39966FF",
    x"39964A5",
    x"399624C",
    x"3995FF4",
    x"3995D9C",
    x"3995B45",
    x"39958EF",
    x"3995699",
    x"3995444",
    x"39951EF",
    x"3994F9B",
    x"3994D47",
    x"3994AF4",
    x"39948A1",
    x"3994650",
    x"39943FE",
    x"39941AE",
    x"3993F5D",
    x"3993D0E",
    x"3993ABF",
    x"3993871",
    x"3993623",
    x"39933D5",
    x"3993189",
    x"3992F3D",
    x"3992CF1",
    x"3992AA6",
    x"399285C",
    x"3992612",
    x"39923C9",
    x"3992180",
    x"3991F38",
    x"3991CF1",
    x"3991AAA",
    x"3991863",
    x"399161D",
    x"39913D8",
    x"3991193",
    x"3990F4F",
    x"3990D0C",
    x"3990AC9",
    x"3990886",
    x"3990645",
    x"3990403",
    x"39901C3",
    x"398FF82",
    x"398FD43",
    x"398FB04",
    x"398F8C5",
    x"398F687",
    x"398F44A",
    x"398F20D",
    x"398EFD1",
    x"398ED95",
    x"398EB5A",
    x"398E920",
    x"398E6E6",
    x"398E4AC",
    x"398E273",
    x"398E03B",
    x"398DE03",
    x"398DBCC",
    x"398D995",
    x"398D75F",
    x"398D52A",
    x"398D2F5",
    x"398D0C0",
    x"398CE8C",
    x"398CC59",
    x"398CA26",
    x"398C7F4",
    x"398C5C2",
    x"398C391",
    x"398C160",
    x"398BF30",
    x"398BD01",
    x"398BAD2",
    x"398B8A3",
    x"398B675",
    x"398B448",
    x"398B21B",
    x"398AFEF",
    x"398ADC3",
    x"398AB98",
    x"398A96D",
    x"398A743",
    x"398A51A",
    x"398A2F1",
    x"398A0C8",
    x"3989EA0",
    x"3989C79",
    x"3989A52",
    x"398982C",
    x"3989606",
    x"39893E1",
    x"39891BC",
    x"3988F98",
    x"3988D74",
    x"3988B51",
    x"398892F",
    x"398870D",
    x"39884EB",
    x"39882CA",
    x"39880AA",
    x"3987E8A",
    x"3987C6B",
    x"3987A4C",
    x"398782D",
    x"3987610",
    x"39873F2",
    x"39871D6",
    x"3986FB9",
    x"3986D9E",
    x"3986B83",
    x"3986968",
    x"398674E",
    x"3986534",
    x"398631B",
    x"3986103",
    x"3985EEB",
    x"3985CD3",
    x"3985ABC",
    x"39858A6",
    x"3985690",
    x"398547B",
    x"3985266",
    x"3985051",
    x"3984E3E",
    x"3984C2A",
    x"3984A18",
    x"3984805",
    x"39845F4",
    x"39843E2",
    x"39841D2",
    x"3983FC1",
    x"3983DB2",
    x"3983BA3",
    x"3983994",
    x"3983786",
    x"3983578",
    x"398336B",
    x"398315E",
    x"3982F52",
    x"3982D47",
    x"3982B3C",
    x"3982931",
    x"3982727",
    x"398251E",
    x"3982315",
    x"398210C",
    x"3981F04",
    x"3981CFD",
    x"3981AF6",
    x"39818EF",
    x"39816E9",
    x"39814E4",
    x"39812DF",
    x"39810DA",
    x"3980ED6",
    x"3980CD3",
    x"3980AD0",
    x"39808CD",
    x"39806CB",
    x"39804CA",
    x"39802C9",
    x"39800C9",
    x"397FD92",
    x"397F993",
    x"397F595",
    x"397F198",
    x"397ED9C",
    x"397E9A1",
    x"397E5A7",
    x"397E1AE",
    x"397DDB6",
    x"397D9C0",
    x"397D5CA",
    x"397D1D5",
    x"397CDE1",
    x"397C9EE",
    x"397C5FC",
    x"397C20B",
    x"397BE1B",
    x"397BA2C",
    x"397B63E",
    x"397B251",
    x"397AE64",
    x"397AA79",
    x"397A68F",
    x"397A2A6",
    x"3979EBE",
    x"3979AD7",
    x"39796F0",
    x"397930B",
    x"3978F27",
    x"3978B44",
    x"3978761",
    x"3978380",
    x"3977FA0",
    x"3977BC0",
    x"39777E2",
    x"3977404",
    x"3977028",
    x"3976C4C",
    x"3976871",
    x"3976498",
    x"39760BF",
    x"3975CE7",
    x"3975911",
    x"397553B",
    x"3975166",
    x"3974D92",
    x"39749BF",
    x"39745ED",
    x"397421C",
    x"3973E4C",
    x"3973A7D",
    x"39736AF",
    x"39732E2",
    x"3972F16",
    x"3972B4A",
    x"3972780",
    x"39723B7",
    x"3971FEE",
    x"3971C27",
    x"3971860",
    x"397149A",
    x"39710D6",
    x"3970D12",
    x"397094F",
    x"397058D",
    x"39701CC",
    x"396FE0C",
    x"396FA4D",
    x"396F68F",
    x"396F2D2",
    x"396EF16",
    x"396EB5B",
    x"396E7A0",
    x"396E3E7",
    x"396E02E",
    x"396DC77",
    x"396D8C0",
    x"396D50A",
    x"396D156",
    x"396CDA2",
    x"396C9EF",
    x"396C63D",
    x"396C28C",
    x"396BEDB",
    x"396BB2C",
    x"396B77E",
    x"396B3D0",
    x"396B024",
    x"396AC78",
    x"396A8CE",
    x"396A524",
    x"396A17B",
    x"3969DD3",
    x"3969A2C",
    x"3969686",
    x"39692E1",
    x"3968F3D",
    x"3968B99",
    x"39687F7",
    x"3968455",
    x"39680B5",
    x"3967D15",
    x"3967976",
    x"39675D8",
    x"396723B",
    x"3966E9F",
    x"3966B04",
    x"396676A",
    x"39663D0",
    x"3966038",
    x"3965CA0",
    x"3965909",
    x"3965574",
    x"39651DF",
    x"3964E4B",
    x"3964AB8",
    x"3964725",
    x"3964394",
    x"3964003",
    x"3963C74",
    x"39638E5",
    x"3963557",
    x"39631CB",
    x"3962E3F",
    x"3962AB3",
    x"3962729",
    x"39623A0",
    x"3962017",
    x"3961C90",
    x"3961909",
    x"3961583",
    x"39611FE",
    x"3960E7A",
    x"3960AF7",
    x"3960775",
    x"39603F3",
    x"3960073",
    x"395FCF3",
    x"395F974",
    x"395F5F6",
    x"395F279",
    x"395EEFD",
    x"395EB82",
    x"395E807",
    x"395E48E",
    x"395E115",
    x"395DD9D",
    x"395DA26",
    x"395D6B0",
    x"395D33B",
    x"395CFC7",
    x"395CC53",
    x"395C8E0",
    x"395C56F",
    x"395C1FE",
    x"395BE8E",
    x"395BB1E",
    x"395B7B0",
    x"395B443",
    x"395B0D6",
    x"395AD6A",
    x"395A9FF",
    x"395A695",
    x"395A32C",
    x"3959FC4",
    x"3959C5C",
    x"39598F5",
    x"3959590",
    x"395922B",
    x"3958EC7",
    x"3958B63",
    x"3958801",
    x"395849F",
    x"395813F",
    x"3957DDF",
    x"3957A80",
    x"3957721",
    x"39573C4",
    x"3957068",
    x"3956D0C",
    x"39569B1",
    x"3956657",
    x"39562FE",
    x"3955FA6",
    x"3955C4E",
    x"39558F7",
    x"39555A2",
    x"395524D",
    x"3954EF8",
    x"3954BA5",
    x"3954853",
    x"3954501",
    x"39541B0",
    x"3953E60",
    x"3953B11",
    x"39537C3",
    x"3953475",
    x"3953128",
    x"3952DDC",
    x"3952A91",
    x"3952747",
    x"39523FE",
    x"39520B5",
    x"3951D6D",
    x"3951A26",
    x"39516E0",
    x"395139B",
    x"3951056",
    x"3950D13",
    x"39509D0",
    x"395068E",
    x"395034D",
    x"395000C",
    x"394FCCD",
    x"394F98E",
    x"394F650",
    x"394F313",
    x"394EFD6",
    x"394EC9B",
    x"394E960",
    x"394E626",
    x"394E2ED",
    x"394DFB5",
    x"394DC7D",
    x"394D946",
    x"394D610",
    x"394D2DB",
    x"394CFA7",
    x"394CC73",
    x"394C941",
    x"394C60F",
    x"394C2DE",
    x"394BFAD",
    x"394BC7E",
    x"394B94F",
    x"394B621",
    x"394B2F4",
    x"394AFC8",
    x"394AC9C",
    x"394A971",
    x"394A648",
    x"394A31E",
    x"3949FF6",
    x"3949CCE",
    x"39499A8",
    x"3949682",
    x"394935C",
    x"3949038",
    x"3948D14",
    x"39489F1",
    x"39486CF",
    x"39483AE",
    x"394808D",
    x"3947D6E",
    x"3947A4F",
    x"3947730",
    x"3947413",
    x"39470F6",
    x"3946DDB",
    x"3946ABF",
    x"39467A5",
    x"394648C",
    x"3946173",
    x"3945E5B",
    x"3945B44",
    x"394582D",
    x"3945518",
    x"3945203",
    x"3944EEF",
    x"3944BDB",
    x"39448C9",
    x"39445B7",
    x"39442A6",
    x"3943F96",
    x"3943C86",
    x"3943977",
    x"3943669",
    x"394335C",
    x"3943050",
    x"3942D44",
    x"3942A39",
    x"394272F",
    x"3942425",
    x"394211D",
    x"3941E15",
    x"3941B0E",
    x"3941807",
    x"3941502",
    x"39411FD",
    x"3940EF9",
    x"3940BF5",
    x"39408F3",
    x"39405F1",
    x"39402F0",
    x"393FFEF",
    x"393FCF0",
    x"393F9F1",
    x"393F6F3",
    x"393F3F5",
    x"393F0F9",
    x"393EDFD",
    x"393EB02",
    x"393E807",
    x"393E50E",
    x"393E215",
    x"393DF1D",
    x"393DC25",
    x"393D92F",
    x"393D639",
    x"393D344",
    x"393D04F",
    x"393CD5B",
    x"393CA68",
    x"393C776",
    x"393C485",
    x"393C194",
    x"393BEA4",
    x"393BBB5",
    x"393B8C6",
    x"393B5D8",
    x"393B2EB",
    x"393AFFF",
    x"393AD13",
    x"393AA28",
    x"393A73E",
    x"393A455",
    x"393A16C",
    x"3939E84",
    x"3939B9D",
    x"39398B6",
    x"39395D0",
    x"39392EB",
    x"3939007",
    x"3938D23",
    x"3938A40",
    x"393875E",
    x"393847D",
    x"393819C",
    x"3937EBC",
    x"3937BDC",
    x"39378FE",
    x"3937620",
    x"3937343",
    x"3937066",
    x"3936D8B",
    x"3936AB0",
    x"39367D5",
    x"39364FC",
    x"3936223",
    x"3935F4B",
    x"3935C73",
    x"393599C",
    x"39356C6",
    x"39353F1",
    x"393511C",
    x"3934E48",
    x"3934B75",
    x"39348A3",
    x"39345D1",
    x"3934300",
    x"393402F",
    x"3933D60",
    x"3933A91",
    x"39337C2",
    x"39334F5",
    x"3933228",
    x"3932F5C",
    x"3932C90",
    x"39329C5",
    x"39326FB",
    x"3932432",
    x"3932169",
    x"3931EA1",
    x"3931BDA",
    x"3931913",
    x"393164D",
    x"3931388",
    x"39310C4",
    x"3930E00",
    x"3930B3D",
    x"393087A",
    x"39305B8",
    x"39302F7",
    x"3930037",
    x"392FD77",
    x"392FAB8",
    x"392F7FA",
    x"392F53C",
    x"392F27F",
    x"392EFC3",
    x"392ED07",
    x"392EA4C",
    x"392E792",
    x"392E4D9",
    x"392E220",
    x"392DF68",
    x"392DCB0",
    x"392D9F9",
    x"392D743",
    x"392D48E",
    x"392D1D9",
    x"392CF25",
    x"392CC71",
    x"392C9BE",
    x"392C70C",
    x"392C45B",
    x"392C1AA",
    x"392BEFA",
    x"392BC4B",
    x"392B99C",
    x"392B6EE",
    x"392B440",
    x"392B194",
    x"392AEE8",
    x"392AC3C",
    x"392A992",
    x"392A6E7",
    x"392A43E",
    x"392A195",
    x"3929EED",
    x"3929C46",
    x"392999F",
    x"39296F9",
    x"3929454",
    x"39291AF",
    x"3928F0B",
    x"3928C67",
    x"39289C5",
    x"3928723",
    x"3928481",
    x"39281E0",
    x"3927F40",
    x"3927CA1",
    x"3927A02",
    x"3927764",
    x"39274C6",
    x"3927229",
    x"3926F8D",
    x"3926CF1",
    x"3926A57",
    x"39267BC",
    x"3926523",
    x"392628A",
    x"3925FF1",
    x"3925D5A",
    x"3925AC3",
    x"392582C",
    x"3925597",
    x"3925302",
    x"392506D",
    x"3924DD9",
    x"3924B46",
    x"39248B4",
    x"3924622",
    x"3924391",
    x"3924100",
    x"3923E70",
    x"3923BE1",
    x"3923952",
    x"39236C4",
    x"3923437",
    x"39231AA",
    x"3922F1E",
    x"3922C93",
    x"3922A08",
    x"392277E",
    x"39224F4",
    x"392226B",
    x"3921FE3",
    x"3921D5B",
    x"3921AD4",
    x"392184E",
    x"39215C8",
    x"3921343",
    x"39210BE",
    x"3920E3A",
    x"3920BB7",
    x"3920935",
    x"39206B3",
    x"3920431",
    x"39201B0",
    x"391FF30",
    x"391FCB1",
    x"391FA32",
    x"391F7B4",
    x"391F536",
    x"391F2B9",
    x"391F03D",
    x"391EDC1",
    x"391EB46",
    x"391E8CB",
    x"391E652",
    x"391E3D8",
    x"391E160",
    x"391DEE8",
    x"391DC70",
    x"391D9F9",
    x"391D783",
    x"391D50E",
    x"391D299",
    x"391D024",
    x"391CDB1",
    x"391CB3D",
    x"391C8CB",
    x"391C659",
    x"391C3E8",
    x"391C177",
    x"391BF07",
    x"391BC98",
    x"391BA29",
    x"391B7BB",
    x"391B54D",
    x"391B2E0",
    x"391B073",
    x"391AE08",
    x"391AB9C",
    x"391A932",
    x"391A6C8",
    x"391A45E",
    x"391A1F6",
    x"3919F8D",
    x"3919D26",
    x"3919ABF",
    x"3919858",
    x"39195F3",
    x"391938E",
    x"3919129",
    x"3918EC5",
    x"3918C62",
    x"39189FF",
    x"391879D",
    x"391853B",
    x"39182DA",
    x"391807A",
    x"3917E1A",
    x"3917BBA",
    x"391795C",
    x"39176FE",
    x"39174A0",
    x"3917243",
    x"3916FE7",
    x"3916D8C",
    x"3916B30",
    x"39168D6",
    x"391667C",
    x"3916423",
    x"39161CA",
    x"3915F72",
    x"3915D1A",
    x"3915AC3",
    x"391586D",
    x"3915617",
    x"39153C2",
    x"391516D",
    x"3914F19",
    x"3914CC6",
    x"3914A73",
    x"3914820",
    x"39145CF",
    x"391437D",
    x"391412D",
    x"3913EDD",
    x"3913C8D",
    x"3913A3F",
    x"39137F0",
    x"39135A3",
    x"3913355",
    x"3913109",
    x"3912EBD",
    x"3912C72",
    x"3912A27",
    x"39127DD",
    x"3912593",
    x"391234A",
    x"3912101",
    x"3911EB9",
    x"3911C72",
    x"3911A2B",
    x"39117E5",
    x"391159F",
    x"391135A",
    x"3911115",
    x"3910ED1",
    x"3910C8E",
    x"3910A4B",
    x"3910809",
    x"39105C7",
    x"3910386",
    x"3910145",
    x"390FF05",
    x"390FCC6",
    x"390FA87",
    x"390F849",
    x"390F60B",
    x"390F3CE",
    x"390F191",
    x"390EF55",
    x"390ED19",
    x"390EADE",
    x"390E8A4",
    x"390E66A",
    x"390E431",
    x"390E1F8",
    x"390DFC0",
    x"390DD88",
    x"390DB51",
    x"390D91A",
    x"390D6E4",
    x"390D4AF",
    x"390D27A",
    x"390D046",
    x"390CE12",
    x"390CBDF",
    x"390C9AC",
    x"390C77A",
    x"390C548",
    x"390C317",
    x"390C0E7",
    x"390BEB7",
    x"390BC87",
    x"390BA58",
    x"390B82A",
    x"390B5FC",
    x"390B3CF",
    x"390B1A2",
    x"390AF76",
    x"390AD4B",
    x"390AB20",
    x"390A8F5",
    x"390A6CB",
    x"390A4A2",
    x"390A279",
    x"390A050",
    x"3909E29",
    x"3909C01",
    x"39099DB",
    x"39097B4",
    x"390958F",
    x"390936A",
    x"3909145",
    x"3908F21",
    x"3908CFD",
    x"3908ADA",
    x"39088B8",
    x"3908696",
    x"3908475",
    x"3908254",
    x"3908034",
    x"3907E14",
    x"3907BF5",
    x"39079D6",
    x"39077B8",
    x"390759A",
    x"390737D",
    x"3907160",
    x"3906F44",
    x"3906D29",
    x"3906B0E",
    x"39068F3",
    x"39066D9",
    x"39064C0",
    x"39062A7",
    x"390608E",
    x"3905E76",
    x"3905C5F",
    x"3905A48",
    x"3905832",
    x"390561C",
    x"3905407",
    x"39051F2",
    x"3904FDE",
    x"3904DCA",
    x"3904BB7",
    x"39049A4",
    x"3904792",
    x"3904581",
    x"390436F",
    x"390415F",
    x"3903F4F",
    x"3903D3F",
    x"3903B30",
    x"3903922",
    x"3903714",
    x"3903506",
    x"39032F9",
    x"39030ED",
    x"3902EE1",
    x"3902CD5",
    x"3902ACA",
    x"39028C0",
    x"39026B6",
    x"39024AC",
    x"39022A3",
    x"390209B",
    x"3901E93",
    x"3901C8C",
    x"3901A85",
    x"390187E",
    x"3901679",
    x"3901473",
    x"390126E",
    x"390106A",
    x"3900E66",
    x"3900C63",
    x"3900A60",
    x"390085E",
    x"390065C",
    x"390045A",
    x"390025A",
    x"3900059",
    x"38FFCB3",
    x"38FF8B5",
    x"38FF4B7",
    x"38FF0BA",
    x"38FECBF",
    x"38FE8C4",
    x"38FE4CA",
    x"38FE0D2",
    x"38FDCDA",
    x"38FD8E3",
    x"38FD4ED",
    x"38FD0F9",
    x"38FCD05",
    x"38FC912",
    x"38FC520",
    x"38FC130",
    x"38FBD40",
    x"38FB951",
    x"38FB563",
    x"38FB176",
    x"38FAD8A",
    x"38FA99F",
    x"38FA5B6",
    x"38FA1CD",
    x"38F9DE5",
    x"38F99FE",
    x"38F9618",
    x"38F9233",
    x"38F8E4F",
    x"38F8A6B",
    x"38F8689",
    x"38F82A8",
    x"38F7EC8",
    x"38F7AE9",
    x"38F770B",
    x"38F732D",
    x"38F6F51",
    x"38F6B76",
    x"38F679B",
    x"38F63C2",
    x"38F5FE9",
    x"38F5C12",
    x"38F583B",
    x"38F5466",
    x"38F5091",
    x"38F4CBD",
    x"38F48EB",
    x"38F4519",
    x"38F4148",
    x"38F3D78",
    x"38F39A9",
    x"38F35DC",
    x"38F320F",
    x"38F2E43",
    x"38F2A77",
    x"38F26AD",
    x"38F22E4",
    x"38F1F1C",
    x"38F1B55",
    x"38F178E",
    x"38F13C9",
    x"38F1004",
    x"38F0C41",
    x"38F087E",
    x"38F04BC",
    x"38F00FC",
    x"38EFD3C",
    x"38EF97D",
    x"38EF5BF",
    x"38EF202",
    x"38EEE46",
    x"38EEA8B",
    x"38EE6D1",
    x"38EE318",
    x"38EDF5F",
    x"38EDBA8",
    x"38ED7F2",
    x"38ED43C",
    x"38ED087",
    x"38ECCD4",
    x"38EC921",
    x"38EC56F",
    x"38EC1BE",
    x"38EBE0E",
    x"38EBA5F",
    x"38EB6B1",
    x"38EB304",
    x"38EAF58",
    x"38EABAC",
    x"38EA802",
    x"38EA458",
    x"38EA0B0",
    x"38E9D08",
    x"38E9961",
    x"38E95BB",
    x"38E9216",
    x"38E8E72",
    x"38E8ACF",
    x"38E872D",
    x"38E838B",
    x"38E7FEB",
    x"38E7C4B",
    x"38E78AD",
    x"38E750F",
    x"38E7172",
    x"38E6DD6",
    x"38E6A3B",
    x"38E66A1",
    x"38E6308",
    x"38E5F70",
    x"38E5BD8",
    x"38E5842",
    x"38E54AC",
    x"38E5118",
    x"38E4D84",
    x"38E49F1",
    x"38E465F",
    x"38E42CE",
    x"38E3F3D",
    x"38E3BAE",
    x"38E381F",
    x"38E3492",
    x"38E3105",
    x"38E2D79",
    x"38E29EE",
    x"38E2664",
    x"38E22DB",
    x"38E1F53",
    x"38E1BCC",
    x"38E1845",
    x"38E14BF",
    x"38E113B",
    x"38E0DB7",
    x"38E0A34",
    x"38E06B2",
    x"38E0331",
    x"38DFFB0",
    x"38DFC31",
    x"38DF8B2",
    x"38DF534",
    x"38DF1B7",
    x"38DEE3B",
    x"38DEAC0",
    x"38DE746",
    x"38DE3CD",
    x"38DE054",
    x"38DDCDD",
    x"38DD966",
    x"38DD5F0",
    x"38DD27B",
    x"38DCF07",
    x"38DCB93",
    x"38DC821",
    x"38DC4AF",
    x"38DC13E",
    x"38DBDCF",
    x"38DBA60",
    x"38DB6F1",
    x"38DB384",
    x"38DB018",
    x"38DACAC",
    x"38DA941",
    x"38DA5D7",
    x"38DA26E",
    x"38D9F06",
    x"38D9B9F",
    x"38D9838",
    x"38D94D3",
    x"38D916E",
    x"38D8E0A",
    x"38D8AA7",
    x"38D8745",
    x"38D83E3",
    x"38D8083",
    x"38D7D23",
    x"38D79C4",
    x"38D7666",
    x"38D7309",
    x"38D6FAD",
    x"38D6C51",
    x"38D68F6",
    x"38D659D",
    x"38D6244",
    x"38D5EEC",
    x"38D5B94",
    x"38D583E",
    x"38D54E8",
    x"38D5193",
    x"38D4E3F",
    x"38D4AEC",
    x"38D479A",
    x"38D4448",
    x"38D40F8",
    x"38D3DA8",
    x"38D3A59",
    x"38D370B",
    x"38D33BD",
    x"38D3071",
    x"38D2D25",
    x"38D29DA",
    x"38D2690",
    x"38D2347",
    x"38D1FFF",
    x"38D1CB7",
    x"38D1970",
    x"38D162A",
    x"38D12E5",
    x"38D0FA1",
    x"38D0C5D",
    x"38D091B",
    x"38D05D9",
    x"38D0298",
    x"38CFF57",
    x"38CFC18",
    x"38CF8D9",
    x"38CF59C",
    x"38CF25F",
    x"38CEF22",
    x"38CEBE7",
    x"38CE8AC",
    x"38CE573",
    x"38CE23A",
    x"38CDF02",
    x"38CDBCA",
    x"38CD894",
    x"38CD55E",
    x"38CD229",
    x"38CCEF5",
    x"38CCBC2",
    x"38CC88F",
    x"38CC55D",
    x"38CC22C",
    x"38CBEFC",
    x"38CBBCD",
    x"38CB89E",
    x"38CB571",
    x"38CB244",
    x"38CAF17",
    x"38CABEC",
    x"38CA8C1",
    x"38CA598",
    x"38CA26F",
    x"38C9F46",
    x"38C9C1F",
    x"38C98F8",
    x"38C95D2",
    x"38C92AD",
    x"38C8F89",
    x"38C8C66",
    x"38C8943",
    x"38C8621",
    x"38C8300",
    x"38C7FE0",
    x"38C7CC0",
    x"38C79A1",
    x"38C7683",
    x"38C7366",
    x"38C7049",
    x"38C6D2E",
    x"38C6A13",
    x"38C66F9",
    x"38C63DF",
    x"38C60C7",
    x"38C5DAF",
    x"38C5A98",
    x"38C5782",
    x"38C546C",
    x"38C5157",
    x"38C4E43",
    x"38C4B30",
    x"38C481E",
    x"38C450C",
    x"38C41FB",
    x"38C3EEB",
    x"38C3BDC",
    x"38C38CD",
    x"38C35C0",
    x"38C32B2",
    x"38C2FA6",
    x"38C2C9B",
    x"38C2990",
    x"38C2686",
    x"38C237D",
    x"38C2074",
    x"38C1D6C",
    x"38C1A65",
    x"38C175F",
    x"38C145A",
    x"38C1155",
    x"38C0E51",
    x"38C0B4E",
    x"38C084B",
    x"38C054A",
    x"38C0249",
    x"38BFF49",
    x"38BFC49",
    x"38BF94A",
    x"38BF64C",
    x"38BF34F",
    x"38BF053",
    x"38BED57",
    x"38BEA5C",
    x"38BE762",
    x"38BE468",
    x"38BE170",
    x"38BDE78",
    x"38BDB80",
    x"38BD88A",
    x"38BD594",
    x"38BD29F",
    x"38BCFAB",
    x"38BCCB7",
    x"38BC9C5",
    x"38BC6D2",
    x"38BC3E1",
    x"38BC0F1",
    x"38BBE01",
    x"38BBB12",
    x"38BB823",
    x"38BB535",
    x"38BB249",
    x"38BAF5C",
    x"38BAC71",
    x"38BA986",
    x"38BA69C",
    x"38BA3B3",
    x"38BA0CA",
    x"38B9DE2",
    x"38B9AFB",
    x"38B9815",
    x"38B952F",
    x"38B924A",
    x"38B8F66",
    x"38B8C83",
    x"38B89A0",
    x"38B86BE",
    x"38B83DC",
    x"38B80FC",
    x"38B7E1C",
    x"38B7B3D",
    x"38B785E",
    x"38B7581",
    x"38B72A4",
    x"38B6FC7",
    x"38B6CEC",
    x"38B6A11",
    x"38B6737",
    x"38B645D",
    x"38B6184",
    x"38B5EAC",
    x"38B5BD5",
    x"38B58FF",
    x"38B5629",
    x"38B5353",
    x"38B507F",
    x"38B4DAB",
    x"38B4AD8",
    x"38B4806",
    x"38B4534",
    x"38B4263",
    x"38B3F93",
    x"38B3CC3",
    x"38B39F5",
    x"38B3726",
    x"38B3459",
    x"38B318C",
    x"38B2EC0",
    x"38B2BF5",
    x"38B292A",
    x"38B2660",
    x"38B2397",
    x"38B20CE",
    x"38B1E07",
    x"38B1B3F",
    x"38B1879",
    x"38B15B3",
    x"38B12EE",
    x"38B102A",
    x"38B0D66",
    x"38B0AA3",
    x"38B07E1",
    x"38B051F",
    x"38B025E",
    x"38AFF9E",
    x"38AFCDE",
    x"38AFA1F",
    x"38AF761",
    x"38AF4A4",
    x"38AF1E7",
    x"38AEF2B",
    x"38AEC6F",
    x"38AE9B5",
    x"38AE6FB",
    x"38AE441",
    x"38AE188",
    x"38ADED0",
    x"38ADC19",
    x"38AD962",
    x"38AD6AC",
    x"38AD3F7",
    x"38AD142",
    x"38ACE8E",
    x"38ACBDB",
    x"38AC928",
    x"38AC676",
    x"38AC3C5",
    x"38AC115",
    x"38ABE65",
    x"38ABBB5",
    x"38AB907",
    x"38AB659",
    x"38AB3AC",
    x"38AB0FF",
    x"38AAE53",
    x"38AABA8",
    x"38AA8FD",
    x"38AA653",
    x"38AA3AA",
    x"38AA102",
    x"38A9E5A",
    x"38A9BB2",
    x"38A990C",
    x"38A9666",
    x"38A93C1",
    x"38A911C",
    x"38A8E78",
    x"38A8BD5",
    x"38A8932",
    x"38A8690",
    x"38A83EF",
    x"38A814E",
    x"38A7EAE",
    x"38A7C0F",
    x"38A7970",
    x"38A76D2",
    x"38A7435",
    x"38A7198",
    x"38A6EFC",
    x"38A6C61",
    x"38A69C6",
    x"38A672C",
    x"38A6492",
    x"38A61F9",
    x"38A5F61",
    x"38A5CCA",
    x"38A5A33",
    x"38A579D",
    x"38A5507",
    x"38A5272",
    x"38A4FDE",
    x"38A4D4A",
    x"38A4AB7",
    x"38A4825",
    x"38A4593",
    x"38A4302",
    x"38A4072",
    x"38A3DE2",
    x"38A3B53",
    x"38A38C4",
    x"38A3636",
    x"38A33A9",
    x"38A311C",
    x"38A2E90",
    x"38A2C05",
    x"38A297A",
    x"38A26F0",
    x"38A2467",
    x"38A21DE",
    x"38A1F56",
    x"38A1CCE",
    x"38A1A48",
    x"38A17C1",
    x"38A153C",
    x"38A12B7",
    x"38A1032",
    x"38A0DAF",
    x"38A0B2C",
    x"38A08A9",
    x"38A0627",
    x"38A03A6",
    x"38A0125",
    x"389FEA5",
    x"389FC26",
    x"389F9A7",
    x"389F729",
    x"389F4AC",
    x"389F22F",
    x"389EFB3",
    x"389ED37",
    x"389EABC",
    x"389E842",
    x"389E5C8",
    x"389E34F",
    x"389E0D6",
    x"389DE5E",
    x"389DBE7",
    x"389D970",
    x"389D6FA",
    x"389D485",
    x"389D210",
    x"389CF9C",
    x"389CD28",
    x"389CAB5",
    x"389C843",
    x"389C5D1",
    x"389C360",
    x"389C0EF",
    x"389BE80",
    x"389BC10",
    x"389B9A1",
    x"389B733",
    x"389B4C6",
    x"389B259",
    x"389AFED",
    x"389AD81",
    x"389AB16",
    x"389A8AB",
    x"389A642",
    x"389A3D8",
    x"389A170",
    x"3899F08",
    x"3899CA0",
    x"3899A39",
    x"38997D3",
    x"389956D",
    x"3899308",
    x"38990A4",
    x"3898E40",
    x"3898BDD",
    x"389897A",
    x"3898718",
    x"38984B7",
    x"3898256",
    x"3897FF5",
    x"3897D96",
    x"3897B37",
    x"38978D8",
    x"389767A",
    x"389741D",
    x"38971C0",
    x"3896F64",
    x"3896D08",
    x"3896AAD",
    x"3896853",
    x"38965F9",
    x"38963A0",
    x"3896147",
    x"3895EEF",
    x"3895C98",
    x"3895A41",
    x"38957EB",
    x"3895595",
    x"3895340",
    x"38950EC",
    x"3894E98",
    x"3894C44",
    x"38949F1",
    x"389479F",
    x"389454E",
    x"38942FD",
    x"38940AC",
    x"3893E5C",
    x"3893C0D",
    x"38939BE",
    x"3893770",
    x"3893523",
    x"38932D6",
    x"3893089",
    x"3892E3D",
    x"3892BF2",
    x"38929A7",
    x"389275D",
    x"3892514",
    x"38922CB",
    x"3892082",
    x"3891E3A",
    x"3891BF3",
    x"38919AC",
    x"3891766",
    x"3891521",
    x"38912DC",
    x"3891097",
    x"3890E53",
    x"3890C10",
    x"38909CD",
    x"389078B",
    x"389054A",
    x"3890309",
    x"38900C8",
    x"388FE88",
    x"388FC49",
    x"388FA0A",
    x"388F7CC",
    x"388F58E",
    x"388F351",
    x"388F114",
    x"388EED8",
    x"388EC9D",
    x"388EA62",
    x"388E828",
    x"388E5EE",
    x"388E3B5",
    x"388E17C",
    x"388DF44",
    x"388DD0D",
    x"388DAD6",
    x"388D89F",
    x"388D669",
    x"388D434",
    x"388D1FF",
    x"388CFCB",
    x"388CD97",
    x"388CB64",
    x"388C932",
    x"388C700",
    x"388C4CE",
    x"388C29D",
    x"388C06D",
    x"388BE3D",
    x"388BC0E",
    x"388B9DF",
    x"388B7B1",
    x"388B583",
    x"388B356",
    x"388B129",
    x"388AEFD",
    x"388ACD2",
    x"388AAA7",
    x"388A87D",
    x"388A653",
    x"388A429",
    x"388A201",
    x"3889FD8",
    x"3889DB1",
    x"3889B8A",
    x"3889963",
    x"388973D",
    x"3889517",
    x"38892F2",
    x"38890CE",
    x"3888EAA",
    x"3888C87",
    x"3888A64",
    x"3888841",
    x"3888620",
    x"38883FE",
    x"38881DE",
    x"3887FBD",
    x"3887D9E",
    x"3887B7F",
    x"3887960",
    x"3887742",
    x"3887524",
    x"3887307",
    x"38870EB",
    x"3886ECF",
    x"3886CB3",
    x"3886A98",
    x"388687E",
    x"3886664",
    x"388644B",
    x"3886232",
    x"388601A",
    x"3885E02",
    x"3885BEB",
    x"38859D4",
    x"38857BE",
    x"38855A8",
    x"3885393",
    x"388517E",
    x"3884F6A",
    x"3884D57",
    x"3884B44",
    x"3884931",
    x"388471F",
    x"388450E",
    x"38842FD",
    x"38840EC",
    x"3883EDC",
    x"3883CCD",
    x"3883ABE",
    x"38838AF",
    x"38836A1",
    x"3883494",
    x"3883287",
    x"388307B",
    x"3882E6F",
    x"3882C63",
    x"3882A59",
    x"388284E",
    x"3882644",
    x"388243B",
    x"3882232",
    x"388202A",
    x"3881E22",
    x"3881C1B",
    x"3881A14",
    x"388180E",
    x"3881608",
    x"3881403",
    x"38811FE",
    x"3880FFA",
    x"3880DF6",
    x"3880BF3",
    x"38809F0",
    x"38807EE",
    x"38805EC",
    x"38803EB",
    x"38801EA",
    x"387FFD5",
    x"387FBD5",
    x"387F7D7",
    x"387F3D9",
    x"387EFDD",
    x"387EBE1",
    x"387E7E7",
    x"387E3ED",
    x"387DFF5",
    x"387DBFD",
    x"387D807",
    x"387D411",
    x"387D01D",
    x"387CC29",
    x"387C837",
    x"387C445",
    x"387C055",
    x"387BC65",
    x"387B876",
    x"387B489",
    x"387B09C",
    x"387ACB0",
    x"387A8C6",
    x"387A4DC",
    x"387A0F3",
    x"3879D0C",
    x"3879925",
    x"387953F",
    x"387915A",
    x"3878D76",
    x"3878993",
    x"38785B1",
    x"38781D1",
    x"3877DF1",
    x"3877A12",
    x"3877634",
    x"3877256",
    x"3876E7A",
    x"3876A9F",
    x"38766C5",
    x"38762EC",
    x"3875F14",
    x"3875B3C",
    x"3875766",
    x"3875391",
    x"3874FBC",
    x"3874BE9",
    x"3874816",
    x"3874445",
    x"3874074",
    x"3873CA4",
    x"38738D6",
    x"3873508",
    x"387313B",
    x"3872D6F",
    x"38729A5",
    x"38725DB",
    x"3872212",
    x"3871E4A",
    x"3871A82",
    x"38716BC",
    x"38712F7",
    x"3870F33",
    x"3870B6F",
    x"38707AD",
    x"38703EC",
    x"387002B",
    x"386FC6C",
    x"386F8AD",
    x"386F4EF",
    x"386F132",
    x"386ED77",
    x"386E9BC",
    x"386E602",
    x"386E249",
    x"386DE91",
    x"386DAD9",
    x"386D723",
    x"386D36E",
    x"386CFB9",
    x"386CC06",
    x"386C853",
    x"386C4A2",
    x"386C0F1",
    x"386BD41",
    x"386B993",
    x"386B5E5",
    x"386B238",
    x"386AE8B",
    x"386AAE0",
    x"386A736",
    x"386A38D",
    x"3869FE4",
    x"3869C3D",
    x"3869896",
    x"38694F0",
    x"386914C",
    x"3868DA8",
    x"3868A05",
    x"3868663",
    x"38682C2",
    x"3867F21",
    x"3867B82",
    x"38677E4",
    x"3867446",
    x"38670AA",
    x"3866D0E",
    x"3866973",
    x"38665D9",
    x"3866240",
    x"3865EA8",
    x"3865B11",
    x"386577A",
    x"38653E5",
    x"3865050",
    x"3864CBD",
    x"386492A",
    x"3864598",
    x"3864207",
    x"3863E77",
    x"3863AE8",
    x"386375A",
    x"38633CC",
    x"3863040",
    x"3862CB4",
    x"386292A",
    x"38625A0",
    x"3862217",
    x"3861E8F",
    x"3861B07",
    x"3861781",
    x"38613FC",
    x"3861077",
    x"3860CF3",
    x"3860971",
    x"38605EF",
    x"386026E",
    x"385FEEE",
    x"385FB6E",
    x"385F7F0",
    x"385F472",
    x"385F0F6",
    x"385ED7A",
    x"385E9FF",
    x"385E685",
    x"385E30C",
    x"385DF93",
    x"385DC1C",
    x"385D8A5",
    x"385D52F",
    x"385D1BB",
    x"385CE47",
    x"385CAD3",
    x"385C761",
    x"385C3F0",
    x"385C07F",
    x"385BD10",
    x"385B9A1",
    x"385B633",
    x"385B2C6",
    x"385AF59",
    x"385ABEE",
    x"385A883",
    x"385A51A",
    x"385A1B1",
    x"3859E49",
    x"3859AE2",
    x"385977B",
    x"3859416",
    x"38590B1",
    x"3858D4E",
    x"38589EB",
    x"3858689",
    x"3858327",
    x"3857FC7",
    x"3857C67",
    x"3857909",
    x"38575AB",
    x"385724E",
    x"3856EF2",
    x"3856B97",
    x"385683C",
    x"38564E2",
    x"385618A",
    x"3855E32",
    x"3855ADA",
    x"3855784",
    x"385542F",
    x"38550DA",
    x"3854D86",
    x"3854A33",
    x"38546E1",
    x"3854390",
    x"385403F",
    x"3853CF0",
    x"38539A1",
    x"3853653",
    x"3853306",
    x"3852FB9",
    x"3852C6E",
    x"3852923",
    x"38525D9",
    x"3852290",
    x"3851F48",
    x"3851C01",
    x"38518BA",
    x"3851574",
    x"385122F",
    x"3850EEB",
    x"3850BA8",
    x"3850865",
    x"3850524",
    x"38501E3",
    x"384FEA3",
    x"384FB63",
    x"384F825",
    x"384F4E7",
    x"384F1AB",
    x"384EE6F",
    x"384EB33",
    x"384E7F9",
    x"384E4BF",
    x"384E187",
    x"384DE4F",
    x"384DB17",
    x"384D7E1",
    x"384D4AC",
    x"384D177",
    x"384CE43",
    x"384CB10",
    x"384C7DD",
    x"384C4AC",
    x"384C17B",
    x"384BE4B",
    x"384BB1C",
    x"384B7ED",
    x"384B4C0",
    x"384B193",
    x"384AE67",
    x"384AB3C",
    x"384A811",
    x"384A4E8",
    x"384A1BF",
    x"3849E97",
    x"3849B70",
    x"3849849",
    x"3849523",
    x"38491FF",
    x"3848EDA",
    x"3848BB7",
    x"3848895",
    x"3848573",
    x"3848252",
    x"3847F32",
    x"3847C12",
    x"38478F4",
    x"38475D6",
    x"38472B9",
    x"3846F9C",
    x"3846C81",
    x"3846966",
    x"384664C",
    x"3846333",
    x"384601B",
    x"3845D03",
    x"38459EC",
    x"38456D6",
    x"38453C1",
    x"38450AC",
    x"3844D98",
    x"3844A85",
    x"3844773",
    x"3844462",
    x"3844151",
    x"3843E41",
    x"3843B32",
    x"3843823",
    x"3843516",
    x"3843209",
    x"3842EFD",
    x"3842BF1",
    x"38428E7",
    x"38425DD",
    x"38422D4",
    x"3841FCB",
    x"3841CC4",
    x"38419BD",
    x"38416B7",
    x"38413B2",
    x"38410AD",
    x"3840DA9",
    x"3840AA6",
    x"38407A4",
    x"38404A3",
    x"38401A2",
    x"383FEA2",
    x"383FBA2",
    x"383F8A4",
    x"383F5A6",
    x"383F2A9",
    x"383EFAD",
    x"383ECB1",
    x"383E9B6",
    x"383E6BC",
    x"383E3C3",
    x"383E0CB",
    x"383DDD3",
    x"383DADC",
    x"383D7E5",
    x"383D4F0",
    x"383D1FB",
    x"383CF07",
    x"383CC13",
    x"383C921",
    x"383C62F",
    x"383C33E",
    x"383C04D",
    x"383BD5D",
    x"383BA6E",
    x"383B780",
    x"383B493",
    x"383B1A6",
    x"383AEBA",
    x"383ABCE",
    x"383A8E4",
    x"383A5FA",
    x"383A311",
    x"383A029",
    x"3839D41",
    x"3839A5A",
    x"3839774",
    x"383948E",
    x"38391A9",
    x"3838EC5",
    x"3838BE2",
    x"38388FF",
    x"383861E",
    x"383833C",
    x"383805C",
    x"3837D7C",
    x"3837A9D",
    x"38377BF",
    x"38374E1",
    x"3837204",
    x"3836F28",
    x"3836C4D",
    x"3836972",
    x"3836698",
    x"38363BF",
    x"38360E6",
    x"3835E0E",
    x"3835B37",
    x"3835861",
    x"383558B",
    x"38352B6",
    x"3834FE2",
    x"3834D0E",
    x"3834A3B",
    x"3834769",
    x"3834497",
    x"38341C7",
    x"3833EF7",
    x"3833C27",
    x"3833958",
    x"383368A",
    x"38333BD",
    x"38330F1",
    x"3832E25",
    x"3832B5A",
    x"383288F",
    x"38325C5",
    x"38322FC",
    x"3832034",
    x"3831D6C",
    x"3831AA5",
    x"38317DF",
    x"3831519",
    x"3831254",
    x"3830F90",
    x"3830CCC",
    x"3830A0A",
    x"3830747",
    x"3830486",
    x"38301C5",
    x"382FF05",
    x"382FC46",
    x"382F987",
    x"382F6C9",
    x"382F40B",
    x"382F14F",
    x"382EE93",
    x"382EBD8",
    x"382E91D",
    x"382E663",
    x"382E3AA",
    x"382E0F1",
    x"382DE39",
    x"382DB82",
    x"382D8CB",
    x"382D616",
    x"382D360",
    x"382D0AC",
    x"382CDF8",
    x"382CB45",
    x"382C892",
    x"382C5E1",
    x"382C330",
    x"382C07F",
    x"382BDCF",
    x"382BB20",
    x"382B872",
    x"382B5C4",
    x"382B317",
    x"382B06A",
    x"382ADBF",
    x"382AB14",
    x"382A869",
    x"382A5BF",
    x"382A316",
    x"382A06E",
    x"3829DC6",
    x"3829B1F",
    x"3829878",
    x"38295D3",
    x"382932E",
    x"3829089",
    x"3828DE5",
    x"3828B42",
    x"38288A0",
    x"38285FE",
    x"382835D",
    x"38280BC",
    x"3827E1C",
    x"3827B7D",
    x"38278DE",
    x"3827641",
    x"38273A3",
    x"3827107",
    x"3826E6B",
    x"3826BD0",
    x"3826935",
    x"382669B",
    x"3826402",
    x"3826169",
    x"3825ED1",
    x"3825C3A",
    x"38259A3",
    x"382570D",
    x"3825477",
    x"38251E3",
    x"3824F4E",
    x"3824CBB",
    x"3824A28",
    x"3824796",
    x"3824504",
    x"3824273",
    x"3823FE3",
    x"3823D53",
    x"3823AC4",
    x"3823836",
    x"38235A8",
    x"382331B",
    x"382308F",
    x"3822E03",
    x"3822B78",
    x"38228ED",
    x"3822663",
    x"38223DA",
    x"3822151",
    x"3821EC9",
    x"3821C42",
    x"38219BB",
    x"3821735",
    x"38214B0",
    x"382122B",
    x"3820FA6",
    x"3820D23",
    x"3820AA0",
    x"382081E",
    x"382059C",
    x"382031B",
    x"382009A",
    x"381FE1A",
    x"381FB9B",
    x"381F91D",
    x"381F69F",
    x"381F421",
    x"381F1A5",
    x"381EF28",
    x"381ECAD",
    x"381EA32",
    x"381E7B8",
    x"381E53E",
    x"381E2C5",
    x"381E04D",
    x"381DDD5",
    x"381DB5E",
    x"381D8E7",
    x"381D672",
    x"381D3FC",
    x"381D188",
    x"381CF13",
    x"381CCA0",
    x"381CA2D",
    x"381C7BB",
    x"381C549",
    x"381C2D8",
    x"381C068",
    x"381BDF8",
    x"381BB89",
    x"381B91A",
    x"381B6AC",
    x"381B43F",
    x"381B1D2",
    x"381AF66",
    x"381ACFA",
    x"381AA90",
    x"381A825",
    x"381A5BB",
    x"381A352",
    x"381A0EA",
    x"3819E82",
    x"3819C1B",
    x"38199B4",
    x"381974E",
    x"38194E8",
    x"3819283",
    x"381901F",
    x"3818DBB",
    x"3818B58",
    x"38188F5",
    x"3818694",
    x"3818432",
    x"38181D1",
    x"3817F71",
    x"3817D12",
    x"3817AB3",
    x"3817854",
    x"38175F7",
    x"3817399",
    x"381713D",
    x"3816EE1",
    x"3816C85",
    x"3816A2B",
    x"38167D0",
    x"3816577",
    x"381631E",
    x"38160C5",
    x"3815E6D",
    x"3815C16",
    x"38159BF",
    x"3815769",
    x"3815513",
    x"38152BE",
    x"381506A",
    x"3814E16",
    x"3814BC3",
    x"3814970",
    x"381471E",
    x"38144CD",
    x"381427C",
    x"381402C",
    x"3813DDC",
    x"3813B8D",
    x"381393E",
    x"38136F0",
    x"38134A3",
    x"3813256",
    x"3813009",
    x"3812DBE",
    x"3812B72",
    x"3812928",
    x"38126DE",
    x"3812494",
    x"381224C",
    x"3812003",
    x"3811DBC",
    x"3811B74",
    x"381192E",
    x"38116E8",
    x"38114A2",
    x"381125E",
    x"3811019",
    x"3810DD6",
    x"3810B92",
    x"3810950",
    x"381070E",
    x"38104CC",
    x"381028B",
    x"381004B",
    x"380FE0B",
    x"380FBCC",
    x"380F98D",
    x"380F74F",
    x"380F512",
    x"380F2D5",
    x"380F098",
    x"380EE5C",
    x"380EC21",
    x"380E9E6",
    x"380E7AC",
    x"380E572",
    x"380E339",
    x"380E101",
    x"380DEC9",
    x"380DC91",
    x"380DA5B",
    x"380D824",
    x"380D5EE",
    x"380D3B9",
    x"380D185",
    x"380CF50",
    x"380CD1D",
    x"380CAEA",
    x"380C8B7",
    x"380C686",
    x"380C454",
    x"380C223",
    x"380BFF3",
    x"380BDC3",
    x"380BB94",
    x"380B966",
    x"380B738",
    x"380B50A",
    x"380B2DD",
    x"380B0B1",
    x"380AE85",
    x"380AC59",
    x"380AA2E",
    x"380A804",
    x"380A5DA",
    x"380A3B1",
    x"380A189",
    x"3809F61",
    x"3809D39",
    x"3809B12",
    x"38098EB",
    x"38096C5",
    x"38094A0",
    x"380927B",
    x"3809057",
    x"3808E33",
    x"3808C10",
    x"38089ED",
    x"38087CB",
    x"38085A9",
    x"3808388",
    x"3808167",
    x"3807F47",
    x"3807D28",
    x"3807B09",
    x"38078EA",
    x"38076CC",
    x"38074AF",
    x"3807292",
    x"3807075",
    x"3806E5A",
    x"3806C3E",
    x"3806A23",
    x"3806809",
    x"38065EF",
    x"38063D6",
    x"38061BE",
    x"3805FA5",
    x"3805D8E",
    x"3805B77",
    x"3805960",
    x"380574A",
    x"3805534",
    x"380531F",
    x"380510B",
    x"3804EF7",
    x"3804CE3",
    x"3804AD0",
    x"38048BE",
    x"38046AC",
    x"380449B",
    x"380428A",
    x"3804079",
    x"3803E69",
    x"3803C5A",
    x"3803A4B",
    x"380383D",
    x"380362F",
    x"3803422",
    x"3803215",
    x"3803009",
    x"3802DFD",
    x"3802BF2",
    x"38029E7",
    x"38027DD",
    x"38025D3",
    x"38023CA",
    x"38021C1",
    x"3801FB9",
    x"3801DB1",
    x"3801BAA",
    x"38019A4",
    x"380179D",
    x"3801598",
    x"3801393",
    x"380118E",
    x"3800F8A",
    x"3800D86",
    x"3800B83",
    x"3800980",
    x"380077E",
    x"380057D",
    x"380037C",
    x"380017B",
    x"37FFEF6",
    x"37FFAF7",
    x"37FF6F9",
    x"37FF2FB",
    x"37FEEFF",
    x"37FEB04",
    x"37FE70A",
    x"37FE310",
    x"37FDF18",
    x"37FDB21",
    x"37FD72A",
    x"37FD335",
    x"37FCF41",
    x"37FCB4E",
    x"37FC75B",
    x"37FC36A",
    x"37FBF79",
    x"37FBB8A",
    x"37FB79C",
    x"37FB3AE",
    x"37FAFC2",
    x"37FABD6",
    x"37FA7EC",
    x"37FA402",
    x"37FA01A",
    x"37F9C32",
    x"37F984C",
    x"37F9466",
    x"37F9082",
    x"37F8C9E",
    x"37F88BB",
    x"37F84DA",
    x"37F80F9",
    x"37F7D19",
    x"37F793A",
    x"37F755D",
    x"37F7180",
    x"37F6DA4",
    x"37F69C9",
    x"37F65EF",
    x"37F6216",
    x"37F5E3E",
    x"37F5A67",
    x"37F5691",
    x"37F52BB",
    x"37F4EE7",
    x"37F4B14",
    x"37F4742",
    x"37F4370",
    x"37F3FA0",
    x"37F3BD1",
    x"37F3802",
    x"37F3435",
    x"37F3068",
    x"37F2C9C",
    x"37F28D2",
    x"37F2508",
    x"37F213F",
    x"37F1D77",
    x"37F19B0",
    x"37F15EA",
    x"37F1225",
    x"37F0E61",
    x"37F0A9E",
    x"37F06DC",
    x"37F031B",
    x"37EFF5B",
    x"37EFB9B",
    x"37EF7DD",
    x"37EF41F",
    x"37EF063",
    x"37EECA7",
    x"37EE8EC",
    x"37EE533",
    x"37EE17A",
    x"37EDDC2",
    x"37EDA0B",
    x"37ED655",
    x"37ED2A0",
    x"37ECEEC",
    x"37ECB38",
    x"37EC786",
    x"37EC3D4",
    x"37EC024",
    x"37EBC74",
    x"37EB8C6",
    x"37EB518",
    x"37EB16B",
    x"37EADBF",
    x"37EAA14",
    x"37EA66A",
    x"37EA2C1",
    x"37E9F19",
    x"37E9B72",
    x"37E97CB",
    x"37E9426",
    x"37E9081",
    x"37E8CDD",
    x"37E893B",
    x"37E8599",
    x"37E81F8",
    x"37E7E58",
    x"37E7AB9",
    x"37E771A",
    x"37E737D",
    x"37E6FE1",
    x"37E6C45",
    x"37E68AB",
    x"37E6511",
    x"37E6178",
    x"37E5DE0",
    x"37E5A49",
    x"37E56B3",
    x"37E531E",
    x"37E4F89",
    x"37E4BF6",
    x"37E4863",
    x"37E44D2",
    x"37E4141",
    x"37E3DB1",
    x"37E3A22",
    x"37E3694",
    x"37E3307",
    x"37E2F7B",
    x"37E2BEF",
    x"37E2865",
    x"37E24DB",
    x"37E2152",
    x"37E1DCA",
    x"37E1A43",
    x"37E16BD",
    x"37E1338",
    x"37E0FB4",
    x"37E0C30",
    x"37E08AD",
    x"37E052C",
    x"37E01AB",
    x"37DFE2B",
    x"37DFAAC",
    x"37DF72E",
    x"37DF3B0",
    x"37DF034",
    x"37DECB8",
    x"37DE93D",
    x"37DE5C3",
    x"37DE24A",
    x"37DDED2",
    x"37DDB5B",
    x"37DD7E5",
    x"37DD46F",
    x"37DD0FA",
    x"37DCD87",
    x"37DCA14",
    x"37DC6A2",
    x"37DC330",
    x"37DBFC0",
    x"37DBC50",
    x"37DB8E2",
    x"37DB574",
    x"37DB207",
    x"37DAE9B",
    x"37DAB30",
    x"37DA7C5",
    x"37DA45C",
    x"37DA0F3",
    x"37D9D8B",
    x"37D9A24",
    x"37D96BE",
    x"37D9359",
    x"37D8FF5",
    x"37D8C91",
    x"37D892E",
    x"37D85CD",
    x"37D826C",
    x"37D7F0B",
    x"37D7BAC",
    x"37D784D",
    x"37D74F0",
    x"37D7193",
    x"37D6E37",
    x"37D6ADC",
    x"37D6782",
    x"37D6428",
    x"37D60D0",
    x"37D5D78",
    x"37D5A21",
    x"37D56CB",
    x"37D5375",
    x"37D5021",
    x"37D4CCD",
    x"37D497B",
    x"37D4629",
    x"37D42D7",
    x"37D3F87",
    x"37D3C38",
    x"37D38E9",
    x"37D359B",
    x"37D324E",
    x"37D2F02",
    x"37D2BB7",
    x"37D286C",
    x"37D2523",
    x"37D21DA",
    x"37D1E92",
    x"37D1B4A",
    x"37D1804",
    x"37D14BE",
    x"37D117A",
    x"37D0E36",
    x"37D0AF2",
    x"37D07B0",
    x"37D046F",
    x"37D012E",
    x"37CFDEE",
    x"37CFAAF",
    x"37CF771",
    x"37CF433",
    x"37CF0F7",
    x"37CEDBB",
    x"37CEA80",
    x"37CE746",
    x"37CE40C",
    x"37CE0D3",
    x"37CDD9C",
    x"37CDA65",
    x"37CD72E",
    x"37CD3F9",
    x"37CD0C5",
    x"37CCD91",
    x"37CCA5E",
    x"37CC72C",
    x"37CC3FA",
    x"37CC0CA",
    x"37CBD9A",
    x"37CBA6B",
    x"37CB73D",
    x"37CB40F",
    x"37CB0E2",
    x"37CADB7",
    x"37CAA8C",
    x"37CA761",
    x"37CA438",
    x"37CA10F",
    x"37C9DE7",
    x"37C9AC0",
    x"37C979A",
    x"37C9475",
    x"37C9150",
    x"37C8E2C",
    x"37C8B09",
    x"37C87E6",
    x"37C84C5",
    x"37C81A4",
    x"37C7E84",
    x"37C7B65",
    x"37C7846",
    x"37C7529",
    x"37C720C",
    x"37C6EF0",
    x"37C6BD4",
    x"37C68BA",
    x"37C65A0",
    x"37C6287",
    x"37C5F6F",
    x"37C5C57",
    x"37C5940",
    x"37C562A",
    x"37C5315",
    x"37C5001",
    x"37C4CED",
    x"37C49DA",
    x"37C46C8",
    x"37C43B7",
    x"37C40A7",
    x"37C3D97",
    x"37C3A88",
    x"37C3779",
    x"37C346C",
    x"37C315F",
    x"37C2E53",
    x"37C2B48",
    x"37C283E",
    x"37C2534",
    x"37C222B",
    x"37C1F23",
    x"37C1C1B",
    x"37C1915",
    x"37C160F",
    x"37C130A",
    x"37C1005",
    x"37C0D02",
    x"37C09FF",
    x"37C06FD",
    x"37C03FB",
    x"37C00FB",
    x"37BFDFB",
    x"37BFAFC",
    x"37BF7FD",
    x"37BF500",
    x"37BF203",
    x"37BEF07",
    x"37BEC0B",
    x"37BE911",
    x"37BE617",
    x"37BE31E",
    x"37BE025",
    x"37BDD2E",
    x"37BDA37",
    x"37BD741",
    x"37BD44B",
    x"37BD156",
    x"37BCE62",
    x"37BCB6F",
    x"37BC87D",
    x"37BC58B",
    x"37BC29A",
    x"37BBFAA",
    x"37BBCBA",
    x"37BB9CB",
    x"37BB6DD",
    x"37BB3F0",
    x"37BB103",
    x"37BAE17",
    x"37BAB2C",
    x"37BA842",
    x"37BA558",
    x"37BA26F",
    x"37B9F87",
    x"37B9C9F",
    x"37B99B9",
    x"37B96D2",
    x"37B93ED",
    x"37B9109",
    x"37B8E25",
    x"37B8B41",
    x"37B885F",
    x"37B857D",
    x"37B829C",
    x"37B7FBC",
    x"37B7CDC",
    x"37B79FE",
    x"37B771F",
    x"37B7442",
    x"37B7165",
    x"37B6E89",
    x"37B6BAE",
    x"37B68D3",
    x"37B65FA",
    x"37B6320",
    x"37B6048",
    x"37B5D70",
    x"37B5A99",
    x"37B57C3",
    x"37B54ED",
    x"37B5219",
    x"37B4F44",
    x"37B4C71",
    x"37B499E",
    x"37B46CC",
    x"37B43FB",
    x"37B412A",
    x"37B3E5A",
    x"37B3B8B",
    x"37B38BC",
    x"37B35EF",
    x"37B3321",
    x"37B3055",
    x"37B2D89",
    x"37B2ABE",
    x"37B27F4",
    x"37B252A",
    x"37B2261",
    x"37B1F99",
    x"37B1CD1",
    x"37B1A0B",
    x"37B1744",
    x"37B147F",
    x"37B11BA",
    x"37B0EF6",
    x"37B0C33",
    x"37B0970",
    x"37B06AE",
    x"37B03ED",
    x"37B012C",
    x"37AFE6C",
    x"37AFBAD",
    x"37AF8EE",
    x"37AF630",
    x"37AF373",
    x"37AF0B7",
    x"37AEDFB",
    x"37AEB40",
    x"37AE885",
    x"37AE5CB",
    x"37AE312",
    x"37AE05A",
    x"37ADDA2",
    x"37ADAEB",
    x"37AD835",
    x"37AD57F",
    x"37AD2CA",
    x"37AD016",
    x"37ACD62",
    x"37ACAAF",
    x"37AC7FD",
    x"37AC54B",
    x"37AC29A",
    x"37ABFEA",
    x"37ABD3A",
    x"37ABA8B",
    x"37AB7DD",
    x"37AB52F",
    x"37AB282",
    x"37AAFD6",
    x"37AAD2A",
    x"37AAA7F",
    x"37AA7D5",
    x"37AA52B",
    x"37AA282",
    x"37A9FDA",
    x"37A9D32",
    x"37A9A8B",
    x"37A97E5",
    x"37A953F",
    x"37A929A",
    x"37A8FF6",
    x"37A8D52",
    x"37A8AAF",
    x"37A880D",
    x"37A856B",
    x"37A82CA",
    x"37A802A",
    x"37A7D8A",
    x"37A7AEB",
    x"37A784D",
    x"37A75AF",
    x"37A7312",
    x"37A7076",
    x"37A6DDA",
    x"37A6B3F",
    x"37A68A4",
    x"37A660A",
    x"37A6371",
    x"37A60D9",
    x"37A5E41",
    x"37A5BAA",
    x"37A5913",
    x"37A567D",
    x"37A53E8",
    x"37A5153",
    x"37A4EBF",
    x"37A4C2C",
    x"37A4999",
    x"37A4707",
    x"37A4475",
    x"37A41E5",
    x"37A3F54",
    x"37A3CC5",
    x"37A3A36",
    x"37A37A8",
    x"37A351A",
    x"37A328D",
    x"37A3001",
    x"37A2D75",
    x"37A2AEA",
    x"37A2860",
    x"37A25D6",
    x"37A234D",
    x"37A20C4",
    x"37A1E3D",
    x"37A1BB5",
    x"37A192F",
    x"37A16A9",
    x"37A1423",
    x"37A119F",
    x"37A0F1B",
    x"37A0C97",
    x"37A0A14",
    x"37A0792",
    x"37A0510",
    x"37A028F",
    x"37A000F",
    x"379FD8F",
    x"379FB10",
    x"379F892",
    x"379F614",
    x"379F397",
    x"379F11A",
    x"379EE9E",
    x"379EC23",
    x"379E9A8",
    x"379E72E",
    x"379E4B5",
    x"379E23C",
    x"379DFC4",
    x"379DD4C",
    x"379DAD5",
    x"379D85E",
    x"379D5E9",
    x"379D374",
    x"379D0FF",
    x"379CE8B",
    x"379CC18",
    x"379C9A5",
    x"379C733",
    x"379C4C1",
    x"379C251",
    x"379BFE0",
    x"379BD71",
    x"379BB02",
    x"379B893",
    x"379B625",
    x"379B3B8",
    x"379B14B",
    x"379AEDF",
    x"379AC74",
    x"379AA09",
    x"379A79F",
    x"379A535",
    x"379A2CC",
    x"379A064",
    x"3799DFC",
    x"3799B95",
    x"379992E",
    x"37996C8",
    x"3799463",
    x"37991FE",
    x"3798F9A",
    x"3798D36",
    x"3798AD3",
    x"3798871",
    x"379860F",
    x"37983AE",
    x"379814D",
    x"3797EED",
    x"3797C8E",
    x"3797A2F",
    x"37977D1",
    x"3797573",
    x"3797316",
    x"37970B9",
    x"3796E5E",
    x"3796C02",
    x"37969A8",
    x"379674D",
    x"37964F4",
    x"379629B",
    x"3796043",
    x"3795DEB",
    x"3795B94",
    x"379593D",
    x"37956E7",
    x"3795492",
    x"379523D",
    x"3794FE9",
    x"3794D95",
    x"3794B42",
    x"37948EF",
    x"379469D",
    x"379444C",
    x"37941FB",
    x"3793FAB",
    x"3793D5B",
    x"3793B0C",
    x"37938BE",
    x"3793670",
    x"3793423",
    x"37931D6",
    x"3792F8A",
    x"3792D3E",
    x"3792AF3",
    x"37928A9",
    x"379265F",
    x"3792415",
    x"37921CD",
    x"3791F84",
    x"3791D3D",
    x"3791AF6",
    x"37918AF",
    x"3791669",
    x"3791424",
    x"37911DF",
    x"3790F9B",
    x"3790D58",
    x"3790B15",
    x"37908D2",
    x"3790690",
    x"379044F",
    x"379020E",
    x"378FFCE",
    x"378FD8E",
    x"378FB4F",
    x"378F910",
    x"378F6D2",
    x"378F495",
    x"378F258",
    x"378F01C",
    x"378EDE0",
    x"378EBA5",
    x"378E96A",
    x"378E730",
    x"378E4F7",
    x"378E2BE",
    x"378E085",
    x"378DE4D",
    x"378DC16",
    x"378D9DF",
    x"378D7A9",
    x"378D574",
    x"378D33E",
    x"378D10A",
    x"378CED6",
    x"378CCA3",
    x"378CA70",
    x"378C83D",
    x"378C60C",
    x"378C3DA",
    x"378C1AA",
    x"378BF79",
    x"378BD4A",
    x"378BB1B",
    x"378B8EC",
    x"378B6BE",
    x"378B491",
    x"378B264",
    x"378B038",
    x"378AE0C",
    x"378ABE1",
    x"378A9B6",
    x"378A78C",
    x"378A562",
    x"378A339",
    x"378A111",
    x"3789EE9",
    x"3789CC1",
    x"3789A9A",
    x"3789874",
    x"378964E",
    x"3789429",
    x"3789204",
    x"3788FE0",
    x"3788DBC",
    x"3788B99",
    x"3788976",
    x"3788754",
    x"3788533",
    x"3788312",
    x"37880F1",
    x"3787ED1",
    x"3787CB2",
    x"3787A93",
    x"3787874",
    x"3787656",
    x"3787439",
    x"378721C",
    x"3787000",
    x"3786DE4",
    x"3786BC9",
    x"37869AE",
    x"3786794",
    x"378657B",
    x"3786362",
    x"3786149",
    x"3785F31",
    x"3785D19",
    x"3785B02",
    x"37858EC",
    x"37856D6",
    x"37854C0",
    x"37852AC",
    x"3785097",
    x"3784E83",
    x"3784C70",
    x"3784A5D",
    x"378484B",
    x"3784639",
    x"3784428",
    x"3784217",
    x"3784007",
    x"3783DF7",
    x"3783BE8",
    x"37839D9",
    x"37837CB",
    x"37835BD",
    x"37833B0",
    x"37831A3",
    x"3782F97",
    x"3782D8B",
    x"3782B80",
    x"3782976",
    x"378276B",
    x"3782562",
    x"3782359",
    x"3782150",
    x"3781F48",
    x"3781D40",
    x"3781B39",
    x"3781933",
    x"378172D",
    x"3781527",
    x"3781322",
    x"378111E",
    x"3780F1A",
    x"3780D16",
    x"3780B13",
    x"3780911",
    x"378070F",
    x"378050D",
    x"378030C",
    x"378010C",
    x"377FE18",
    x"377FA19",
    x"377F61B",
    x"377F21E",
    x"377EE22",
    x"377EA26",
    x"377E62C",
    x"377E233",
    x"377DE3B",
    x"377DA44",
    x"377D64E",
    x"377D259",
    x"377CE65",
    x"377CA72",
    x"377C680",
    x"377C28F",
    x"377BE9F",
    x"377BAAF",
    x"377B6C1",
    x"377B2D4",
    x"377AEE8",
    x"377AAFD",
    x"377A712",
    x"377A329",
    x"3779F41",
    x"3779B59",
    x"3779773",
    x"377938E",
    x"3778FA9",
    x"3778BC6",
    x"37787E3",
    x"3778402",
    x"3778021",
    x"3777C42",
    x"3777863",
    x"3777486",
    x"37770A9",
    x"3776CCD",
    x"37768F3",
    x"3776519",
    x"3776140",
    x"3775D68",
    x"3775991",
    x"37755BB",
    x"37751E6",
    x"3774E12",
    x"3774A3F",
    x"377466D",
    x"377429C",
    x"3773ECC",
    x"3773AFD",
    x"377372E",
    x"3773361",
    x"3772F95",
    x"3772BC9",
    x"37727FF",
    x"3772435",
    x"377206D",
    x"3771CA5",
    x"37718DE",
    x"3771519",
    x"3771154",
    x"3770D90",
    x"37709CD",
    x"377060B",
    x"377024A",
    x"376FE8A",
    x"376FACB",
    x"376F70D",
    x"376F34F",
    x"376EF93",
    x"376EBD8",
    x"376E81D",
    x"376E463",
    x"376E0AB",
    x"376DCF3",
    x"376D93C",
    x"376D587",
    x"376D1D2",
    x"376CE1E",
    x"376CA6B",
    x"376C6B8",
    x"376C307",
    x"376BF57",
    x"376BBA8",
    x"376B7F9",
    x"376B44C",
    x"376B09F",
    x"376ACF3",
    x"376A948",
    x"376A59F",
    x"376A1F6",
    x"3769E4E",
    x"3769AA6",
    x"3769700",
    x"376935B",
    x"3768FB7",
    x"3768C13",
    x"3768871",
    x"37684CF",
    x"376812E",
    x"3767D8E",
    x"37679EF",
    x"3767651",
    x"37672B4",
    x"3766F18",
    x"3766B7D",
    x"37667E2",
    x"3766449",
    x"37660B0",
    x"3765D18",
    x"3765982",
    x"37655EC",
    x"3765257",
    x"3764EC2",
    x"3764B2F",
    x"376479D",
    x"376440B",
    x"376407B",
    x"3763CEB",
    x"376395C",
    x"37635CE",
    x"3763241",
    x"3762EB5",
    x"3762B2A",
    x"37627A0",
    x"3762416",
    x"376208E",
    x"3761D06",
    x"376197F",
    x"37615F9",
    x"3761274",
    x"3760EF0",
    x"3760B6D",
    x"37607EA",
    x"3760469",
    x"37600E8",
    x"375FD68",
    x"375F9E9",
    x"375F66B",
    x"375F2EE",
    x"375EF72",
    x"375EBF6",
    x"375E87C",
    x"375E502",
    x"375E189",
    x"375DE11",
    x"375DA9A",
    x"375D724",
    x"375D3AF",
    x"375D03A",
    x"375CCC7",
    x"375C954",
    x"375C5E2",
    x"375C271",
    x"375BF01",
    x"375BB91",
    x"375B823",
    x"375B4B5",
    x"375B149",
    x"375ADDD",
    x"375AA72",
    x"375A708",
    x"375A39E",
    x"375A036",
    x"3759CCE",
    x"3759967",
    x"3759601",
    x"375929C",
    x"3758F38",
    x"3758BD5",
    x"3758872",
    x"3758510",
    x"37581B0",
    x"3757E50",
    x"3757AF0",
    x"3757792",
    x"3757435",
    x"37570D8",
    x"3756D7C",
    x"3756A21",
    x"37566C7",
    x"375636E",
    x"3756016",
    x"3755CBE",
    x"3755967",
    x"3755611",
    x"37552BC",
    x"3754F68",
    x"3754C14",
    x"37548C2",
    x"3754570",
    x"375421F",
    x"3753ECF",
    x"3753B80",
    x"3753831",
    x"37534E4",
    x"3753197",
    x"3752E4B",
    x"3752B00",
    x"37527B5",
    x"375246C",
    x"3752123",
    x"3751DDB",
    x"3751A94",
    x"375174E",
    x"3751408",
    x"37510C4",
    x"3750D80",
    x"3750A3D",
    x"37506FB",
    x"37503BA",
    x"3750079",
    x"374FD39",
    x"374F9FA",
    x"374F6BC",
    x"374F37F",
    x"374F043",
    x"374ED07",
    x"374E9CC",
    x"374E692",
    x"374E359",
    x"374E020",
    x"374DCE9",
    x"374D9B2",
    x"374D67C",
    x"374D347",
    x"374D012",
    x"374CCDF",
    x"374C9AC",
    x"374C67A",
    x"374C349",
    x"374C018",
    x"374BCE9",
    x"374B9BA",
    x"374B68C",
    x"374B35E",
    x"374B032",
    x"374AD06",
    x"374A9DC",
    x"374A6B1",
    x"374A388",
    x"374A060",
    x"3749D38",
    x"3749A11",
    x"37496EB",
    x"37493C6",
    x"37490A1",
    x"3748D7D",
    x"3748A5A",
    x"3748738",
    x"3748417",
    x"37480F6",
    x"3747DD6",
    x"3747AB7",
    x"3747799",
    x"374747B",
    x"374715F",
    x"3746E43",
    x"3746B27",
    x"374680D",
    x"37464F3",
    x"37461DB",
    x"3745EC3",
    x"3745BAB",
    x"3745895",
    x"374557F",
    x"374526A",
    x"3744F56",
    x"3744C42",
    x"3744930",
    x"374461E",
    x"374430D",
    x"3743FFC",
    x"3743CED",
    x"37439DE",
    x"37436D0",
    x"37433C2",
    x"37430B6",
    x"3742DAA",
    x"3742A9F",
    x"3742795",
    x"374248B",
    x"3742182",
    x"3741E7A",
    x"3741B73",
    x"374186D",
    x"3741567",
    x"3741262",
    x"3740F5E",
    x"3740C5A",
    x"3740958",
    x"3740656",
    x"3740354",
    x"3740054",
    x"373FD54",
    x"373FA55",
    x"373F757",
    x"373F45A",
    x"373F15D",
    x"373EE61",
    x"373EB66",
    x"373E86B",
    x"373E571",
    x"373E278",
    x"373DF80",
    x"373DC89",
    x"373D992",
    x"373D69C",
    x"373D3A7",
    x"373D0B2",
    x"373CDBE",
    x"373CACB",
    x"373C7D9",
    x"373C4E7",
    x"373C1F6",
    x"373BF06",
    x"373BC17",
    x"373B928",
    x"373B63A",
    x"373B34D",
    x"373B061",
    x"373AD75",
    x"373AA8A",
    x"373A7A0",
    x"373A4B6",
    x"373A1CD",
    x"3739EE5",
    x"3739BFE",
    x"3739917",
    x"3739631",
    x"373934C",
    x"3739068",
    x"3738D84",
    x"3738AA1",
    x"37387BF",
    x"37384DD",
    x"37381FC",
    x"3737F1C",
    x"3737C3D",
    x"373795E",
    x"3737680",
    x"37373A3",
    x"37370C6",
    x"3736DEA",
    x"3736B0F",
    x"3736835",
    x"373655B",
    x"3736282",
    x"3735FAA",
    x"3735CD2",
    x"37359FB",
    x"3735725",
    x"3735450",
    x"373517B",
    x"3734EA7",
    x"3734BD4",
    x"3734901",
    x"373462F",
    x"373435E",
    x"373408E",
    x"3733DBE",
    x"3733AEF",
    x"3733820",
    x"3733553",
    x"3733286",
    x"3732FB9",
    x"3732CEE",
    x"3732A23",
    x"3732759",
    x"373248F",
    x"37321C6",
    x"3731EFE",
    x"3731C37",
    x"3731970",
    x"37316AA",
    x"37313E5",
    x"3731120",
    x"3730E5C",
    x"3730B99",
    x"37308D7",
    x"3730615",
    x"3730354",
    x"3730093",
    x"372FDD3",
    x"372FB14",
    x"372F856",
    x"372F598",
    x"372F2DB",
    x"372F01F",
    x"372ED63",
    x"372EAA8",
    x"372E7EE",
    x"372E534",
    x"372E27B",
    x"372DFC3",
    x"372DD0B",
    x"372DA54",
    x"372D79E",
    x"372D4E8",
    x"372D233",
    x"372CF7F",
    x"372CCCC",
    x"372CA19",
    x"372C767",
    x"372C4B5",
    x"372C204",
    x"372BF54",
    x"372BCA5",
    x"372B9F6",
    x"372B748",
    x"372B49A",
    x"372B1ED",
    x"372AF41",
    x"372AC96",
    x"372A9EB",
    x"372A741",
    x"372A497",
    x"372A1EE",
    x"3729F46",
    x"3729C9F",
    x"37299F8",
    x"3729752",
    x"37294AC",
    x"3729207",
    x"3728F63",
    x"3728CC0",
    x"3728A1D",
    x"372877B",
    x"37284D9",
    x"3728238",
    x"3727F98",
    x"3727CF8",
    x"3727A5A",
    x"37277BB",
    x"372751E",
    x"3727281",
    x"3726FE4",
    x"3726D49",
    x"3726AAE",
    x"3726813",
    x"372657A",
    x"37262E1",
    x"3726048",
    x"3725DB1",
    x"3725B19",
    x"3725883",
    x"37255ED",
    x"3725358",
    x"37250C4",
    x"3724E30",
    x"3724B9C",
    x"372490A",
    x"3724678",
    x"37243E7",
    x"3724156",
    x"3723EC6",
    x"3723C37",
    x"37239A8",
    x"372371A",
    x"372348C",
    x"37231FF",
    x"3722F73",
    x"3722CE8",
    x"3722A5D",
    x"37227D3",
    x"3722549",
    x"37222C0",
    x"3722038",
    x"3721DB0",
    x"3721B29",
    x"37218A2",
    x"372161C",
    x"3721397",
    x"3721113",
    x"3720E8F",
    x"3720C0B",
    x"3720989",
    x"3720707",
    x"3720485",
    x"3720204",
    x"371FF84",
    x"371FD05",
    x"371FA86",
    x"371F807",
    x"371F58A",
    x"371F30D",
    x"371F090",
    x"371EE14",
    x"371EB99",
    x"371E91E",
    x"371E6A4",
    x"371E42B",
    x"371E1B2",
    x"371DF3A",
    x"371DCC3",
    x"371DA4C",
    x"371D7D6",
    x"371D560",
    x"371D2EB",
    x"371D076",
    x"371CE03",
    x"371CB8F",
    x"371C91D",
    x"371C6AB",
    x"371C43A",
    x"371C1C9",
    x"371BF59",
    x"371BCE9",
    x"371BA7A",
    x"371B80C",
    x"371B59E",
    x"371B331",
    x"371B0C5",
    x"371AE59",
    x"371ABED",
    x"371A983",
    x"371A719",
    x"371A4AF",
    x"371A246",
    x"3719FDE",
    x"3719D76",
    x"3719B0F",
    x"37198A9",
    x"3719643",
    x"37193DE",
    x"3719179",
    x"3718F15",
    x"3718CB2",
    x"3718A4F",
    x"37187EC",
    x"371858B",
    x"371832A",
    x"37180C9",
    x"3717E69",
    x"3717C0A",
    x"37179AB",
    x"371774D",
    x"37174F0",
    x"3717293",
    x"3717036",
    x"3716DDA",
    x"3716B7F",
    x"3716925",
    x"37166CB",
    x"3716471",
    x"3716219",
    x"3715FC0",
    x"3715D69",
    x"3715B12",
    x"37158BB",
    x"3715665",
    x"3715410",
    x"37151BB",
    x"3714F67",
    x"3714D13",
    x"3714AC0",
    x"371486E",
    x"371461C",
    x"37143CB",
    x"371417A",
    x"3713F2A",
    x"3713CDB",
    x"3713A8C",
    x"371383E",
    x"37135F0",
    x"37133A3",
    x"3713156",
    x"3712F0A",
    x"3712CBE",
    x"3712A74",
    x"3712829",
    x"37125DF",
    x"3712396",
    x"371214E",
    x"3711F06",
    x"3711CBE",
    x"3711A77",
    x"3711831",
    x"37115EB",
    x"37113A6",
    x"3711161",
    x"3710F1D",
    x"3710CDA",
    x"3710A97",
    x"3710854",
    x"3710613",
    x"37103D1",
    x"3710191",
    x"370FF51",
    x"370FD11",
    x"370FAD2",
    x"370F894",
    x"370F656",
    x"370F418",
    x"370F1DC",
    x"370EFA0",
    x"370ED64",
    x"370EB29",
    x"370E8EE",
    x"370E6B4",
    x"370E47B",
    x"370E242",
    x"370E00A",
    x"370DDD2",
    x"370DB9B",
    x"370D964",
    x"370D72E",
    x"370D4F9",
    x"370D2C4",
    x"370D08F",
    x"370CE5B",
    x"370CC28",
    x"370C9F5",
    x"370C7C3",
    x"370C592",
    x"370C360",
    x"370C130",
    x"370BF00",
    x"370BCD0",
    x"370BAA1",
    x"370B873",
    x"370B645",
    x"370B418",
    x"370B1EB",
    x"370AFBF",
    x"370AD93",
    x"370AB68",
    x"370A93E",
    x"370A714",
    x"370A4EA",
    x"370A2C1",
    x"370A099",
    x"3709E71",
    x"3709C49",
    x"3709A23",
    x"37097FC",
    x"37095D7",
    x"37093B1",
    x"370918D",
    x"3708F69",
    x"3708D45",
    x"3708B22",
    x"3708900",
    x"37086DE",
    x"37084BC",
    x"370829B",
    x"370807B",
    x"3707E5B",
    x"3707C3C",
    x"3707A1D",
    x"37077FF",
    x"37075E1",
    x"37073C4",
    x"37071A7",
    x"3706F8B",
    x"3706D6F",
    x"3706B54",
    x"3706939",
    x"370671F",
    x"3706506",
    x"37062ED",
    x"37060D4",
    x"3705EBD",
    x"3705CA5",
    x"3705A8E",
    x"3705878",
    x"3705662",
    x"370544D",
    x"3705238",
    x"3705023",
    x"3704E10",
    x"3704BFC",
    x"37049EA",
    x"37047D8",
    x"37045C6",
    x"37043B5",
    x"37041A4",
    x"3703F94",
    x"3703D84",
    x"3703B75",
    x"3703966",
    x"3703758",
    x"370354B",
    x"370333E",
    x"3703131",
    x"3702F25",
    x"3702D1A",
    x"3702B0F",
    x"3702904",
    x"37026FA",
    x"37024F1",
    x"37022E8",
    x"37020DF",
    x"3701ED7",
    x"3701CD0",
    x"3701AC9",
    x"37018C2",
    x"37016BC",
    x"37014B7",
    x"37012B2",
    x"37010AE",
    x"3700EAA",
    x"3700CA6",
    x"3700AA3",
    x"37008A1",
    x"370069F",
    x"370049E",
    x"370029D",
    x"370009C",
    x"36FFD39",
    x"36FF93A",
    x"36FF53D",
    x"36FF140",
    x"36FED44",
    x"36FE949",
    x"36FE54F",
    x"36FE157",
    x"36FDD5F",
    x"36FD968",
    x"36FD572",
    x"36FD17D",
    x"36FCD89",
    x"36FC996",
    x"36FC5A4",
    x"36FC1B4",
    x"36FBDC4",
    x"36FB9D5",
    x"36FB5E7",
    x"36FB1FA",
    x"36FAE0E",
    x"36FAA23",
    x"36FA639",
    x"36FA250",
    x"36F9E67",
    x"36F9A80",
    x"36F969A",
    x"36F92B5",
    x"36F8ED1",
    x"36F8AEE",
    x"36F870B",
    x"36F832A",
    x"36F7F4A",
    x"36F7B6A",
    x"36F778C",
    x"36F73AF",
    x"36F6FD2",
    x"36F6BF7",
    x"36F681C",
    x"36F6443",
    x"36F606A",
    x"36F5C93",
    x"36F58BC",
    x"36F54E6",
    x"36F5111",
    x"36F4D3E",
    x"36F496B",
    x"36F4599",
    x"36F41C8",
    x"36F3DF8",
    x"36F3A29",
    x"36F365B",
    x"36F328E",
    x"36F2EC2",
    x"36F2AF6",
    x"36F272C",
    x"36F2363",
    x"36F1F9A",
    x"36F1BD3",
    x"36F180D",
    x"36F1447",
    x"36F1082",
    x"36F0CBF",
    x"36F08FC",
    x"36F053A",
    x"36F0179",
    x"36EFDBA",
    x"36EF9FB",
    x"36EF63D",
    x"36EF27F",
    x"36EEEC3",
    x"36EEB08",
    x"36EE74E",
    x"36EE394",
    x"36EDFDC",
    x"36EDC24",
    x"36ED86E",
    x"36ED4B8",
    x"36ED104",
    x"36ECD50",
    x"36EC99D",
    x"36EC5EB",
    x"36EC23A",
    x"36EBE8A",
    x"36EBADB",
    x"36EB72C",
    x"36EB37F",
    x"36EAFD3",
    x"36EAC27",
    x"36EA87D",
    x"36EA4D3",
    x"36EA12A",
    x"36E9D82",
    x"36E99DB",
    x"36E9635",
    x"36E9290",
    x"36E8EEC",
    x"36E8B49",
    x"36E87A6",
    x"36E8405",
    x"36E8064",
    x"36E7CC5",
    x"36E7926",
    x"36E7588",
    x"36E71EB",
    x"36E6E4F",
    x"36E6AB4",
    x"36E671A",
    x"36E6381",
    x"36E5FE8",
    x"36E5C51",
    x"36E58BA",
    x"36E5524",
    x"36E518F",
    x"36E4DFB",
    x"36E4A68",
    x"36E46D6",
    x"36E4345",
    x"36E3FB5",
    x"36E3C25",
    x"36E3897",
    x"36E3509",
    x"36E317C",
    x"36E2DF0",
    x"36E2A65",
    x"36E26DB",
    x"36E2352",
    x"36E1FC9",
    x"36E1C42",
    x"36E18BB",
    x"36E1535",
    x"36E11B1",
    x"36E0E2D",
    x"36E0AA9",
    x"36E0727",
    x"36E03A6",
    x"36E0025",
    x"36DFCA6",
    x"36DF927",
    x"36DF5A9",
    x"36DF22C",
    x"36DEEB0",
    x"36DEB35",
    x"36DE7BB",
    x"36DE441",
    x"36DE0C8",
    x"36DDD51",
    x"36DD9DA",
    x"36DD664",
    x"36DD2EF",
    x"36DCF7A",
    x"36DCC07",
    x"36DC894",
    x"36DC523",
    x"36DC1B2",
    x"36DBE42",
    x"36DBAD3",
    x"36DB764",
    x"36DB3F7",
    x"36DB08A",
    x"36DAD1F",
    x"36DA9B4",
    x"36DA64A",
    x"36DA2E1",
    x"36D9F78",
    x"36D9C11",
    x"36D98AA",
    x"36D9544",
    x"36D91E0",
    x"36D8E7C",
    x"36D8B18",
    x"36D87B6",
    x"36D8455",
    x"36D80F4",
    x"36D7D94",
    x"36D7A35",
    x"36D76D7",
    x"36D737A",
    x"36D701D",
    x"36D6CC2",
    x"36D6967",
    x"36D660D",
    x"36D62B4",
    x"36D5F5C",
    x"36D5C04",
    x"36D58AE",
    x"36D5558",
    x"36D5203",
    x"36D4EAF",
    x"36D4B5B",
    x"36D4809",
    x"36D44B7",
    x"36D4167",
    x"36D3E17",
    x"36D3AC8",
    x"36D3779",
    x"36D342C",
    x"36D30DF",
    x"36D2D93",
    x"36D2A49",
    x"36D26FE",
    x"36D23B5",
    x"36D206C",
    x"36D1D25",
    x"36D19DE",
    x"36D1698",
    x"36D1353",
    x"36D100E",
    x"36D0CCB",
    x"36D0988",
    x"36D0646",
    x"36D0305",
    x"36CFFC4",
    x"36CFC85",
    x"36CF946",
    x"36CF608",
    x"36CF2CB",
    x"36CEF8F",
    x"36CEC53",
    x"36CE919",
    x"36CE5DF",
    x"36CE2A6",
    x"36CDF6D",
    x"36CDC36",
    x"36CD8FF",
    x"36CD5C9",
    x"36CD294",
    x"36CCF60",
    x"36CCC2D",
    x"36CC8FA",
    x"36CC5C8",
    x"36CC297",
    x"36CBF67",
    x"36CBC37",
    x"36CB909",
    x"36CB5DB",
    x"36CB2AE",
    x"36CAF82",
    x"36CAC56",
    x"36CA92B",
    x"36CA602",
    x"36CA2D8",
    x"36C9FB0",
    x"36C9C89",
    x"36C9962",
    x"36C963C",
    x"36C9317",
    x"36C8FF2",
    x"36C8CCF",
    x"36C89AC",
    x"36C868A",
    x"36C8369",
    x"36C8048",
    x"36C7D29",
    x"36C7A0A",
    x"36C76EC",
    x"36C73CE",
    x"36C70B2",
    x"36C6D96",
    x"36C6A7B",
    x"36C6761",
    x"36C6447",
    x"36C612E",
    x"36C5E17",
    x"36C5AFF",
    x"36C57E9",
    x"36C54D3",
    x"36C51BF",
    x"36C4EAB",
    x"36C4B97",
    x"36C4885",
    x"36C4573",
    x"36C4262",
    x"36C3F52",
    x"36C3C42",
    x"36C3934",
    x"36C3626",
    x"36C3319",
    x"36C300C",
    x"36C2D01",
    x"36C29F6",
    x"36C26EC",
    x"36C23E2",
    x"36C20DA",
    x"36C1DD2",
    x"36C1ACB",
    x"36C17C4",
    x"36C14BF",
    x"36C11BA",
    x"36C0EB6",
    x"36C0BB3",
    x"36C08B0",
    x"36C05AE",
    x"36C02AD",
    x"36BFFAD",
    x"36BFCAD",
    x"36BF9AF",
    x"36BF6B1",
    x"36BF3B3",
    x"36BF0B7",
    x"36BEDBB",
    x"36BEAC0",
    x"36BE7C6",
    x"36BE4CC",
    x"36BE1D3",
    x"36BDEDB",
    x"36BDBE4",
    x"36BD8ED",
    x"36BD5F7",
    x"36BD302",
    x"36BD00E",
    x"36BCD1A",
    x"36BCA27",
    x"36BC735",
    x"36BC444",
    x"36BC153",
    x"36BBE63",
    x"36BBB74",
    x"36BB885",
    x"36BB597",
    x"36BB2AA",
    x"36BAFBE",
    x"36BACD3",
    x"36BA9E8",
    x"36BA6FE",
    x"36BA414",
    x"36BA12C",
    x"36B9E44",
    x"36B9B5C",
    x"36B9876",
    x"36B9590",
    x"36B92AB",
    x"36B8FC7",
    x"36B8CE3",
    x"36B8A00",
    x"36B871E",
    x"36B843D",
    x"36B815C",
    x"36B7E7C",
    x"36B7B9D",
    x"36B78BE",
    x"36B75E1",
    x"36B7303",
    x"36B7027",
    x"36B6D4B",
    x"36B6A70",
    x"36B6796",
    x"36B64BD",
    x"36B61E4",
    x"36B5F0C",
    x"36B5C34",
    x"36B595E",
    x"36B5688",
    x"36B53B2",
    x"36B50DE",
    x"36B4E0A",
    x"36B4B37",
    x"36B4864",
    x"36B4593",
    x"36B42C1",
    x"36B3FF1",
    x"36B3D22",
    x"36B3A53",
    x"36B3784",
    x"36B34B7",
    x"36B31EA",
    x"36B2F1E",
    x"36B2C52",
    x"36B2988",
    x"36B26BE",
    x"36B23F4",
    x"36B212C",
    x"36B1E64",
    x"36B1B9C",
    x"36B18D6",
    x"36B1610",
    x"36B134B",
    x"36B1086",
    x"36B0DC3",
    x"36B0B00",
    x"36B083D",
    x"36B057B",
    x"36B02BA",
    x"36AFFFA",
    x"36AFD3A",
    x"36AFA7B",
    x"36AF7BD",
    x"36AF500",
    x"36AF243",
    x"36AEF86",
    x"36AECCB",
    x"36AEA10",
    x"36AE756",
    x"36AE49C",
    x"36AE1E4",
    x"36ADF2B",
    x"36ADC74",
    x"36AD9BD",
    x"36AD707",
    x"36AD452",
    x"36AD19D",
    x"36ACEE9",
    x"36ACC35",
    x"36AC983",
    x"36AC6D1",
    x"36AC41F",
    x"36AC16F",
    x"36ABEBF",
    x"36ABC0F",
    x"36AB961",
    x"36AB6B3",
    x"36AB405",
    x"36AB159",
    x"36AAEAD",
    x"36AAC01",
    x"36AA957",
    x"36AA6AD",
    x"36AA403",
    x"36AA15B",
    x"36A9EB3",
    x"36A9C0B",
    x"36A9965",
    x"36A96BF",
    x"36A9419",
    x"36A9174",
    x"36A8ED0",
    x"36A8C2D",
    x"36A898A",
    x"36A86E8",
    x"36A8447",
    x"36A81A6",
    x"36A7F06",
    x"36A7C67",
    x"36A79C8",
    x"36A772A",
    x"36A748C",
    x"36A71EF",
    x"36A6F53",
    x"36A6CB8",
    x"36A6A1D",
    x"36A6783",
    x"36A64E9",
    x"36A6250",
    x"36A5FB8",
    x"36A5D20",
    x"36A5A89",
    x"36A57F3",
    x"36A555D",
    x"36A52C8",
    x"36A5034",
    x"36A4DA0",
    x"36A4B0D",
    x"36A487B",
    x"36A45E9",
    x"36A4358",
    x"36A40C7",
    x"36A3E38",
    x"36A3BA8",
    x"36A391A",
    x"36A368C",
    x"36A33FE",
    x"36A3172",
    x"36A2EE6",
    x"36A2C5A",
    x"36A29CF",
    x"36A2745",
    x"36A24BC",
    x"36A2233",
    x"36A1FAB",
    x"36A1D23",
    x"36A1A9C",
    x"36A1816",
    x"36A1590",
    x"36A130B",
    x"36A1087",
    x"36A0E03",
    x"36A0B80",
    x"36A08FD",
    x"36A067B",
    x"36A03FA",
    x"36A0179",
    x"369FEF9",
    x"369FC7A",
    x"369F9FB",
    x"369F77D",
    x"369F4FF",
    x"369F282",
    x"369F006",
    x"369ED8A",
    x"369EB0F",
    x"369E895",
    x"369E61B",
    x"369E3A2",
    x"369E129",
    x"369DEB1",
    x"369DC3A",
    x"369D9C3",
    x"369D74D",
    x"369D4D7",
    x"369D262",
    x"369CFEE",
    x"369CD7A",
    x"369CB07",
    x"369C895",
    x"369C623",
    x"369C3B2",
    x"369C141",
    x"369BED1",
    x"369BC62",
    x"369B9F3",
    x"369B785",
    x"369B517",
    x"369B2AA",
    x"369B03E",
    x"369ADD2",
    x"369AB67",
    x"369A8FC",
    x"369A692",
    x"369A429",
    x"369A1C0",
    x"3699F58",
    x"3699CF1",
    x"3699A8A",
    x"3699823",
    x"36995BE",
    x"3699359",
    x"36990F4",
    x"3698E90",
    x"3698C2D",
    x"36989CA",
    x"3698768",
    x"3698506",
    x"36982A5",
    x"3698045",
    x"3697DE5",
    x"3697B86",
    x"3697927",
    x"36976C9",
    x"369746C",
    x"369720F",
    x"3696FB3",
    x"3696D57",
    x"3696AFC",
    x"36968A2",
    x"3696648",
    x"36963EF",
    x"3696196",
    x"3695F3E",
    x"3695CE6",
    x"3695A8F",
    x"3695839",
    x"36955E3",
    x"369538E",
    x"369513A",
    x"3694EE6",
    x"3694C92",
    x"3694A3F",
    x"36947ED",
    x"369459B",
    x"369434A",
    x"36940FA",
    x"3693EAA",
    x"3693C5A",
    x"3693A0C",
    x"36937BD",
    x"3693570",
    x"3693323",
    x"36930D6",
    x"3692E8A",
    x"3692C3F",
    x"36929F4",
    x"36927AA",
    x"3692560",
    x"3692317",
    x"36920CF",
    x"3691E87",
    x"3691C3F",
    x"36919F9",
    x"36917B2",
    x"369156D",
    x"3691328",
    x"36910E3",
    x"3690E9F",
    x"3690C5C",
    x"3690A19",
    x"36907D7",
    x"3690595",
    x"3690354",
    x"3690114",
    x"368FED4",
    x"368FC94",
    x"368FA55",
    x"368F817",
    x"368F5D9",
    x"368F39C",
    x"368F15F",
    x"368EF23",
    x"368ECE8",
    x"368EAAD",
    x"368E872",
    x"368E639",
    x"368E3FF",
    x"368E1C7",
    x"368DF8E",
    x"368DD57",
    x"368DB20",
    x"368D8E9",
    x"368D6B3",
    x"368D47E",
    x"368D249",
    x"368D015",
    x"368CDE1",
    x"368CBAE",
    x"368C97B",
    x"368C749",
    x"368C518",
    x"368C2E7",
    x"368C0B6",
    x"368BE86",
    x"368BC57",
    x"368BA28",
    x"368B7FA",
    x"368B5CC",
    x"368B39F",
    x"368B172",
    x"368AF46",
    x"368AD1B",
    x"368AAF0",
    x"368A8C5",
    x"368A69B",
    x"368A472",
    x"368A249",
    x"368A021",
    x"3689DF9",
    x"3689BD2",
    x"36899AB",
    x"3689785",
    x"368955F",
    x"368933A",
    x"3689116",
    x"3688EF2",
    x"3688CCE",
    x"3688AAB",
    x"3688889",
    x"3688667",
    x"3688446",
    x"3688225",
    x"3688005",
    x"3687DE5",
    x"3687BC6",
    x"36879A7",
    x"3687789",
    x"368756B",
    x"368734E",
    x"3687131",
    x"3686F15",
    x"3686CFA",
    x"3686ADF",
    x"36868C5",
    x"36866AB",
    x"3686491",
    x"3686278",
    x"3686060",
    x"3685E48",
    x"3685C31",
    x"3685A1A",
    x"3685804",
    x"36855EE",
    x"36853D9",
    x"36851C4",
    x"3684FB0",
    x"3684D9C",
    x"3684B89",
    x"3684976",
    x"3684764",
    x"3684553",
    x"3684342",
    x"3684131",
    x"3683F21",
    x"3683D12",
    x"3683B03",
    x"36838F4",
    x"36836E6",
    x"36834D9",
    x"36832CC",
    x"36830BF",
    x"3682EB3",
    x"3682CA8",
    x"3682A9D",
    x"3682893",
    x"3682689",
    x"368247F",
    x"3682276",
    x"368206E",
    x"3681E66",
    x"3681C5F",
    x"3681A58",
    x"3681852",
    x"368164C",
    x"3681447",
    x"3681242",
    x"368103D",
    x"3680E3A",
    x"3680C36",
    x"3680A33",
    x"3680831",
    x"368062F",
    x"368042E",
    x"368022D",
    x"368002D",
    x"367FC5B",
    x"367F85C",
    x"367F45F",
    x"367F062",
    x"367EC67",
    x"367E86C",
    x"367E472",
    x"367E07A",
    x"367DC82",
    x"367D88B",
    x"367D496",
    x"367D0A1",
    x"367CCAD",
    x"367C8BB",
    x"367C4C9",
    x"367C0D8",
    x"367BCE9",
    x"367B8FA",
    x"367B50C",
    x"367B11F",
    x"367AD34",
    x"367A949",
    x"367A55F",
    x"367A176",
    x"3679D8E",
    x"36799A7",
    x"36795C1",
    x"36791DC",
    x"3678DF9",
    x"3678A16",
    x"3678633",
    x"3678252",
    x"3677E72",
    x"3677A93",
    x"36776B5",
    x"36772D8",
    x"3676EFC",
    x"3676B20",
    x"3676746",
    x"367636D",
    x"3675F94",
    x"3675BBD",
    x"36757E6",
    x"3675411",
    x"367503C",
    x"3674C69",
    x"3674896",
    x"36744C5",
    x"36740F4",
    x"3673D24",
    x"3673955",
    x"3673587",
    x"36731BA",
    x"3672DEF",
    x"3672A24",
    x"3672659",
    x"3672290",
    x"3671EC8",
    x"3671B01",
    x"367173B",
    x"3671375",
    x"3670FB1",
    x"3670BED",
    x"367082B",
    x"3670469",
    x"36700A9",
    x"366FCE9",
    x"366F92A",
    x"366F56C",
    x"366F1B0",
    x"366EDF4",
    x"366EA39",
    x"366E67F",
    x"366E2C5",
    x"366DF0D",
    x"366DB56",
    x"366D79F",
    x"366D3EA",
    x"366D036",
    x"366CC82",
    x"366C8CF",
    x"366C51E",
    x"366C16D",
    x"366BDBD",
    x"366BA0E",
    x"366B660",
    x"366B2B3",
    x"366AF06",
    x"366AB5B",
    x"366A7B1",
    x"366A407",
    x"366A05F",
    x"3669CB7",
    x"3669910",
    x"366956B",
    x"36691C6",
    x"3668E22",
    x"3668A7F",
    x"36686DC",
    x"366833B",
    x"3667F9B",
    x"3667BFB",
    x"366785D",
    x"36674BF",
    x"3667122",
    x"3666D87",
    x"36669EC",
    x"3666652",
    x"36662B9",
    x"3665F20",
    x"3665B89",
    x"36657F3",
    x"366545D",
    x"36650C8",
    x"3664D35",
    x"36649A2",
    x"3664610",
    x"366427F",
    x"3663EEF",
    x"3663B5F",
    x"36637D1",
    x"3663443",
    x"36630B7",
    x"3662D2B",
    x"36629A0",
    x"3662616",
    x"366228D",
    x"3661F05",
    x"3661B7E",
    x"36617F7",
    x"3661472",
    x"36610ED",
    x"3660D69",
    x"36609E6",
    x"3660664",
    x"36602E3",
    x"365FF63",
    x"365FBE3",
    x"365F865",
    x"365F4E7",
    x"365F16A",
    x"365EDEE",
    x"365EA73",
    x"365E6F9",
    x"365E380",
    x"365E007",
    x"365DC90",
    x"365D919",
    x"365D5A3",
    x"365D22E",
    x"365CEBA",
    x"365CB47",
    x"365C7D5",
    x"365C463",
    x"365C0F2",
    x"365BD83",
    x"365BA14",
    x"365B6A6",
    x"365B338",
    x"365AFCC",
    x"365AC60",
    x"365A8F6",
    x"365A58C",
    x"365A223",
    x"3659EBB",
    x"3659B54",
    x"36597ED",
    x"3659488",
    x"3659123",
    x"3658DBF",
    x"3658A5C",
    x"36586FA",
    x"3658399",
    x"3658038",
    x"3657CD8",
    x"365797A",
    x"365761C",
    x"36572BF",
    x"3656F62",
    x"3656C07",
    x"36568AC",
    x"3656553",
    x"36561FA",
    x"3655EA2",
    x"3655B4A",
    x"36557F4",
    x"365549E",
    x"365514A",
    x"3654DF6",
    x"3654AA3",
    x"3654750",
    x"36543FF",
    x"36540AE",
    x"3653D5F",
    x"3653A10",
    x"36536C2",
    x"3653374",
    x"3653028",
    x"3652CDC",
    x"3652991",
    x"3652647",
    x"36522FE",
    x"3651FB6",
    x"3651C6E",
    x"3651928",
    x"36515E2",
    x"365129D",
    x"3650F59",
    x"3650C15",
    x"36508D3",
    x"3650591",
    x"3650250",
    x"364FF10",
    x"364FBD0",
    x"364F892",
    x"364F554",
    x"364F217",
    x"364EEDB",
    x"364EBA0",
    x"364E865",
    x"364E52B",
    x"364E1F2",
    x"364DEBA",
    x"364DB83",
    x"364D84D",
    x"364D517",
    x"364D1E2",
    x"364CEAE",
    x"364CB7B",
    x"364C848",
    x"364C517",
    x"364C1E6",
    x"364BEB6",
    x"364BB86",
    x"364B858",
    x"364B52A",
    x"364B1FD",
    x"364AED1",
    x"364ABA6",
    x"364A87B",
    x"364A552",
    x"364A229",
    x"3649F01",
    x"3649BD9",
    x"36498B3",
    x"364958D",
    x"3649268",
    x"3648F44",
    x"3648C20",
    x"36488FE",
    x"36485DC",
    x"36482BB",
    x"3647F9A",
    x"3647C7B",
    x"364795C",
    x"364763E",
    x"3647321",
    x"3647005",
    x"3646CE9",
    x"36469CE",
    x"36466B4",
    x"364639B",
    x"3646082",
    x"3645D6B",
    x"3645A54",
    x"364573D",
    x"3645428",
    x"3645113",
    x"3644DFF",
    x"3644AEC",
    x"36447DA",
    x"36444C8",
    x"36441B8",
    x"3643EA8",
    x"3643B98",
    x"364388A",
    x"364357C",
    x"364326F",
    x"3642F63",
    x"3642C57",
    x"364294D",
    x"3642643",
    x"3642339",
    x"3642031",
    x"3641D29",
    x"3641A22",
    x"364171C",
    x"3641417",
    x"3641112",
    x"3640E0E",
    x"3640B0B",
    x"3640809",
    x"3640507",
    x"3640206",
    x"363FF06",
    x"363FC07",
    x"363F908",
    x"363F60A",
    x"363F30D",
    x"363F011",
    x"363ED15",
    x"363EA1A",
    x"363E720",
    x"363E427",
    x"363E12E",
    x"363DE36",
    x"363DB3F",
    x"363D848",
    x"363D553",
    x"363D25E",
    x"363CF6A",
    x"363CC76",
    x"363C983",
    x"363C691",
    x"363C3A0",
    x"363C0AF",
    x"363BDC0",
    x"363BAD1",
    x"363B7E2",
    x"363B4F5",
    x"363B208",
    x"363AF1C",
    x"363AC30",
    x"363A946",
    x"363A65C",
    x"363A372",
    x"363A08A",
    x"3639DA2",
    x"3639ABB",
    x"36397D5",
    x"36394EF",
    x"363920A",
    x"3638F26",
    x"3638C43",
    x"3638960",
    x"363867E",
    x"363839D",
    x"36380BC",
    x"3637DDC",
    x"3637AFD",
    x"363781F",
    x"3637541",
    x"3637264",
    x"3636F88",
    x"3636CAC",
    x"36369D2",
    x"36366F8",
    x"363641E",
    x"3636146",
    x"3635E6E",
    x"3635B96",
    x"36358C0",
    x"36355EA",
    x"3635315",
    x"3635040",
    x"3634D6D",
    x"3634A9A",
    x"36347C7",
    x"36344F6",
    x"3634225",
    x"3633F55",
    x"3633C85",
    x"36339B6",
    x"36336E8",
    x"363341B",
    x"363314E",
    x"3632E82",
    x"3632BB7",
    x"36328EC",
    x"3632623",
    x"3632359",
    x"3632091",
    x"3631DC9",
    x"3631B02",
    x"363183C",
    x"3631576",
    x"36312B1",
    x"3630FED",
    x"3630D29",
    x"3630A66",
    x"36307A4",
    x"36304E2",
    x"3630221",
    x"362FF61",
    x"362FCA2",
    x"362F9E3",
    x"362F725",
    x"362F467",
    x"362F1AA",
    x"362EEEE",
    x"362EC33",
    x"362E978",
    x"362E6BE",
    x"362E405",
    x"362E14C",
    x"362DE94",
    x"362DBDD",
    x"362D926",
    x"362D670",
    x"362D3BB",
    x"362D107",
    x"362CE53",
    x"362CB9F",
    x"362C8ED",
    x"362C63B",
    x"362C38A",
    x"362C0D9",
    x"362BE29",
    x"362BB7A",
    x"362B8CB",
    x"362B61E",
    x"362B370",
    x"362B0C4",
    x"362AE18",
    x"362AB6D",
    x"362A8C2",
    x"362A618",
    x"362A36F",
    x"362A0C7",
    x"3629E1F",
    x"3629B78",
    x"36298D1",
    x"362962B",
    x"3629386",
    x"36290E2",
    x"3628E3E",
    x"3628B9A",
    x"36288F8",
    x"3628656",
    x"36283B5",
    x"3628114",
    x"3627E74",
    x"3627BD5",
    x"3627936",
    x"3627698",
    x"36273FB",
    x"362715E",
    x"3626EC2",
    x"3626C27",
    x"362698C",
    x"36266F2",
    x"3626459",
    x"36261C0",
    x"3625F28",
    x"3625C90",
    x"36259FA",
    x"3625763",
    x"36254CE",
    x"3625239",
    x"3624FA5",
    x"3624D11",
    x"3624A7E",
    x"36247EC",
    x"362455A",
    x"36242C9",
    x"3624039",
    x"3623DA9",
    x"3623B1A",
    x"362388C",
    x"36235FE",
    x"3623371",
    x"36230E4",
    x"3622E58",
    x"3622BCD",
    x"3622942",
    x"36226B8",
    x"362242F",
    x"36221A6",
    x"3621F1E",
    x"3621C97",
    x"3621A10",
    x"3621789",
    x"3621504",
    x"362127F",
    x"3620FFB",
    x"3620D77",
    x"3620AF4",
    x"3620872",
    x"36205F0",
    x"362036F",
    x"36200EE",
    x"361FE6E",
    x"361FBEF",
    x"361F970",
    x"361F6F2",
    x"361F475",
    x"361F1F8",
    x"361EF7C",
    x"361ED00",
    x"361EA85",
    x"361E80B",
    x"361E591",
    x"361E318",
    x"361E0A0",
    x"361DE28",
    x"361DBB1",
    x"361D93A",
    x"361D6C4",
    x"361D44F",
    x"361D1DA",
    x"361CF66",
    x"361CCF2",
    x"361CA7F",
    x"361C80D",
    x"361C59B",
    x"361C32A",
    x"361C0BA",
    x"361BE4A",
    x"361BBDA",
    x"361B96C",
    x"361B6FE",
    x"361B490",
    x"361B223",
    x"361AFB7",
    x"361AD4C",
    x"361AAE0",
    x"361A876",
    x"361A60C",
    x"361A3A3",
    x"361A13A",
    x"3619ED2",
    x"3619C6B",
    x"3619A04",
    x"361979E",
    x"3619538",
    x"36192D3",
    x"361906F",
    x"3618E0B",
    x"3618BA8",
    x"3618945",
    x"36186E3",
    x"3618482",
    x"3618221",
    x"3617FC1",
    x"3617D61",
    x"3617B02",
    x"36178A4",
    x"3617646",
    x"36173E9",
    x"361718C",
    x"3616F30",
    x"3616CD4",
    x"3616A79",
    x"361681F",
    x"36165C5",
    x"361636C",
    x"3616114",
    x"3615EBC",
    x"3615C64",
    x"3615A0D",
    x"36157B7",
    x"3615562",
    x"361530D",
    x"36150B8",
    x"3614E64",
    x"3614C11",
    x"36149BE",
    x"361476C",
    x"361451A",
    x"36142C9",
    x"3614079",
    x"3613E29",
    x"3613BDA",
    x"361398B",
    x"361373D",
    x"36134F0",
    x"36132A3",
    x"3613056",
    x"3612E0B",
    x"3612BBF",
    x"3612975",
    x"361272B",
    x"36124E1",
    x"3612298",
    x"3612050",
    x"3611E08",
    x"3611BC1",
    x"361197A",
    x"3611734",
    x"36114EE",
    x"36112AA",
    x"3611065",
    x"3610E21",
    x"3610BDE",
    x"361099B",
    x"3610759",
    x"3610518",
    x"36102D7",
    x"3610096",
    x"360FE56",
    x"360FC17",
    x"360F9D8",
    x"360F79A",
    x"360F55D",
    x"360F320",
    x"360F0E3",
    x"360EEA7",
    x"360EC6C",
    x"360EA31",
    x"360E7F7",
    x"360E5BD",
    x"360E384",
    x"360E14B",
    x"360DF13",
    x"360DCDC",
    x"360DAA5",
    x"360D86E",
    x"360D638",
    x"360D403",
    x"360D1CE",
    x"360CF9A",
    x"360CD67",
    x"360CB34",
    x"360C901",
    x"360C6CF",
    x"360C49E",
    x"360C26D",
    x"360C03C",
    x"360BE0D",
    x"360BBDD",
    x"360B9AF",
    x"360B781",
    x"360B553",
    x"360B326",
    x"360B0F9",
    x"360AECD",
    x"360ACA2",
    x"360AA77",
    x"360A84D",
    x"360A623",
    x"360A3FA",
    x"360A1D1",
    x"3609FA9",
    x"3609D81",
    x"3609B5A",
    x"3609933",
    x"360970D",
    x"36094E8",
    x"36092C3",
    x"360909F",
    x"3608E7B",
    x"3608C57",
    x"3608A34",
    x"3608812",
    x"36085F0",
    x"36083CF",
    x"36081AF",
    x"3607F8E",
    x"3607D6F",
    x"3607B50",
    x"3607931",
    x"3607713",
    x"36074F6",
    x"36072D9",
    x"36070BC",
    x"3606EA0",
    x"3606C85",
    x"3606A6A",
    x"3606850",
    x"3606636",
    x"360641C",
    x"3606204",
    x"3605FEB",
    x"3605DD4",
    x"3605BBD",
    x"36059A6",
    x"3605790",
    x"360557A",
    x"3605365",
    x"3605150",
    x"3604F3C",
    x"3604D29",
    x"3604B16",
    x"3604903",
    x"36046F1",
    x"36044E0",
    x"36042CF",
    x"36040BE",
    x"3603EAE",
    x"3603C9F",
    x"3603A90",
    x"3603882",
    x"3603674",
    x"3603467",
    x"360325A",
    x"360304D",
    x"3602E42",
    x"3602C36",
    x"3602A2B",
    x"3602821",
    x"3602617",
    x"360240E",
    x"3602205",
    x"3601FFD",
    x"3601DF5",
    x"3601BEE",
    x"36019E7",
    x"36017E1",
    x"36015DB",
    x"36013D6",
    x"36011D1",
    x"3600FCD",
    x"3600DCA",
    x"3600BC6",
    x"36009C4",
    x"36007C2",
    x"36005C0",
    x"36003BF",
    x"36001BE",
    x"35FFF7C",
    x"35FFB7D",
    x"35FF77E",
    x"35FF381",
    x"35FEF85",
    x"35FEB89",
    x"35FE78F",
    x"35FE395",
    x"35FDF9D",
    x"35FDBA6",
    x"35FD7AF",
    x"35FD3BA",
    x"35FCFC5",
    x"35FCBD2",
    x"35FC7DF",
    x"35FC3EE",
    x"35FBFFD",
    x"35FBC0E",
    x"35FB81F",
    x"35FB432",
    x"35FB045",
    x"35FAC5A",
    x"35FA86F",
    x"35FA485",
    x"35FA09D",
    x"35F9CB5",
    x"35F98CE",
    x"35F94E9",
    x"35F9104",
    x"35F8D20",
    x"35F893D",
    x"35F855C",
    x"35F817B",
    x"35F7D9B",
    x"35F79BC",
    x"35F75DE",
    x"35F7201",
    x"35F6E25",
    x"35F6A4A",
    x"35F6670",
    x"35F6297",
    x"35F5EBF",
    x"35F5AE7",
    x"35F5711",
    x"35F533C",
    x"35F4F67",
    x"35F4B94",
    x"35F47C2",
    x"35F43F0",
    x"35F4020",
    x"35F3C50",
    x"35F3882",
    x"35F34B4",
    x"35F30E7",
    x"35F2D1B",
    x"35F2951",
    x"35F2587",
    x"35F21BE",
    x"35F1DF6",
    x"35F1A2F",
    x"35F1669",
    x"35F12A4",
    x"35F0EE0",
    x"35F0B1C",
    x"35F075A",
    x"35F0399",
    x"35EFFD8",
    x"35EFC19",
    x"35EF85A",
    x"35EF49C",
    x"35EF0E0",
    x"35EED24",
    x"35EE969",
    x"35EE5AF",
    x"35EE1F6",
    x"35EDE3E",
    x"35EDA87",
    x"35ED6D1",
    x"35ED31C",
    x"35ECF68",
    x"35ECBB4",
    x"35EC802",
    x"35EC450",
    x"35EC0A0",
    x"35EBCF0",
    x"35EB941",
    x"35EB593",
    x"35EB1E6",
    x"35EAE3A",
    x"35EAA8F",
    x"35EA6E5",
    x"35EA33C",
    x"35E9F93",
    x"35E9BEC",
    x"35E9845",
    x"35E94A0",
    x"35E90FB",
    x"35E8D57",
    x"35E89B4",
    x"35E8612",
    x"35E8271",
    x"35E7ED1",
    x"35E7B32",
    x"35E7794",
    x"35E73F6",
    x"35E705A",
    x"35E6CBE",
    x"35E6923",
    x"35E6589",
    x"35E61F0",
    x"35E5E58",
    x"35E5AC1",
    x"35E572B",
    x"35E5396",
    x"35E5001",
    x"35E4C6E",
    x"35E48DB",
    x"35E4549",
    x"35E41B8",
    x"35E3E28",
    x"35E3A99",
    x"35E370B",
    x"35E337E",
    x"35E2FF1",
    x"35E2C66",
    x"35E28DB",
    x"35E2551",
    x"35E21C9",
    x"35E1E41",
    x"35E1AB9",
    x"35E1733",
    x"35E13AE",
    x"35E1029",
    x"35E0CA6",
    x"35E0923",
    x"35E05A1",
    x"35E0220",
    x"35DFEA0",
    x"35DFB21",
    x"35DF7A3",
    x"35DF425",
    x"35DF0A8",
    x"35DED2D",
    x"35DE9B2",
    x"35DE638",
    x"35DE2BF",
    x"35DDF46",
    x"35DDBCF",
    x"35DD859",
    x"35DD4E3",
    x"35DD16E",
    x"35DCDFA",
    x"35DCA87",
    x"35DC715",
    x"35DC3A4",
    x"35DC033",
    x"35DBCC4",
    x"35DB955",
    x"35DB5E7",
    x"35DB27A",
    x"35DAF0E",
    x"35DABA2",
    x"35DA838",
    x"35DA4CE",
    x"35DA165",
    x"35D9DFD",
    x"35D9A96",
    x"35D9730",
    x"35D93CB",
    x"35D9066",
    x"35D8D03",
    x"35D89A0",
    x"35D863E",
    x"35D82DD",
    x"35D7F7C",
    x"35D7C1D",
    x"35D78BE",
    x"35D7561",
    x"35D7204",
    x"35D6EA8",
    x"35D6B4C",
    x"35D67F2",
    x"35D6498",
    x"35D6140",
    x"35D5DE8",
    x"35D5A91",
    x"35D573A",
    x"35D53E5",
    x"35D5090",
    x"35D4D3D",
    x"35D49EA",
    x"35D4698",
    x"35D4347",
    x"35D3FF6",
    x"35D3CA7",
    x"35D3958",
    x"35D360A",
    x"35D32BD",
    x"35D2F71",
    x"35D2C25",
    x"35D28DA",
    x"35D2591",
    x"35D2248",
    x"35D1EFF",
    x"35D1BB8",
    x"35D1872",
    x"35D152C",
    x"35D11E7",
    x"35D0EA3",
    x"35D0B60",
    x"35D081D",
    x"35D04DC",
    x"35D019B",
    x"35CFE5B",
    x"35CFB1C",
    x"35CF7DD",
    x"35CF4A0",
    x"35CF163",
    x"35CEE27",
    x"35CEAEC",
    x"35CE7B2",
    x"35CE478",
    x"35CE13F",
    x"35CDE07",
    x"35CDAD0",
    x"35CD79A",
    x"35CD465",
    x"35CD130",
    x"35CCDFC",
    x"35CCAC9",
    x"35CC797",
    x"35CC465",
    x"35CC134",
    x"35CBE04",
    x"35CBAD5",
    x"35CB7A7",
    x"35CB47A",
    x"35CB14D",
    x"35CAE21",
    x"35CAAF6",
    x"35CA7CB",
    x"35CA4A2",
    x"35CA179",
    x"35C9E51",
    x"35C9B2A",
    x"35C9803",
    x"35C94DE",
    x"35C91B9",
    x"35C8E95",
    x"35C8B72",
    x"35C884F",
    x"35C852E",
    x"35C820D",
    x"35C7EED",
    x"35C7BCD",
    x"35C78AF",
    x"35C7591",
    x"35C7274",
    x"35C6F58",
    x"35C6C3C",
    x"35C6922",
    x"35C6608",
    x"35C62EF",
    x"35C5FD6",
    x"35C5CBF",
    x"35C59A8",
    x"35C5692",
    x"35C537D",
    x"35C5068",
    x"35C4D54",
    x"35C4A41",
    x"35C472F",
    x"35C441E",
    x"35C410D",
    x"35C3DFD",
    x"35C3AEE",
    x"35C37E0",
    x"35C34D2",
    x"35C31C5",
    x"35C2EB9",
    x"35C2BAE",
    x"35C28A3",
    x"35C259A",
    x"35C2291",
    x"35C1F88",
    x"35C1C81",
    x"35C197A",
    x"35C1674",
    x"35C136F",
    x"35C106A",
    x"35C0D67",
    x"35C0A64",
    x"35C0762",
    x"35C0460",
    x"35C015F",
    x"35BFE5F",
    x"35BFB60",
    x"35BF862",
    x"35BF564",
    x"35BF267",
    x"35BEF6B",
    x"35BEC6F",
    x"35BE975",
    x"35BE67B",
    x"35BE381",
    x"35BE089",
    x"35BDD91",
    x"35BDA9A",
    x"35BD7A4",
    x"35BD4AE",
    x"35BD1B9",
    x"35BCEC5",
    x"35BCBD2",
    x"35BC8DF",
    x"35BC5EE",
    x"35BC2FC",
    x"35BC00C",
    x"35BBD1C",
    x"35BBA2E",
    x"35BB73F",
    x"35BB452",
    x"35BB165",
    x"35BAE79",
    x"35BAB8E",
    x"35BA8A3",
    x"35BA5BA",
    x"35BA2D1",
    x"35B9FE8",
    x"35B9D01",
    x"35B9A1A",
    x"35B9734",
    x"35B944E",
    x"35B9169",
    x"35B8E85",
    x"35B8BA2",
    x"35B88C0",
    x"35B85DE",
    x"35B82FD",
    x"35B801C",
    x"35B7D3D",
    x"35B7A5E",
    x"35B777F",
    x"35B74A2",
    x"35B71C5",
    x"35B6EE9",
    x"35B6C0E",
    x"35B6933",
    x"35B6659",
    x"35B6380",
    x"35B60A7",
    x"35B5DCF",
    x"35B5AF8",
    x"35B5822",
    x"35B554C",
    x"35B5277",
    x"35B4FA3",
    x"35B4CD0",
    x"35B49FD",
    x"35B472B",
    x"35B4459",
    x"35B4188",
    x"35B3EB8",
    x"35B3BE9",
    x"35B391A",
    x"35B364C",
    x"35B337F",
    x"35B30B3",
    x"35B2DE7",
    x"35B2B1C",
    x"35B2851",
    x"35B2588",
    x"35B22BF",
    x"35B1FF6",
    x"35B1D2F",
    x"35B1A68",
    x"35B17A1",
    x"35B14DC",
    x"35B1217",
    x"35B0F53",
    x"35B0C8F",
    x"35B09CC",
    x"35B070A",
    x"35B0449",
    x"35B0188",
    x"35AFEC8",
    x"35AFC09",
    x"35AF94A",
    x"35AF68C",
    x"35AF3CF",
    x"35AF112",
    x"35AEE56",
    x"35AEB9B",
    x"35AE8E1",
    x"35AE627",
    x"35AE36D",
    x"35AE0B5",
    x"35ADDFD",
    x"35ADB46",
    x"35AD88F",
    x"35AD5DA",
    x"35AD325",
    x"35AD070",
    x"35ACDBC",
    x"35ACB09",
    x"35AC857",
    x"35AC5A5",
    x"35AC2F4",
    x"35AC044",
    x"35ABD94",
    x"35ABAE5",
    x"35AB836",
    x"35AB589",
    x"35AB2DC",
    x"35AB02F",
    x"35AAD84",
    x"35AAAD8",
    x"35AA82E",
    x"35AA584",
    x"35AA2DB",
    x"35AA033",
    x"35A9D8B",
    x"35A9AE4",
    x"35A983E",
    x"35A9598",
    x"35A92F3",
    x"35A904F",
    x"35A8DAB",
    x"35A8B08",
    x"35A8865",
    x"35A85C4",
    x"35A8322",
    x"35A8082",
    x"35A7DE2",
    x"35A7B43",
    x"35A78A5",
    x"35A7607",
    x"35A736A",
    x"35A70CD",
    x"35A6E31",
    x"35A6B96",
    x"35A68FB",
    x"35A6661",
    x"35A63C8",
    x"35A6130",
    x"35A5E98",
    x"35A5C00",
    x"35A596A",
    x"35A56D4",
    x"35A543E",
    x"35A51A9",
    x"35A4F15",
    x"35A4C82",
    x"35A49EF",
    x"35A475D",
    x"35A44CB",
    x"35A423B",
    x"35A3FAA",
    x"35A3D1B",
    x"35A3A8C",
    x"35A37FD",
    x"35A3570",
    x"35A32E3",
    x"35A3056",
    x"35A2DCB",
    x"35A2B3F",
    x"35A28B5",
    x"35A262B",
    x"35A23A2",
    x"35A2119",
    x"35A1E91",
    x"35A1C0A",
    x"35A1983",
    x"35A16FD",
    x"35A1478",
    x"35A11F3",
    x"35A0F6F",
    x"35A0CEB",
    x"35A0A68",
    x"35A07E6",
    x"35A0564",
    x"35A02E3",
    x"35A0063",
    x"359FDE3",
    x"359FB64",
    x"359F8E5",
    x"359F668",
    x"359F3EA",
    x"359F16E",
    x"359EEF2",
    x"359EC76",
    x"359E9FB",
    x"359E781",
    x"359E508",
    x"359E28F",
    x"359E016",
    x"359DD9F",
    x"359DB27",
    x"359D8B1",
    x"359D63B",
    x"359D3C6",
    x"359D151",
    x"359CEDD",
    x"359CC6A",
    x"359C9F7",
    x"359C785",
    x"359C513",
    x"359C2A2",
    x"359C032",
    x"359BDC2",
    x"359BB53",
    x"359B8E4",
    x"359B677",
    x"359B409",
    x"359B19D",
    x"359AF30",
    x"359ACC5",
    x"359AA5A",
    x"359A7F0",
    x"359A586",
    x"359A31D",
    x"359A0B5",
    x"3599E4D",
    x"3599BE5",
    x"359997F",
    x"3599719",
    x"35994B3",
    x"359924E",
    x"3598FEA",
    x"3598D86",
    x"3598B23",
    x"35988C1",
    x"359865F",
    x"35983FE",
    x"359819D",
    x"3597F3D",
    x"3597CDD",
    x"3597A7E",
    x"3597820",
    x"35975C2",
    x"3597365",
    x"3597109",
    x"3596EAD",
    x"3596C51",
    x"35969F6",
    x"359679C",
    x"3596543",
    x"35962EA",
    x"3596091",
    x"3595E39",
    x"3595BE2",
    x"359598B",
    x"3595735",
    x"35954E0",
    x"359528B",
    x"3595037",
    x"3594DE3",
    x"3594B90",
    x"359493D",
    x"35946EB",
    x"3594499",
    x"3594249",
    x"3593FF8",
    x"3593DA9",
    x"3593B5A",
    x"359390B",
    x"35936BD",
    x"3593470",
    x"3593223",
    x"3592FD7",
    x"3592D8B",
    x"3592B40",
    x"35928F5",
    x"35926AB",
    x"3592462",
    x"3592219",
    x"3591FD1",
    x"3591D89",
    x"3591B42",
    x"35918FC",
    x"35916B6",
    x"3591470",
    x"359122B",
    x"3590FE7",
    x"3590DA3",
    x"3590B60",
    x"359091E",
    x"35906DC",
    x"359049A",
    x"3590259",
    x"3590019",
    x"358FDD9",
    x"358FB9A",
    x"358F95C",
    x"358F71E",
    x"358F4E0",
    x"358F2A3",
    x"358F067",
    x"358EE2B",
    x"358EBF0",
    x"358E9B5",
    x"358E77B",
    x"358E541",
    x"358E308",
    x"358E0D0",
    x"358DE98",
    x"358DC60",
    x"358DA2A",
    x"358D7F3",
    x"358D5BE",
    x"358D388",
    x"358D154",
    x"358CF20",
    x"358CCEC",
    x"358CAB9",
    x"358C887",
    x"358C655",
    x"358C424",
    x"358C1F3",
    x"358BFC3",
    x"358BD93",
    x"358BB64",
    x"358B935",
    x"358B707",
    x"358B4DA",
    x"358B2AD",
    x"358B081",
    x"358AE55",
    x"358AC29",
    x"358A9FF",
    x"358A7D4",
    x"358A5AB",
    x"358A382",
    x"358A159",
    x"3589F31",
    x"3589D09",
    x"3589AE2",
    x"35898BC",
    x"3589696",
    x"3589471",
    x"358924C",
    x"3589027",
    x"3588E04",
    x"3588BE0",
    x"35889BE",
    x"358879C",
    x"358857A",
    x"3588359",
    x"3588138",
    x"3587F18",
    x"3587CF9",
    x"3587ADA",
    x"35878BB",
    x"358769D",
    x"3587480",
    x"3587263",
    x"3587047",
    x"3586E2B",
    x"3586C10",
    x"35869F5",
    x"35867DB",
    x"35865C1",
    x"35863A8",
    x"358618F",
    x"3585F77",
    x"3585D5F",
    x"3585B48",
    x"3585932",
    x"358571C",
    x"3585506",
    x"35852F1",
    x"35850DD",
    x"3584EC9",
    x"3584CB5",
    x"3584AA2",
    x"3584890",
    x"358467E",
    x"358446D",
    x"358425C",
    x"358404C",
    x"3583E3C",
    x"3583C2C",
    x"3583A1E",
    x"358380F",
    x"3583602",
    x"35833F4",
    x"35831E8",
    x"3582FDB",
    x"3582DD0",
    x"3582BC5",
    x"35829BA",
    x"35827B0",
    x"35825A6",
    x"358239D",
    x"3582194",
    x"3581F8C",
    x"3581D84",
    x"3581B7D",
    x"3581977",
    x"3581771",
    x"358156B",
    x"3581366",
    x"3581161",
    x"3580F5D",
    x"3580D5A",
    x"3580B57",
    x"3580954",
    x"3580752",
    x"3580550",
    x"358034F",
    x"358014F",
    x"357FE9E",
    x"357FA9E",
    x"357F6A0",
    x"357F2A3",
    x"357EEA7",
    x"357EAAC",
    x"357E6B2",
    x"357E2B8",
    x"357DEC0",
    x"357DAC9",
    x"357D6D3",
    x"357D2DE",
    x"357CEE9",
    x"357CAF6",
    x"357C704",
    x"357C313",
    x"357BF22",
    x"357BB33",
    x"357B745",
    x"357B357",
    x"357AF6B",
    x"357AB80",
    x"357A795",
    x"357A3AC",
    x"3579FC4",
    x"3579BDC",
    x"35797F6",
    x"3579410",
    x"357902C",
    x"3578C48",
    x"3578865",
    x"3578484",
    x"35780A3",
    x"3577CC3",
    x"35778E5",
    x"3577507",
    x"357712A",
    x"3576D4E",
    x"3576974",
    x"357659A",
    x"35761C1",
    x"3575DE9",
    x"3575A12",
    x"357563C",
    x"3575267",
    x"3574E93",
    x"3574ABF",
    x"35746ED",
    x"357431C",
    x"3573F4C",
    x"3573B7C",
    x"35737AE",
    x"35733E0",
    x"3573014",
    x"3572C48",
    x"357287E",
    x"35724B4",
    x"35720EB",
    x"3571D24",
    x"357195D",
    x"3571597",
    x"35711D2",
    x"3570E0E",
    x"3570A4B",
    x"3570689",
    x"35702C8",
    x"356FF08",
    x"356FB48",
    x"356F78A",
    x"356F3CD",
    x"356F010",
    x"356EC55",
    x"356E89A",
    x"356E4E0",
    x"356E127",
    x"356DD70",
    x"356D9B9",
    x"356D603",
    x"356D24E",
    x"356CE9A",
    x"356CAE6",
    x"356C734",
    x"356C383",
    x"356BFD2",
    x"356BC23",
    x"356B874",
    x"356B4C7",
    x"356B11A",
    x"356AD6E",
    x"356A9C3",
    x"356A619",
    x"356A270",
    x"3569EC8",
    x"3569B21",
    x"356977A",
    x"35693D5",
    x"3569031",
    x"3568C8D",
    x"35688EA",
    x"3568548",
    x"35681A8",
    x"3567E08",
    x"3567A69",
    x"35676CA",
    x"356732D",
    x"3566F91",
    x"3566BF5",
    x"356685B",
    x"35664C1",
    x"3566129",
    x"3565D91",
    x"35659FA",
    x"3565664",
    x"35652CF",
    x"3564F3A",
    x"3564BA7",
    x"3564814",
    x"3564483",
    x"35640F2",
    x"3563D62",
    x"35639D3",
    x"3563645",
    x"35632B8",
    x"3562F2C",
    x"3562BA1",
    x"3562816",
    x"356248D",
    x"3562104",
    x"3561D7C",
    x"35619F5",
    x"356166F",
    x"35612EA",
    x"3560F66",
    x"3560BE2",
    x"3560860",
    x"35604DE",
    x"356015D",
    x"355FDDD",
    x"355FA5E",
    x"355F6E0",
    x"355F363",
    x"355EFE7",
    x"355EC6B",
    x"355E8F0",
    x"355E577",
    x"355E1FE",
    x"355DE86",
    x"355DB0E",
    x"355D798",
    x"355D423",
    x"355D0AE",
    x"355CD3A",
    x"355C9C7",
    x"355C655",
    x"355C2E4",
    x"355BF74",
    x"355BC04",
    x"355B896",
    x"355B528",
    x"355B1BB",
    x"355AE4F",
    x"355AAE4",
    x"355A77A",
    x"355A410",
    x"355A0A8",
    x"3559D40",
    x"35599D9",
    x"3559673",
    x"355930E",
    x"3558FAA",
    x"3558C46",
    x"35588E4",
    x"3558582",
    x"3558221",
    x"3557EC1",
    x"3557B61",
    x"3557803",
    x"35574A5",
    x"3557149",
    x"3556DED",
    x"3556A92",
    x"3556737",
    x"35563DE",
    x"3556086",
    x"3555D2E",
    x"35559D7",
    x"3555681",
    x"355532C",
    x"3554FD7",
    x"3554C84",
    x"3554931",
    x"35545DF",
    x"355428E",
    x"3553F3E",
    x"3553BEE",
    x"35538A0",
    x"3553552",
    x"3553205",
    x"3552EB9",
    x"3552B6E",
    x"3552823",
    x"35524DA",
    x"3552191",
    x"3551E49",
    x"3551B02",
    x"35517BC",
    x"3551476",
    x"3551131",
    x"3550DED",
    x"3550AAA",
    x"3550768",
    x"3550427",
    x"35500E6",
    x"354FDA6",
    x"354FA67",
    x"354F729",
    x"354F3EC",
    x"354F0AF",
    x"354ED73",
    x"354EA38",
    x"354E6FE",
    x"354E3C5",
    x"354E08C",
    x"354DD55",
    x"354DA1E",
    x"354D6E7",
    x"354D3B2",
    x"354D07E",
    x"354CD4A",
    x"354CA17",
    x"354C6E5",
    x"354C3B4",
    x"354C083",
    x"354BD53",
    x"354BA24",
    x"354B6F6",
    x"354B3C9",
    x"354B09C",
    x"354AD71",
    x"354AA46",
    x"354A71B",
    x"354A3F2",
    x"354A0C9",
    x"3549DA2",
    x"3549A7B",
    x"3549754",
    x"354942F",
    x"354910A",
    x"3548DE6",
    x"3548AC3",
    x"35487A1",
    x"3548480",
    x"354815F",
    x"3547E3F",
    x"3547B20",
    x"3547801",
    x"35474E4",
    x"35471C7",
    x"3546EAB",
    x"3546B8F",
    x"3546875",
    x"354655B",
    x"3546242",
    x"3545F2A",
    x"3545C13",
    x"35458FC",
    x"35455E6",
    x"35452D1",
    x"3544FBD",
    x"3544CA9",
    x"3544996",
    x"3544684",
    x"3544373",
    x"3544063",
    x"3543D53",
    x"3543A44",
    x"3543736",
    x"3543428",
    x"354311C",
    x"3542E10",
    x"3542B05",
    x"35427FA",
    x"35424F1",
    x"35421E8",
    x"3541EE0",
    x"3541BD9",
    x"35418D2",
    x"35415CC",
    x"35412C7",
    x"3540FC3",
    x"3540CBF",
    x"35409BC",
    x"35406BA",
    x"35403B9",
    x"35400B8",
    x"353FDB9",
    x"353FABA",
    x"353F7BB",
    x"353F4BE",
    x"353F1C1",
    x"353EEC5",
    x"353EBC9",
    x"353E8CF",
    x"353E5D5",
    x"353E2DC",
    x"353DFE4",
    x"353DCEC",
    x"353D9F5",
    x"353D6FF",
    x"353D40A",
    x"353D115",
    x"353CE21",
    x"353CB2E",
    x"353C83C",
    x"353C54A",
    x"353C259",
    x"353BF69",
    x"353BC79",
    x"353B98A",
    x"353B69C",
    x"353B3AF",
    x"353B0C3",
    x"353ADD7",
    x"353AAEC",
    x"353A801",
    x"353A518",
    x"353A22F",
    x"3539F47",
    x"3539C5F",
    x"3539978",
    x"3539692",
    x"35393AD",
    x"35390C9",
    x"3538DE5",
    x"3538B02",
    x"353881F",
    x"353853E",
    x"353825D",
    x"3537F7C",
    x"3537C9D",
    x"35379BE",
    x"35376E0",
    x"3537403",
    x"3537126",
    x"3536E4A",
    x"3536B6F",
    x"3536894",
    x"35365BB",
    x"35362E1",
    x"3536009",
    x"3535D31",
    x"3535A5A",
    x"3535784",
    x"35354AF",
    x"35351DA",
    x"3534F06",
    x"3534C32",
    x"3534960",
    x"353468E",
    x"35343BC",
    x"35340EC",
    x"3533E1C",
    x"3533B4D",
    x"353387E",
    x"35335B1",
    x"35332E3",
    x"3533017",
    x"3532D4B",
    x"3532A80",
    x"35327B6",
    x"35324ED",
    x"3532224",
    x"3531F5C",
    x"3531C94",
    x"35319CD",
    x"3531707",
    x"3531442",
    x"353117D",
    x"3530EB9",
    x"3530BF6",
    x"3530933",
    x"3530671",
    x"35303B0",
    x"35300EF",
    x"352FE2F",
    x"352FB70",
    x"352F8B2",
    x"352F5F4",
    x"352F337",
    x"352F07A",
    x"352EDBE",
    x"352EB03",
    x"352E849",
    x"352E58F",
    x"352E2D6",
    x"352E01E",
    x"352DD66",
    x"352DAAF",
    x"352D7F9",
    x"352D543",
    x"352D28E",
    x"352CFDA",
    x"352CD26",
    x"352CA73",
    x"352C7C1",
    x"352C50F",
    x"352C25E",
    x"352BFAE",
    x"352BCFF",
    x"352BA50",
    x"352B7A1",
    x"352B4F4",
    x"352B247",
    x"352AF9B",
    x"352ACEF",
    x"352AA44",
    x"352A79A",
    x"352A4F0",
    x"352A247",
    x"3529F9F",
    x"3529CF8",
    x"3529A51",
    x"35297AA",
    x"3529505",
    x"3529260",
    x"3528FBC",
    x"3528D18",
    x"3528A75",
    x"35287D3",
    x"3528531",
    x"3528290",
    x"3527FF0",
    x"3527D50",
    x"3527AB1",
    x"3527813",
    x"3527575",
    x"35272D8",
    x"352703C",
    x"3526DA0",
    x"3526B05",
    x"352686B",
    x"35265D1",
    x"3526338",
    x"352609F",
    x"3525E07",
    x"3525B70",
    x"35258DA",
    x"3525644",
    x"35253AF",
    x"352511A",
    x"3524E86",
    x"3524BF3",
    x"3524960",
    x"35246CE",
    x"352443D",
    x"35241AC",
    x"3523F1C",
    x"3523C8C",
    x"35239FD",
    x"352376F",
    x"35234E2",
    x"3523255",
    x"3522FC9",
    x"3522D3D",
    x"3522AB2",
    x"3522828",
    x"352259E",
    x"3522315",
    x"352208C",
    x"3521E05",
    x"3521B7D",
    x"35218F7",
    x"3521671",
    x"35213EC",
    x"3521167",
    x"3520EE3",
    x"3520C5F",
    x"35209DD",
    x"352075B",
    x"35204D9",
    x"3520258",
    x"351FFD8",
    x"351FD58",
    x"351FAD9",
    x"351F85B",
    x"351F5DD",
    x"351F360",
    x"351F0E3",
    x"351EE67",
    x"351EBEC",
    x"351E971",
    x"351E6F7",
    x"351E47E",
    x"351E205",
    x"351DF8D",
    x"351DD15",
    x"351DA9E",
    x"351D828",
    x"351D5B2",
    x"351D33D",
    x"351D0C9",
    x"351CE55",
    x"351CBE2",
    x"351C96F",
    x"351C6FD",
    x"351C48B",
    x"351C21B",
    x"351BFAA",
    x"351BD3B",
    x"351BACC",
    x"351B85D",
    x"351B5F0",
    x"351B382",
    x"351B116",
    x"351AEAA",
    x"351AC3E",
    x"351A9D4",
    x"351A76A",
    x"351A500",
    x"351A297",
    x"351A02F",
    x"3519DC7",
    x"3519B60",
    x"35198F9",
    x"3519693",
    x"351942E",
    x"35191C9",
    x"3518F65",
    x"3518D01",
    x"3518A9F",
    x"351883C",
    x"35185DA",
    x"3518379",
    x"3518119",
    x"3517EB9",
    x"3517C59",
    x"35179FB",
    x"351779C",
    x"351753F",
    x"35172E2",
    x"3517085",
    x"3516E29",
    x"3516BCE",
    x"3516974",
    x"3516719",
    x"35164C0",
    x"3516267",
    x"351600F",
    x"3515DB7",
    x"3515B60",
    x"3515909",
    x"35156B3",
    x"351545E",
    x"3515209",
    x"3514FB5",
    x"3514D61",
    x"3514B0E",
    x"35148BC",
    x"351466A",
    x"3514419",
    x"35141C8",
    x"3513F78",
    x"3513D28",
    x"3513AD9",
    x"351388B",
    x"351363D",
    x"35133F0",
    x"35131A3",
    x"3512F57",
    x"3512D0B",
    x"3512AC0",
    x"3512876",
    x"351262C",
    x"35123E3",
    x"351219A",
    x"3511F52",
    x"3511D0A",
    x"3511AC3",
    x"351187D",
    x"3511637",
    x"35113F2",
    x"35111AD",
    x"3510F69",
    x"3510D26",
    x"3510AE3",
    x"35108A0",
    x"351065E",
    x"351041D",
    x"35101DC",
    x"350FF9C",
    x"350FD5C",
    x"350FB1D",
    x"350F8DF",
    x"350F6A1",
    x"350F463",
    x"350F227",
    x"350EFEA",
    x"350EDAF",
    x"350EB74",
    x"350E939",
    x"350E6FF",
    x"350E4C5",
    x"350E28D",
    x"350E054",
    x"350DE1C",
    x"350DBE5",
    x"350D9AE",
    x"350D778",
    x"350D543",
    x"350D30E",
    x"350D0D9",
    x"350CEA5",
    x"350CC72",
    x"350CA3F",
    x"350C80D",
    x"350C5DB",
    x"350C3AA",
    x"350C179",
    x"350BF49",
    x"350BD1A",
    x"350BAEB",
    x"350B8BC",
    x"350B68E",
    x"350B461",
    x"350B234",
    x"350B008",
    x"350ADDC",
    x"350ABB1",
    x"350A986",
    x"350A75C",
    x"350A532",
    x"350A309",
    x"350A0E1",
    x"3509EB9",
    x"3509C92",
    x"3509A6B",
    x"3509844",
    x"350961F",
    x"35093F9",
    x"35091D5",
    x"3508FB0",
    x"3508D8D",
    x"3508B6A",
    x"3508947",
    x"3508725",
    x"3508503",
    x"35082E2",
    x"35080C2",
    x"3507EA2",
    x"3507C83",
    x"3507A64",
    x"3507845",
    x"3507628",
    x"350740A",
    x"35071EE",
    x"3506FD1",
    x"3506DB6",
    x"3506B9B",
    x"3506980",
    x"3506766",
    x"350654C",
    x"3506333",
    x"350611B",
    x"3505F03",
    x"3505CEB",
    x"3505AD4",
    x"35058BE",
    x"35056A8",
    x"3505492",
    x"350527D",
    x"3505069",
    x"3504E55",
    x"3504C42",
    x"3504A2F",
    x"350481D",
    x"350460B",
    x"35043FA",
    x"35041E9",
    x"3503FD9",
    x"3503DC9",
    x"3503BBA",
    x"35039AB",
    x"350379D",
    x"3503590",
    x"3503382",
    x"3503176",
    x"3502F6A",
    x"3502D5E",
    x"3502B53",
    x"3502948",
    x"350273E",
    x"3502535",
    x"350232C",
    x"3502123",
    x"3501F1B",
    x"3501D14",
    x"3501B0D",
    x"3501906",
    x"3501700",
    x"35014FB",
    x"35012F6",
    x"35010F1",
    x"3500EED",
    x"3500CEA",
    x"3500AE7",
    x"35008E4",
    x"35006E2",
    x"35004E1",
    x"35002E0",
    x"35000DF",
    x"34FFDBF",
    x"34FF9C0",
    x"34FF5C2",
    x"34FF1C5",
    x"34FEDC9",
    x"34FE9CE",
    x"34FE5D4",
    x"34FE1DC",
    x"34FDDE4",
    x"34FD9ED",
    x"34FD5F7",
    x"34FD202",
    x"34FCE0E",
    x"34FCA1B",
    x"34FC629",
    x"34FC237",
    x"34FBE47",
    x"34FBA58",
    x"34FB66A",
    x"34FB27D",
    x"34FAE91",
    x"34FAAA6",
    x"34FA6BC",
    x"34FA2D2",
    x"34F9EEA",
    x"34F9B03",
    x"34F971D",
    x"34F9337",
    x"34F8F53",
    x"34F8B70",
    x"34F878D",
    x"34F83AC",
    x"34F7FCC",
    x"34F7BEC",
    x"34F780E",
    x"34F7430",
    x"34F7054",
    x"34F6C78",
    x"34F689D",
    x"34F64C4",
    x"34F60EB",
    x"34F5D13",
    x"34F593C",
    x"34F5567",
    x"34F5192",
    x"34F4DBE",
    x"34F49EB",
    x"34F4619",
    x"34F4248",
    x"34F3E78",
    x"34F3AA9",
    x"34F36DA",
    x"34F330D",
    x"34F2F41",
    x"34F2B75",
    x"34F27AB",
    x"34F23E2",
    x"34F2019",
    x"34F1C52",
    x"34F188B",
    x"34F14C5",
    x"34F1101",
    x"34F0D3D",
    x"34F097A",
    x"34F05B8",
    x"34F01F7",
    x"34EFE37",
    x"34EFA78",
    x"34EF6BA",
    x"34EF2FD",
    x"34EEF40",
    x"34EEB85",
    x"34EE7CB",
    x"34EE411",
    x"34EE059",
    x"34EDCA1",
    x"34ED8EA",
    x"34ED534",
    x"34ED180",
    x"34ECDCC",
    x"34ECA19",
    x"34EC667",
    x"34EC2B6",
    x"34EBF05",
    x"34EBB56",
    x"34EB7A8",
    x"34EB3FA",
    x"34EB04E",
    x"34EACA2",
    x"34EA8F7",
    x"34EA54E",
    x"34EA1A5",
    x"34E9DFD",
    x"34E9A56",
    x"34E96B0",
    x"34E930A",
    x"34E8F66",
    x"34E8BC3",
    x"34E8820",
    x"34E847F",
    x"34E80DE",
    x"34E7D3E",
    x"34E799F",
    x"34E7601",
    x"34E7264",
    x"34E6EC8",
    x"34E6B2D",
    x"34E6793",
    x"34E63F9",
    x"34E6061",
    x"34E5CC9",
    x"34E5932",
    x"34E559C",
    x"34E5207",
    x"34E4E73",
    x"34E4AE0",
    x"34E474E",
    x"34E43BC",
    x"34E402C",
    x"34E3C9C",
    x"34E390E",
    x"34E3580",
    x"34E31F3",
    x"34E2E67",
    x"34E2ADC",
    x"34E2751",
    x"34E23C8",
    x"34E2040",
    x"34E1CB8",
    x"34E1931",
    x"34E15AB",
    x"34E1226",
    x"34E0EA2",
    x"34E0B1F",
    x"34E079D",
    x"34E041B",
    x"34E009B",
    x"34DFD1B",
    x"34DF99C",
    x"34DF61E",
    x"34DF2A1",
    x"34DEF25",
    x"34DEBA9",
    x"34DE82F",
    x"34DE4B5",
    x"34DE13D",
    x"34DDDC5",
    x"34DDA4E",
    x"34DD6D8",
    x"34DD362",
    x"34DCFEE",
    x"34DCC7A",
    x"34DC908",
    x"34DC596",
    x"34DC225",
    x"34DBEB5",
    x"34DBB46",
    x"34DB7D7",
    x"34DB46A",
    x"34DB0FD",
    x"34DAD91",
    x"34DAA26",
    x"34DA6BC",
    x"34DA353",
    x"34D9FEA",
    x"34D9C83",
    x"34D991C",
    x"34D95B6",
    x"34D9251",
    x"34D8EED",
    x"34D8B8A",
    x"34D8827",
    x"34D84C6",
    x"34D8165",
    x"34D7E05",
    x"34D7AA6",
    x"34D7748",
    x"34D73EA",
    x"34D708E",
    x"34D6D32",
    x"34D69D7",
    x"34D667D",
    x"34D6324",
    x"34D5FCC",
    x"34D5C74",
    x"34D591D",
    x"34D55C7",
    x"34D5272",
    x"34D4F1E",
    x"34D4BCB",
    x"34D4878",
    x"34D4527",
    x"34D41D6",
    x"34D3E86",
    x"34D3B36",
    x"34D37E8",
    x"34D349B",
    x"34D314E",
    x"34D2E02",
    x"34D2AB7",
    x"34D276D",
    x"34D2423",
    x"34D20DA",
    x"34D1D93",
    x"34D1A4C",
    x"34D1705",
    x"34D13C0",
    x"34D107C",
    x"34D0D38",
    x"34D09F5",
    x"34D06B3",
    x"34D0372",
    x"34D0031",
    x"34CFCF2",
    x"34CF9B3",
    x"34CF675",
    x"34CF337",
    x"34CEFFB",
    x"34CECBF",
    x"34CE985",
    x"34CE64B",
    x"34CE312",
    x"34CDFD9",
    x"34CDCA2",
    x"34CD96B",
    x"34CD635",
    x"34CD300",
    x"34CCFCB",
    x"34CCC98",
    x"34CC965",
    x"34CC633",
    x"34CC302",
    x"34CBFD2",
    x"34CBCA2",
    x"34CB973",
    x"34CB645",
    x"34CB318",
    x"34CAFEC",
    x"34CACC0",
    x"34CA995",
    x"34CA66B",
    x"34CA342",
    x"34CA01A",
    x"34C9CF2",
    x"34C99CB",
    x"34C96A5",
    x"34C9380",
    x"34C905C",
    x"34C8D38",
    x"34C8A15",
    x"34C86F3",
    x"34C83D1",
    x"34C80B1",
    x"34C7D91",
    x"34C7A72",
    x"34C7754",
    x"34C7436",
    x"34C711A",
    x"34C6DFE",
    x"34C6AE3",
    x"34C67C8",
    x"34C64AF",
    x"34C6196",
    x"34C5E7E",
    x"34C5B67",
    x"34C5850",
    x"34C553B",
    x"34C5226",
    x"34C4F12",
    x"34C4BFE",
    x"34C48EC",
    x"34C45DA",
    x"34C42C9",
    x"34C3FB8",
    x"34C3CA9",
    x"34C399A",
    x"34C368C",
    x"34C337F",
    x"34C3072",
    x"34C2D67",
    x"34C2A5C",
    x"34C2751",
    x"34C2448",
    x"34C213F",
    x"34C1E37",
    x"34C1B30",
    x"34C182A",
    x"34C1524",
    x"34C121F",
    x"34C0F1B",
    x"34C0C18",
    x"34C0915",
    x"34C0613",
    x"34C0312",
    x"34C0012",
    x"34BFD12",
    x"34BFA13",
    x"34BF715",
    x"34BF417",
    x"34BF11B",
    x"34BEE1F",
    x"34BEB24",
    x"34BE829",
    x"34BE530",
    x"34BE237",
    x"34BDF3F",
    x"34BDC47",
    x"34BD950",
    x"34BD65A",
    x"34BD365",
    x"34BD071",
    x"34BCD7D",
    x"34BCA8A",
    x"34BC798",
    x"34BC4A6",
    x"34BC1B5",
    x"34BBEC5",
    x"34BBBD6",
    x"34BB8E7",
    x"34BB5FA",
    x"34BB30C",
    x"34BB020",
    x"34BAD34",
    x"34BAA49",
    x"34BA75F",
    x"34BA476",
    x"34BA18D",
    x"34B9EA5",
    x"34B9BBE",
    x"34B98D7",
    x"34B95F1",
    x"34B930C",
    x"34B9028",
    x"34B8D44",
    x"34B8A61",
    x"34B877F",
    x"34B849D",
    x"34B81BD",
    x"34B7EDC",
    x"34B7BFD",
    x"34B791E",
    x"34B7641",
    x"34B7363",
    x"34B7087",
    x"34B6DAB",
    x"34B6AD0",
    x"34B67F6",
    x"34B651C",
    x"34B6243",
    x"34B5F6B",
    x"34B5C93",
    x"34B59BD",
    x"34B56E7",
    x"34B5411",
    x"34B513D",
    x"34B4E69",
    x"34B4B95",
    x"34B48C3",
    x"34B45F1",
    x"34B4320",
    x"34B404F",
    x"34B3D80",
    x"34B3AB1",
    x"34B37E2",
    x"34B3515",
    x"34B3248",
    x"34B2F7C",
    x"34B2CB0",
    x"34B29E5",
    x"34B271B",
    x"34B2452",
    x"34B2189",
    x"34B1EC1",
    x"34B1BFA",
    x"34B1933",
    x"34B166D",
    x"34B13A8",
    x"34B10E3",
    x"34B0E1F",
    x"34B0B5C",
    x"34B089A",
    x"34B05D8",
    x"34B0317",
    x"34B0056",
    x"34AFD96",
    x"34AFAD7",
    x"34AF819",
    x"34AF55B",
    x"34AF29E",
    x"34AEFE2",
    x"34AED26",
    x"34AEA6B",
    x"34AE7B1",
    x"34AE4F8",
    x"34AE23F",
    x"34ADF86",
    x"34ADCCF",
    x"34ADA18",
    x"34AD762",
    x"34AD4AC",
    x"34AD1F8",
    x"34ACF43",
    x"34ACC90",
    x"34AC9DD",
    x"34AC72B",
    x"34AC47A",
    x"34AC1C9",
    x"34ABF19",
    x"34ABC69",
    x"34AB9BA",
    x"34AB70C",
    x"34AB45F",
    x"34AB1B2",
    x"34AAF06",
    x"34AAC5B",
    x"34AA9B0",
    x"34AA706",
    x"34AA45C",
    x"34AA1B4",
    x"34A9F0C",
    x"34A9C64",
    x"34A99BD",
    x"34A9717",
    x"34A9472",
    x"34A91CD",
    x"34A8F29",
    x"34A8C85",
    x"34A89E3",
    x"34A8740",
    x"34A849F",
    x"34A81FE",
    x"34A7F5E",
    x"34A7CBE",
    x"34A7A20",
    x"34A7781",
    x"34A74E4",
    x"34A7247",
    x"34A6FAB",
    x"34A6D0F",
    x"34A6A74",
    x"34A67DA",
    x"34A6540",
    x"34A62A7",
    x"34A600F",
    x"34A5D77",
    x"34A5AE0",
    x"34A584A",
    x"34A55B4",
    x"34A531F",
    x"34A508A",
    x"34A4DF7",
    x"34A4B63",
    x"34A48D1",
    x"34A463F",
    x"34A43AE",
    x"34A411D",
    x"34A3E8D",
    x"34A3BFE",
    x"34A396F",
    x"34A36E1",
    x"34A3454",
    x"34A31C7",
    x"34A2F3B",
    x"34A2CAF",
    x"34A2A25",
    x"34A279A",
    x"34A2511",
    x"34A2288",
    x"34A2000",
    x"34A1D78",
    x"34A1AF1",
    x"34A186A",
    x"34A15E5",
    x"34A135F",
    x"34A10DB",
    x"34A0E57",
    x"34A0BD4",
    x"34A0951",
    x"34A06CF",
    x"34A044E",
    x"34A01CD",
    x"349FF4D",
    x"349FCCD",
    x"349FA4E",
    x"349F7D0",
    x"349F552",
    x"349F2D5",
    x"349F059",
    x"349EDDD",
    x"349EB62",
    x"349E8E8",
    x"349E66E",
    x"349E3F4",
    x"349E17C",
    x"349DF04",
    x"349DC8C",
    x"349DA15",
    x"349D79F",
    x"349D52A",
    x"349D2B5",
    x"349D040",
    x"349CDCC",
    x"349CB59",
    x"349C8E7",
    x"349C675",
    x"349C404",
    x"349C193",
    x"349BF23",
    x"349BCB3",
    x"349BA44",
    x"349B7D6",
    x"349B568",
    x"349B2FB",
    x"349B08F",
    x"349AE23",
    x"349ABB8",
    x"349A94D",
    x"349A6E3",
    x"349A47A",
    x"349A211",
    x"3499FA9",
    x"3499D41",
    x"3499ADA",
    x"3499874",
    x"349960E",
    x"34993A9",
    x"3499144",
    x"3498EE0",
    x"3498C7D",
    x"3498A1A",
    x"34987B8",
    x"3498556",
    x"34982F5",
    x"3498095",
    x"3497E35",
    x"3497BD5",
    x"3497977",
    x"3497719",
    x"34974BB",
    x"349725E",
    x"3497002",
    x"3496DA6",
    x"3496B4B",
    x"34968F1",
    x"3496697",
    x"349643D",
    x"34961E5",
    x"3495F8C",
    x"3495D35",
    x"3495ADE",
    x"3495887",
    x"3495632",
    x"34953DC",
    x"3495188",
    x"3494F34",
    x"3494CE0",
    x"3494A8D",
    x"349483B",
    x"34945E9",
    x"3494398",
    x"3494147",
    x"3493EF7",
    x"3493CA8",
    x"3493A59",
    x"349380B",
    x"34935BD",
    x"3493370",
    x"3493123",
    x"3492ED7",
    x"3492C8C",
    x"3492A41",
    x"34927F7",
    x"34925AD",
    x"3492364",
    x"349211B",
    x"3491ED3",
    x"3491C8C",
    x"3491A45",
    x"34917FF",
    x"34915B9",
    x"3491374",
    x"349112F",
    x"3490EEB",
    x"3490CA8",
    x"3490A65",
    x"3490822",
    x"34905E1",
    x"34903A0",
    x"349015F",
    x"348FF1F",
    x"348FCDF",
    x"348FAA0",
    x"348F862",
    x"348F624",
    x"348F3E7",
    x"348F1AA",
    x"348EF6E",
    x"348ED33",
    x"348EAF8",
    x"348E8BD",
    x"348E683",
    x"348E44A",
    x"348E211",
    x"348DFD9",
    x"348DDA1",
    x"348DB6A",
    x"348D933",
    x"348D6FD",
    x"348D4C8",
    x"348D293",
    x"348D05F",
    x"348CE2B",
    x"348CBF8",
    x"348C9C5",
    x"348C793",
    x"348C561",
    x"348C330",
    x"348C0FF",
    x"348BECF",
    x"348BCA0",
    x"348BA71",
    x"348B843",
    x"348B615",
    x"348B3E8",
    x"348B1BB",
    x"348AF8F",
    x"348AD63",
    x"348AB38",
    x"348A90E",
    x"348A6E4",
    x"348A4BA",
    x"348A291",
    x"348A069",
    x"3489E41",
    x"3489C1A",
    x"34899F3",
    x"34897CD",
    x"34895A7",
    x"3489382",
    x"348915D",
    x"3488F39",
    x"3488D16",
    x"3488AF3",
    x"34888D0",
    x"34886AE",
    x"348848D",
    x"348826C",
    x"348804C",
    x"3487E2C",
    x"3487C0D",
    x"34879EE",
    x"34877D0",
    x"34875B2",
    x"3487395",
    x"3487178",
    x"3486F5C",
    x"3486D41",
    x"3486B25",
    x"348690B",
    x"34866F1",
    x"34864D7",
    x"34862BF",
    x"34860A6",
    x"3485E8E",
    x"3485C77",
    x"3485A60",
    x"348584A",
    x"3485634",
    x"348541F",
    x"348520A",
    x"3484FF6",
    x"3484DE2",
    x"3484BCF",
    x"34849BC",
    x"34847AA",
    x"3484598",
    x"3484387",
    x"3484176",
    x"3483F66",
    x"3483D57",
    x"3483B48",
    x"3483939",
    x"348372B",
    x"348351D",
    x"3483310",
    x"3483104",
    x"3482EF8",
    x"3482CEC",
    x"3482AE1",
    x"34828D7",
    x"34826CD",
    x"34824C3",
    x"34822BB",
    x"34820B2",
    x"3481EAA",
    x"3481CA3",
    x"3481A9C",
    x"3481895",
    x"3481690",
    x"348148A",
    x"3481285",
    x"3481081",
    x"3480E7D",
    x"3480C7A",
    x"3480A77",
    x"3480874",
    x"3480673",
    x"3480471",
    x"3480270",
    x"3480070",
    x"347FCE1",
    x"347F8E2",
    x"347F4E4",
    x"347F0E8",
    x"347ECEC",
    x"347E8F1",
    x"347E4F7",
    x"347E0FF",
    x"347DD07",
    x"347D910",
    x"347D51A",
    x"347D126",
    x"347CD32",
    x"347C93F",
    x"347C54D",
    x"347C15C",
    x"347BD6D",
    x"347B97E",
    x"347B590",
    x"347B1A3",
    x"347ADB7",
    x"347A9CC",
    x"347A5E2",
    x"347A1F9",
    x"3479E11",
    x"3479A2A",
    x"3479644",
    x"347925F",
    x"3478E7B",
    x"3478A98",
    x"34786B5",
    x"34782D4",
    x"3477EF4",
    x"3477B15",
    x"3477737",
    x"3477359",
    x"3476F7D",
    x"3476BA1",
    x"34767C7",
    x"34763EE",
    x"3476015",
    x"3475C3E",
    x"3475867",
    x"3475491",
    x"34750BD",
    x"3474CE9",
    x"3474916",
    x"3474544",
    x"3474174",
    x"3473DA4",
    x"34739D5",
    x"3473607",
    x"347323A",
    x"3472E6E",
    x"3472AA3",
    x"34726D8",
    x"347230F",
    x"3471F47",
    x"3471B7F",
    x"34717B9",
    x"34713F4",
    x"347102F",
    x"3470C6C",
    x"34708A9",
    x"34704E7",
    x"3470126",
    x"346FD67",
    x"346F9A8",
    x"346F5EA",
    x"346F22D",
    x"346EE71",
    x"346EAB6",
    x"346E6FB",
    x"346E342",
    x"346DF8A",
    x"346DBD2",
    x"346D81C",
    x"346D466",
    x"346D0B2",
    x"346CCFE",
    x"346C94B",
    x"346C599",
    x"346C1E8",
    x"346BE38",
    x"346BA89",
    x"346B6DB",
    x"346B32E",
    x"346AF81",
    x"346ABD6",
    x"346A82B",
    x"346A482",
    x"346A0D9",
    x"3469D31",
    x"346998B",
    x"34695E5",
    x"3469240",
    x"3468E9C",
    x"3468AF8",
    x"3468756",
    x"34683B5",
    x"3468014",
    x"3467C75",
    x"34678D6",
    x"3467538",
    x"346719B",
    x"3466DFF",
    x"3466A64",
    x"34666CA",
    x"3466331",
    x"3465F99",
    x"3465C01",
    x"346586B",
    x"34654D5",
    x"3465140",
    x"3464DAC",
    x"3464A19",
    x"3464687",
    x"34642F6",
    x"3463F66",
    x"3463BD6",
    x"3463848",
    x"34634BA",
    x"346312E",
    x"3462DA2",
    x"3462A17",
    x"346268D",
    x"3462303",
    x"3461F7B",
    x"3461BF4",
    x"346186D",
    x"34614E8",
    x"3461163",
    x"3460DDF",
    x"3460A5C",
    x"34606DA",
    x"3460358",
    x"345FFD8",
    x"345FC58",
    x"345F8DA",
    x"345F55C",
    x"345F1DF",
    x"345EE63",
    x"345EAE8",
    x"345E76E",
    x"345E3F4",
    x"345E07C",
    x"345DD04",
    x"345D98D",
    x"345D617",
    x"345D2A2",
    x"345CF2E",
    x"345CBBA",
    x"345C848",
    x"345C4D6",
    x"345C166",
    x"345BDF6",
    x"345BA87",
    x"345B718",
    x"345B3AB",
    x"345B03F",
    x"345ACD3",
    x"345A968",
    x"345A5FE",
    x"345A295",
    x"3459F2D",
    x"3459BC6",
    x"345985F",
    x"34594F9",
    x"3459195",
    x"3458E31",
    x"3458ACD",
    x"345876B",
    x"345840A",
    x"34580A9",
    x"3457D49",
    x"34579EB",
    x"345768C",
    x"345732F",
    x"3456FD3",
    x"3456C77",
    x"345691D",
    x"34565C3",
    x"345626A",
    x"3455F12",
    x"3455BBA",
    x"3455864",
    x"345550E",
    x"34551B9",
    x"3454E65",
    x"3454B12",
    x"34547C0",
    x"345446E",
    x"345411D",
    x"3453DCE",
    x"3453A7E",
    x"3453730",
    x"34533E3",
    x"3453096",
    x"3452D4B",
    x"3452A00",
    x"34526B6",
    x"345236C",
    x"3452024",
    x"3451CDC",
    x"3451995",
    x"345164F",
    x"345130A",
    x"3450FC6",
    x"3450C82",
    x"3450940",
    x"34505FE",
    x"34502BD",
    x"344FF7C",
    x"344FC3D",
    x"344F8FE",
    x"344F5C0",
    x"344F283",
    x"344EF47",
    x"344EC0C",
    x"344E8D1",
    x"344E597",
    x"344E25E",
    x"344DF26",
    x"344DBEF",
    x"344D8B8",
    x"344D582",
    x"344D24D",
    x"344CF19",
    x"344CBE6",
    x"344C8B3",
    x"344C582",
    x"344C251",
    x"344BF20",
    x"344BBF1",
    x"344B8C2",
    x"344B595",
    x"344B268",
    x"344AF3B",
    x"344AC10",
    x"344A8E5",
    x"344A5BC",
    x"344A293",
    x"3449F6A",
    x"3449C43",
    x"344991C",
    x"34495F6",
    x"34492D1",
    x"3448FAD",
    x"3448C89",
    x"3448967",
    x"3448645",
    x"3448323",
    x"3448003",
    x"3447CE3",
    x"34479C5",
    x"34476A7",
    x"3447389",
    x"344706D",
    x"3446D51",
    x"3446A36",
    x"344671C",
    x"3446403",
    x"34460EA",
    x"3445DD2",
    x"3445ABB",
    x"34457A5",
    x"344548F",
    x"344517A",
    x"3444E66",
    x"3444B53",
    x"3444841",
    x"344452F",
    x"344421E",
    x"3443F0E",
    x"3443BFF",
    x"34438F0",
    x"34435E2",
    x"34432D5",
    x"3442FC9",
    x"3442CBD",
    x"34429B2",
    x"34426A8",
    x"344239F",
    x"3442097",
    x"3441D8F",
    x"3441A88",
    x"3441782",
    x"344147C",
    x"3441177",
    x"3440E73",
    x"3440B70",
    x"344086E",
    x"344056C",
    x"344026B",
    x"343FF6B",
    x"343FC6B",
    x"343F96C",
    x"343F66E",
    x"343F371",
    x"343F075",
    x"343ED79",
    x"343EA7E",
    x"343E784",
    x"343E48A",
    x"343E191",
    x"343DE99",
    x"343DBA2",
    x"343D8AC",
    x"343D5B6",
    x"343D2C1",
    x"343CFCC",
    x"343CCD9",
    x"343C9E6",
    x"343C6F4",
    x"343C403",
    x"343C112",
    x"343BE22",
    x"343BB33",
    x"343B844",
    x"343B557",
    x"343B26A",
    x"343AF7E",
    x"343AC92",
    x"343A9A7",
    x"343A6BD",
    x"343A3D4",
    x"343A0EB",
    x"3439E03",
    x"3439B1C",
    x"3439836",
    x"3439550",
    x"343926B",
    x"3438F87",
    x"3438CA3",
    x"34389C1",
    x"34386DF",
    x"34383FD",
    x"343811D",
    x"3437E3D",
    x"3437B5D",
    x"343787F",
    x"34375A1",
    x"34372C4",
    x"3436FE8",
    x"3436D0C",
    x"3436A31",
    x"3436757",
    x"343647E",
    x"34361A5",
    x"3435ECD",
    x"3435BF5",
    x"343591F",
    x"3435649",
    x"3435374",
    x"343509F",
    x"3434DCB",
    x"3434AF8",
    x"3434826",
    x"3434554",
    x"3434283",
    x"3433FB3",
    x"3433CE3",
    x"3433A14",
    x"3433746",
    x"3433479",
    x"34331AC",
    x"3432EE0",
    x"3432C15",
    x"343294A",
    x"3432680",
    x"34323B7",
    x"34320EE",
    x"3431E26",
    x"3431B5F",
    x"3431899",
    x"34315D3",
    x"343130E",
    x"3431049",
    x"3430D85",
    x"3430AC2",
    x"3430800",
    x"343053E",
    x"343027D",
    x"342FFBD",
    x"342FCFE",
    x"342FA3F",
    x"342F780",
    x"342F4C3",
    x"342F206",
    x"342EF4A",
    x"342EC8E",
    x"342E9D4",
    x"342E71A",
    x"342E460",
    x"342E1A7",
    x"342DEEF",
    x"342DC38",
    x"342D981",
    x"342D6CB",
    x"342D416",
    x"342D161",
    x"342CEAD",
    x"342CBFA",
    x"342C947",
    x"342C695",
    x"342C3E4",
    x"342C133",
    x"342BE83",
    x"342BBD4",
    x"342B925",
    x"342B677",
    x"342B3CA",
    x"342B11D",
    x"342AE71",
    x"342ABC6",
    x"342A91C",
    x"342A672",
    x"342A3C8",
    x"342A120",
    x"3429E78",
    x"3429BD1",
    x"342992A",
    x"3429684",
    x"34293DF",
    x"342913A",
    x"3428E96",
    x"3428BF3",
    x"3428950",
    x"34286AE",
    x"342840D",
    x"342816C",
    x"3427ECC",
    x"3427C2D",
    x"342798E",
    x"34276F0",
    x"3427452",
    x"34271B6",
    x"3426F1A",
    x"3426C7E",
    x"34269E3",
    x"3426749",
    x"34264B0",
    x"3426217",
    x"3425F7F",
    x"3425CE7",
    x"3425A50",
    x"34257BA",
    x"3425524",
    x"342528F",
    x"3424FFB",
    x"3424D67",
    x"3424AD4",
    x"3424842",
    x"34245B0",
    x"342431F",
    x"342408F",
    x"3423DFF",
    x"3423B70",
    x"34238E1",
    x"3423653",
    x"34233C6",
    x"3423139",
    x"3422EAD",
    x"3422C22",
    x"3422997",
    x"342270D",
    x"3422484",
    x"34221FB",
    x"3421F73",
    x"3421CEB",
    x"3421A64",
    x"34217DE",
    x"3421558",
    x"34212D3",
    x"342104F",
    x"3420DCB",
    x"3420B48",
    x"34208C6",
    x"3420644",
    x"34203C2",
    x"3420142",
    x"341FEC2",
    x"341FC42",
    x"341F9C4",
    x"341F746",
    x"341F4C8",
    x"341F24B",
    x"341EFCF",
    x"341ED53",
    x"341EAD8",
    x"341E85E",
    x"341E5E4",
    x"341E36B",
    x"341E0F2",
    x"341DE7A",
    x"341DC03",
    x"341D98C",
    x"341D716",
    x"341D4A1",
    x"341D22C",
    x"341CFB8",
    x"341CD44",
    x"341CAD1",
    x"341C85F",
    x"341C5ED",
    x"341C37C",
    x"341C10B",
    x"341BE9B",
    x"341BC2C",
    x"341B9BD",
    x"341B74F",
    x"341B4E1",
    x"341B275",
    x"341B008",
    x"341AD9D",
    x"341AB31",
    x"341A8C7",
    x"341A65D",
    x"341A3F4",
    x"341A18B",
    x"3419F23",
    x"3419CBC",
    x"3419A55",
    x"34197EE",
    x"3419589",
    x"3419324",
    x"34190BF",
    x"3418E5B",
    x"3418BF8",
    x"3418995",
    x"3418733",
    x"34184D2",
    x"3418271",
    x"3418010",
    x"3417DB1",
    x"3417B52",
    x"34178F3",
    x"3417695",
    x"3417438",
    x"34171DB",
    x"3416F7F",
    x"3416D23",
    x"3416AC8",
    x"341686E",
    x"3416614",
    x"34163BB",
    x"3416162",
    x"3415F0A",
    x"3415CB3",
    x"3415A5C",
    x"3415805",
    x"34155B0",
    x"341535B",
    x"3415106",
    x"3414EB2",
    x"3414C5F",
    x"3414A0C",
    x"34147BA",
    x"3414568",
    x"3414317",
    x"34140C6",
    x"3413E77",
    x"3413C27",
    x"34139D9",
    x"341378A",
    x"341353D",
    x"34132F0",
    x"34130A3",
    x"3412E57",
    x"3412C0C",
    x"34129C1",
    x"3412777",
    x"341252E",
    x"34122E5",
    x"341209C",
    x"3411E54",
    x"3411C0D",
    x"34119C6",
    x"3411780",
    x"341153B",
    x"34112F6",
    x"34110B1",
    x"3410E6D",
    x"3410C2A",
    x"34109E7",
    x"34107A5",
    x"3410563",
    x"3410322",
    x"34100E2",
    x"340FEA2",
    x"340FC62",
    x"340FA24",
    x"340F7E5",
    x"340F5A8",
    x"340F36A",
    x"340F12E",
    x"340EEF2",
    x"340ECB6",
    x"340EA7C",
    x"340E841",
    x"340E607",
    x"340E3CE",
    x"340E195",
    x"340DF5D",
    x"340DD26",
    x"340DAEF",
    x"340D8B8",
    x"340D682",
    x"340D44D",
    x"340D218",
    x"340CFE4",
    x"340CDB0",
    x"340CB7D",
    x"340C94B",
    x"340C719",
    x"340C4E7",
    x"340C2B6",
    x"340C086",
    x"340BE56",
    x"340BC27",
    x"340B9F8",
    x"340B7CA",
    x"340B59C",
    x"340B36F",
    x"340B142",
    x"340AF16",
    x"340ACEB",
    x"340AAC0",
    x"340A895",
    x"340A66B",
    x"340A442",
    x"340A219",
    x"3409FF1",
    x"3409DC9",
    x"3409BA2",
    x"340997B",
    x"3409755",
    x"3409530",
    x"340930B",
    x"34090E6",
    x"3408EC2",
    x"3408C9F",
    x"3408A7C",
    x"340885A",
    x"3408638",
    x"3408417",
    x"34081F6",
    x"3407FD6",
    x"3407DB6",
    x"3407B97",
    x"3407978",
    x"340775A",
    x"340753C",
    x"340731F",
    x"3407103",
    x"3406EE7",
    x"3406CCB",
    x"3406AB0",
    x"3406896",
    x"340667C",
    x"3406463",
    x"340624A",
    x"3406032",
    x"3405E1A",
    x"3405C03",
    x"34059EC",
    x"34057D6",
    x"34055C0",
    x"34053AB",
    x"3405196",
    x"3404F82",
    x"3404D6E",
    x"3404B5B",
    x"3404949",
    x"3404737",
    x"3404525",
    x"3404314",
    x"3404103",
    x"3403EF3",
    x"3403CE4",
    x"3403AD5",
    x"34038C7",
    x"34036B9",
    x"34034AB",
    x"340329E",
    x"3403092",
    x"3402E86",
    x"3402C7B",
    x"3402A70",
    x"3402865",
    x"340265C",
    x"3402452",
    x"3402249",
    x"3402041",
    x"3401E39",
    x"3401C32",
    x"3401A2B",
    x"3401825",
    x"340161F",
    x"340141A",
    x"3401215",
    x"3401011",
    x"3400E0D",
    x"3400C0A",
    x"3400A07",
    x"3400805",
    x"3400603",
    x"3400402",
    x"3400201",
    x"3400001",
    x"33FFC02",
    x"33FF804",
    x"33FF406",
    x"33FF00A",
    x"33FEC0E",
    x"33FE814",
    x"33FE41A",
    x"33FE022",
    x"33FDC2A",
    x"33FD834",
    x"33FD43E",
    x"33FD04A",
    x"33FCC56",
    x"33FC864",
    x"33FC472",
    x"33FC081",
    x"33FBC92",
    x"33FB8A3",
    x"33FB4B5",
    x"33FB0C9",
    x"33FACDD",
    x"33FA8F2",
    x"33FA508",
    x"33FA120",
    x"33F9D38",
    x"33F9951",
    x"33F956B",
    x"33F9186",
    x"33F8DA2",
    x"33F89C0",
    x"33F85DE",
    x"33F81FD",
    x"33F7E1D",
    x"33F7A3E",
    x"33F765F",
    x"33F7282",
    x"33F6EA6",
    x"33F6ACB",
    x"33F66F1",
    x"33F6318",
    x"33F5F3F",
    x"33F5B68",
    x"33F5792",
    x"33F53BC",
    x"33F4FE8",
    x"33F4C14",
    x"33F4842",
    x"33F4470",
    x"33F409F",
    x"33F3CD0",
    x"33F3901",
    x"33F3533",
    x"33F3166",
    x"33F2D9B",
    x"33F29D0",
    x"33F2606",
    x"33F223D",
    x"33F1E75",
    x"33F1AAD",
    x"33F16E7",
    x"33F1322",
    x"33F0F5E",
    x"33F0B9A",
    x"33F07D8",
    x"33F0416",
    x"33F0056",
    x"33EFC96",
    x"33EF8D7",
    x"33EF51A",
    x"33EF15D",
    x"33EEDA1",
    x"33EE9E6",
    x"33EE62C",
    x"33EE273",
    x"33EDEBB",
    x"33EDB04",
    x"33ED74D",
    x"33ED398",
    x"33ECFE4",
    x"33ECC30",
    x"33EC87D",
    x"33EC4CC",
    x"33EC11B",
    x"33EBD6B",
    x"33EB9BC",
    x"33EB60E",
    x"33EB261",
    x"33EAEB5",
    x"33EAB0A",
    x"33EA760",
    x"33EA3B6",
    x"33EA00E",
    x"33E9C66",
    x"33E98C0",
    x"33E951A",
    x"33E9175",
    x"33E8DD1",
    x"33E8A2E",
    x"33E868C",
    x"33E82EB",
    x"33E7F4B",
    x"33E7BAB",
    x"33E780D",
    x"33E746F",
    x"33E70D3",
    x"33E6D37",
    x"33E699C",
    x"33E6602",
    x"33E6269",
    x"33E5ED1",
    x"33E5B3A",
    x"33E57A3",
    x"33E540E",
    x"33E5079",
    x"33E4CE5",
    x"33E4953",
    x"33E45C1",
    x"33E4230",
    x"33E3EA0",
    x"33E3B11",
    x"33E3782",
    x"33E33F5",
    x"33E3068",
    x"33E2CDD",
    x"33E2952",
    x"33E25C8",
    x"33E223F",
    x"33E1EB7",
    x"33E1B30",
    x"33E17A9",
    x"33E1424",
    x"33E109F",
    x"33E0D1B",
    x"33E0999",
    x"33E0617",
    x"33E0296",
    x"33DFF15",
    x"33DFB96",
    x"33DF818",
    x"33DF49A",
    x"33DF11D",
    x"33DEDA1",
    x"33DEA26",
    x"33DE6AC",
    x"33DE333",
    x"33DDFBB",
    x"33DDC43",
    x"33DD8CD",
    x"33DD557",
    x"33DD1E2",
    x"33DCE6E",
    x"33DCAFB",
    x"33DC788",
    x"33DC417",
    x"33DC0A6",
    x"33DBD37",
    x"33DB9C8",
    x"33DB65A",
    x"33DB2ED",
    x"33DAF80",
    x"33DAC15",
    x"33DA8AA",
    x"33DA540",
    x"33DA1D8",
    x"33D9E70",
    x"33D9B08",
    x"33D97A2",
    x"33D943D",
    x"33D90D8",
    x"33D8D74",
    x"33D8A11",
    x"33D86AF",
    x"33D834E",
    x"33D7FED",
    x"33D7C8E",
    x"33D792F",
    x"33D75D1",
    x"33D7274",
    x"33D6F18",
    x"33D6BBD",
    x"33D6862",
    x"33D6508",
    x"33D61B0",
    x"33D5E58",
    x"33D5B00",
    x"33D57AA",
    x"33D5455",
    x"33D5100",
    x"33D4DAC",
    x"33D4A59",
    x"33D4707",
    x"33D43B6",
    x"33D4065",
    x"33D3D15",
    x"33D39C7",
    x"33D3679",
    x"33D332B",
    x"33D2FDF",
    x"33D2C93",
    x"33D2949",
    x"33D25FF",
    x"33D22B6",
    x"33D1F6D",
    x"33D1C26",
    x"33D18DF",
    x"33D1599",
    x"33D1254",
    x"33D0F10",
    x"33D0BCD",
    x"33D088A",
    x"33D0549",
    x"33D0208",
    x"33CFEC8",
    x"33CFB88",
    x"33CF84A",
    x"33CF50C",
    x"33CF1CF",
    x"33CEE93",
    x"33CEB58",
    x"33CE81E",
    x"33CE4E4",
    x"33CE1AB",
    x"33CDE73",
    x"33CDB3C",
    x"33CD806",
    x"33CD4D0",
    x"33CD19B",
    x"33CCE67",
    x"33CCB34",
    x"33CC802",
    x"33CC4D0",
    x"33CC19F",
    x"33CBE6F",
    x"33CBB40",
    x"33CB812",
    x"33CB4E4",
    x"33CB1B7",
    x"33CAE8B",
    x"33CAB60",
    x"33CA835",
    x"33CA50C",
    x"33CA1E3",
    x"33C9EBB",
    x"33C9B93",
    x"33C986D",
    x"33C9547",
    x"33C9222",
    x"33C8EFE",
    x"33C8BDB",
    x"33C88B8",
    x"33C8596",
    x"33C8275",
    x"33C7F55",
    x"33C7C36",
    x"33C7917",
    x"33C75F9",
    x"33C72DC",
    x"33C6FC0",
    x"33C6CA4",
    x"33C6989",
    x"33C6670",
    x"33C6356",
    x"33C603E",
    x"33C5D26",
    x"33C5A0F",
    x"33C56F9",
    x"33C53E4",
    x"33C50CF",
    x"33C4DBB",
    x"33C4AA8",
    x"33C4796",
    x"33C4485",
    x"33C4174",
    x"33C3E64",
    x"33C3B55",
    x"33C3846",
    x"33C3538",
    x"33C322C",
    x"33C2F1F",
    x"33C2C14",
    x"33C2909",
    x"33C25FF",
    x"33C22F6",
    x"33C1FEE",
    x"33C1CE6",
    x"33C19DF",
    x"33C16D9",
    x"33C13D4",
    x"33C10CF",
    x"33C0DCC",
    x"33C0AC9",
    x"33C07C6",
    x"33C04C5",
    x"33C01C4",
    x"33BFEC4",
    x"33BFBC5",
    x"33BF8C6",
    x"33BF5C8",
    x"33BF2CB",
    x"33BEFCF",
    x"33BECD3",
    x"33BE9D8",
    x"33BE6DE",
    x"33BE3E5",
    x"33BE0EC",
    x"33BDDF4",
    x"33BDAFD",
    x"33BD807",
    x"33BD511",
    x"33BD21C",
    x"33BCF28",
    x"33BCC35",
    x"33BC942",
    x"33BC650",
    x"33BC35F",
    x"33BC06E",
    x"33BBD7F",
    x"33BBA90",
    x"33BB7A1",
    x"33BB4B4",
    x"33BB1C7",
    x"33BAEDB",
    x"33BABF0",
    x"33BA905",
    x"33BA61B",
    x"33BA332",
    x"33BA04A",
    x"33B9D62",
    x"33B9A7B",
    x"33B9795",
    x"33B94AF",
    x"33B91CA",
    x"33B8EE6",
    x"33B8C03",
    x"33B8920",
    x"33B863E",
    x"33B835D",
    x"33B807D",
    x"33B7D9D",
    x"33B7ABE",
    x"33B77DF",
    x"33B7502",
    x"33B7225",
    x"33B6F49",
    x"33B6C6D",
    x"33B6993",
    x"33B66B9",
    x"33B63DF",
    x"33B6107",
    x"33B5E2F",
    x"33B5B57",
    x"33B5881",
    x"33B55AB",
    x"33B52D6",
    x"33B5002",
    x"33B4D2E",
    x"33B4A5B",
    x"33B4789",
    x"33B44B7",
    x"33B41E7",
    x"33B3F16",
    x"33B3C47",
    x"33B3978",
    x"33B36AA",
    x"33B33DD",
    x"33B3110",
    x"33B2E44",
    x"33B2B79",
    x"33B28AF",
    x"33B25E5",
    x"33B231C",
    x"33B2053",
    x"33B1D8C",
    x"33B1AC5",
    x"33B17FE",
    x"33B1539",
    x"33B1274",
    x"33B0FAF",
    x"33B0CEC",
    x"33B0A29",
    x"33B0767",
    x"33B04A5",
    x"33B01E4",
    x"33AFF24",
    x"33AFC65",
    x"33AF9A6",
    x"33AF6E8",
    x"33AF42B",
    x"33AF16E",
    x"33AEEB2",
    x"33AEBF7",
    x"33AE93C",
    x"33AE682",
    x"33AE3C9",
    x"33AE110",
    x"33ADE58",
    x"33ADBA1",
    x"33AD8EA",
    x"33AD634",
    x"33AD37F",
    x"33AD0CB",
    x"33ACE17",
    x"33ACB64",
    x"33AC8B1",
    x"33AC5FF",
    x"33AC34E",
    x"33AC09E",
    x"33ABDEE",
    x"33ABB3F",
    x"33AB890",
    x"33AB5E2",
    x"33AB335",
    x"33AB089",
    x"33AADDD",
    x"33AAB32",
    x"33AA887",
    x"33AA5DE",
    x"33AA334",
    x"33AA08C",
    x"33A9DE4",
    x"33A9B3D",
    x"33A9897",
    x"33A95F1",
    x"33A934C",
    x"33A90A7",
    x"33A8E03",
    x"33A8B60",
    x"33A88BE",
    x"33A861C",
    x"33A837A",
    x"33A80DA",
    x"33A7E3A",
    x"33A7B9B",
    x"33A78FC",
    x"33A765E",
    x"33A73C1",
    x"33A7124",
    x"33A6E89",
    x"33A6BED",
    x"33A6953",
    x"33A66B9",
    x"33A641F",
    x"33A6186",
    x"33A5EEE",
    x"33A5C57",
    x"33A59C0",
    x"33A572A",
    x"33A5495",
    x"33A5200",
    x"33A4F6C",
    x"33A4CD8",
    x"33A4A45",
    x"33A47B3",
    x"33A4521",
    x"33A4290",
    x"33A4000",
    x"33A3D70",
    x"33A3AE1",
    x"33A3853",
    x"33A35C5",
    x"33A3338",
    x"33A30AC",
    x"33A2E20",
    x"33A2B95",
    x"33A290A",
    x"33A2680",
    x"33A23F7",
    x"33A216E",
    x"33A1EE6",
    x"33A1C5F",
    x"33A19D8",
    x"33A1752",
    x"33A14CC",
    x"33A1247",
    x"33A0FC3",
    x"33A0D3F",
    x"33A0ABC",
    x"33A083A",
    x"33A05B8",
    x"33A0337",
    x"33A00B7",
    x"339FE37",
    x"339FBB8",
    x"339F939",
    x"339F6BB",
    x"339F43E",
    x"339F1C1",
    x"339EF45",
    x"339ECC9",
    x"339EA4E",
    x"339E7D4",
    x"339E55A",
    x"339E2E1",
    x"339E069",
    x"339DDF1",
    x"339DB7A",
    x"339D903",
    x"339D68D",
    x"339D418",
    x"339D1A3",
    x"339CF2F",
    x"339CCBC",
    x"339CA49",
    x"339C7D7",
    x"339C565",
    x"339C2F4",
    x"339C084",
    x"339BE14",
    x"339BBA5",
    x"339B936",
    x"339B6C8",
    x"339B45B",
    x"339B1EE",
    x"339AF82",
    x"339AD16",
    x"339AAAB",
    x"339A841",
    x"339A5D7",
    x"339A36E",
    x"339A105",
    x"3399E9D",
    x"3399C36",
    x"33999CF",
    x"3399769",
    x"3399503",
    x"339929E",
    x"339903A",
    x"3398DD6",
    x"3398B73",
    x"3398911",
    x"33986AF",
    x"339844D",
    x"33981EC",
    x"3397F8C",
    x"3397D2D",
    x"3397ACE",
    x"339786F",
    x"3397611",
    x"33973B4",
    x"3397158",
    x"3396EFC",
    x"3396CA0",
    x"3396A45",
    x"33967EB",
    x"3396591",
    x"3396338",
    x"33960E0",
    x"3395E88",
    x"3395C30",
    x"33959DA",
    x"3395784",
    x"339552E",
    x"33952D9",
    x"3395085",
    x"3394E31",
    x"3394BDD",
    x"339498B",
    x"3394739",
    x"33944E7",
    x"3394296",
    x"3394046",
    x"3393DF6",
    x"3393BA7",
    x"3393958",
    x"339370A",
    x"33934BD",
    x"3393270",
    x"3393023",
    x"3392DD8",
    x"3392B8D",
    x"3392942",
    x"33926F8",
    x"33924AE",
    x"3392266",
    x"339201D",
    x"3391DD6",
    x"3391B8E",
    x"3391948",
    x"3391702",
    x"33914BC",
    x"3391277",
    x"3391033",
    x"3390DEF",
    x"3390BAC",
    x"3390969",
    x"3390727",
    x"33904E6",
    x"33902A5",
    x"3390065",
    x"338FE25",
    x"338FBE5",
    x"338F9A7",
    x"338F769",
    x"338F52B",
    x"338F2EE",
    x"338F0B2",
    x"338EE76",
    x"338EC3A",
    x"338EA00",
    x"338E7C5",
    x"338E58C",
    x"338E353",
    x"338E11A",
    x"338DEE2",
    x"338DCAB",
    x"338DA74",
    x"338D83D",
    x"338D608",
    x"338D3D2",
    x"338D19E",
    x"338CF6A",
    x"338CD36",
    x"338CB03",
    x"338C8D0",
    x"338C69E",
    x"338C46D",
    x"338C23C",
    x"338C00C",
    x"338BDDC",
    x"338BBAD",
    x"338B97E",
    x"338B750",
    x"338B523",
    x"338B2F6",
    x"338B0C9",
    x"338AE9D",
    x"338AC72",
    x"338AA47",
    x"338A81D",
    x"338A5F3",
    x"338A3CA",
    x"338A1A1",
    x"3389F79",
    x"3389D51",
    x"3389B2A",
    x"3389904",
    x"33896DE",
    x"33894B8",
    x"3389294",
    x"338906F",
    x"3388E4B",
    x"3388C28",
    x"3388A05",
    x"33887E3",
    x"33885C1",
    x"33883A0",
    x"338817F",
    x"3387F5F",
    x"3387D40",
    x"3387B21",
    x"3387902",
    x"33876E4",
    x"33874C7",
    x"33872AA",
    x"338708D",
    x"3386E72",
    x"3386C56",
    x"3386A3B",
    x"3386821",
    x"3386607",
    x"33863EE",
    x"33861D5",
    x"3385FBD",
    x"3385DA5",
    x"3385B8E",
    x"3385978",
    x"3385762",
    x"338554C",
    x"3385337",
    x"3385122",
    x"3384F0E",
    x"3384CFB",
    x"3384AE8",
    x"33848D5",
    x"33846C3",
    x"33844B2",
    x"33842A1",
    x"3384091",
    x"3383E81",
    x"3383C71",
    x"3383A63",
    x"3383854",
    x"3383646",
    x"3383439",
    x"338322C",
    x"3383020",
    x"3382E14",
    x"3382C09",
    x"33829FE",
    x"33827F4",
    x"33825EA",
    x"33823E1",
    x"33821D8",
    x"3381FD0",
    x"3381DC8",
    x"3381BC1",
    x"33819BB",
    x"33817B4",
    x"33815AF",
    x"33813AA",
    x"33811A5",
    x"3380FA1",
    x"3380D9D",
    x"3380B9A",
    x"3380997",
    x"3380795",
    x"3380593",
    x"3380392",
    x"3380192",
    x"337FF24",
    x"337FB24",
    x"337F726",
    x"337F329",
    x"337EF2C",
    x"337EB31",
    x"337E737",
    x"337E33D",
    x"337DF45",
    x"337DB4E",
    x"337D757",
    x"337D362",
    x"337CF6E",
    x"337CB7A",
    x"337C788",
    x"337C397",
    x"337BFA6",
    x"337BBB7",
    x"337B7C8",
    x"337B3DB",
    x"337AFEE",
    x"337AC03",
    x"337A818",
    x"337A42F",
    x"337A046",
    x"3379C5F",
    x"3379878",
    x"3379493",
    x"33790AE",
    x"3378CCA",
    x"33788E7",
    x"3378506",
    x"3378125",
    x"3377D45",
    x"3377966",
    x"3377588",
    x"33771AC",
    x"3376DD0",
    x"33769F5",
    x"337661B",
    x"3376242",
    x"3375E6A",
    x"3375A92",
    x"33756BC",
    x"33752E7",
    x"3374F13",
    x"3374B40",
    x"337476D",
    x"337439C",
    x"3373FCB",
    x"3373BFC",
    x"337382D",
    x"3373460",
    x"3373093",
    x"3372CC8",
    x"33728FD",
    x"3372533",
    x"337216A",
    x"3371DA2",
    x"33719DB",
    x"3371615",
    x"3371250",
    x"3370E8C",
    x"3370AC9",
    x"3370707",
    x"3370346",
    x"336FF85",
    x"336FBC6",
    x"336F807",
    x"336F44A",
    x"336F08D",
    x"336ECD1",
    x"336E917",
    x"336E55D",
    x"336E1A4",
    x"336DDEC",
    x"336DA35",
    x"336D67F",
    x"336D2CA",
    x"336CF16",
    x"336CB62",
    x"336C7B0",
    x"336C3FE",
    x"336C04E",
    x"336BC9E",
    x"336B8F0",
    x"336B542",
    x"336B195",
    x"336ADE9",
    x"336AA3E",
    x"336A694",
    x"336A2EB",
    x"3369F42",
    x"3369B9B",
    x"33697F5",
    x"336944F",
    x"33690AB",
    x"3368D07",
    x"3368964",
    x"33685C2",
    x"3368221",
    x"3367E81",
    x"3367AE2",
    x"3367744",
    x"33673A6",
    x"336700A",
    x"3366C6E",
    x"33668D4",
    x"336653A",
    x"33661A1",
    x"3365E09",
    x"3365A72",
    x"33656DC",
    x"3365346",
    x"3364FB2",
    x"3364C1F",
    x"336488C",
    x"33644FA",
    x"336416A",
    x"3363DDA",
    x"3363A4B",
    x"33636BD",
    x"336332F",
    x"3362FA3",
    x"3362C17",
    x"336288D",
    x"3362503",
    x"336217A",
    x"3361DF2",
    x"3361A6B",
    x"33616E5",
    x"3361360",
    x"3360FDC",
    x"3360C58",
    x"33608D5",
    x"3360554",
    x"33601D3",
    x"335FE53",
    x"335FAD4",
    x"335F755",
    x"335F3D8",
    x"335F05B",
    x"335ECE0",
    x"335E965",
    x"335E5EB",
    x"335E272",
    x"335DEFA",
    x"335DB82",
    x"335D80C",
    x"335D496",
    x"335D122",
    x"335CDAE",
    x"335CA3B",
    x"335C6C9",
    x"335C357",
    x"335BFE7",
    x"335BC78",
    x"335B909",
    x"335B59B",
    x"335B22E",
    x"335AEC2",
    x"335AB57",
    x"335A7EC",
    x"335A483",
    x"335A11A",
    x"3359DB2",
    x"3359A4B",
    x"33596E5",
    x"3359380",
    x"335901B",
    x"3358CB8",
    x"3358955",
    x"33585F3",
    x"3358292",
    x"3357F32",
    x"3357BD2",
    x"3357874",
    x"3357516",
    x"33571B9",
    x"3356E5D",
    x"3356B02",
    x"33567A8",
    x"335644E",
    x"33560F6",
    x"3355D9E",
    x"3355A47",
    x"33556F1",
    x"335539B",
    x"3355047",
    x"3354CF3",
    x"33549A0",
    x"335464E",
    x"33542FD",
    x"3353FAD",
    x"3353C5D",
    x"335390F",
    x"33535C1",
    x"3353274",
    x"3352F28",
    x"3352BDC",
    x"3352892",
    x"3352548",
    x"33521FF",
    x"3351EB7",
    x"3351B70",
    x"3351829",
    x"33514E4",
    x"335119F",
    x"3350E5B",
    x"3350B18",
    x"33507D5",
    x"3350494",
    x"3350153",
    x"334FE13",
    x"334FAD4",
    x"334F796",
    x"334F458",
    x"334F11B",
    x"334EDE0",
    x"334EAA4",
    x"334E76A",
    x"334E431",
    x"334E0F8",
    x"334DDC0",
    x"334DA89",
    x"334D753",
    x"334D41E",
    x"334D0E9",
    x"334CDB5",
    x"334CA82",
    x"334C750",
    x"334C41E",
    x"334C0EE",
    x"334BDBE",
    x"334BA8F",
    x"334B761",
    x"334B433",
    x"334B107",
    x"334ADDB",
    x"334AAB0",
    x"334A785",
    x"334A45C",
    x"334A133",
    x"3349E0B",
    x"3349AE4",
    x"33497BE",
    x"3349498",
    x"3349174",
    x"3348E50",
    x"3348B2C",
    x"334880A",
    x"33484E8",
    x"33481C8",
    x"3347EA7",
    x"3347B88",
    x"334786A",
    x"334754C",
    x"334722F",
    x"3346F13",
    x"3346BF8",
    x"33468DD",
    x"33465C3",
    x"33462AA",
    x"3345F92",
    x"3345C7A",
    x"3345964",
    x"334564E",
    x"3345338",
    x"3345024",
    x"3344D10",
    x"33449FD",
    x"33446EB",
    x"33443DA",
    x"33440C9",
    x"3343DBA",
    x"3343AAA",
    x"334379C",
    x"334348F",
    x"3343182",
    x"3342E76",
    x"3342B6B",
    x"3342860",
    x"3342557",
    x"334224E",
    x"3341F45",
    x"3341C3E",
    x"3341937",
    x"3341631",
    x"334132C",
    x"3341028",
    x"3340D24",
    x"3340A21",
    x"334071F",
    x"334041E",
    x"334011D",
    x"333FE1D",
    x"333FB1E",
    x"333F81F",
    x"333F522",
    x"333F225",
    x"333EF29",
    x"333EC2D",
    x"333E933",
    x"333E639",
    x"333E340",
    x"333E047",
    x"333DD4F",
    x"333DA58",
    x"333D762",
    x"333D46D",
    x"333D178",
    x"333CE84",
    x"333CB91",
    x"333C89E",
    x"333C5AC",
    x"333C2BB",
    x"333BFCB",
    x"333BCDB",
    x"333B9ED",
    x"333B6FF",
    x"333B411",
    x"333B124",
    x"333AE39",
    x"333AB4D",
    x"333A863",
    x"333A579",
    x"333A290",
    x"3339FA8",
    x"3339CC0",
    x"33399DA",
    x"33396F3",
    x"333940E",
    x"3339129",
    x"3338E45",
    x"3338B62",
    x"3338880",
    x"333859E",
    x"33382BD",
    x"3337FDD",
    x"3337CFD",
    x"3337A1E",
    x"3337740",
    x"3337463",
    x"3337186",
    x"3336EAA",
    x"3336BCE",
    x"33368F4",
    x"333661A",
    x"3336341",
    x"3336068",
    x"3335D91",
    x"3335ABA",
    x"33357E3",
    x"333550E",
    x"3335239",
    x"3334F65",
    x"3334C91",
    x"33349BE",
    x"33346EC",
    x"333441B",
    x"333414A",
    x"3333E7A",
    x"3333BAB",
    x"33338DC",
    x"333360E",
    x"3333341",
    x"3333075",
    x"3332DA9",
    x"3332ADE",
    x"3332814",
    x"333254A",
    x"3332281",
    x"3331FB9",
    x"3331CF1",
    x"3331A2A",
    x"3331764",
    x"333149E",
    x"33311DA",
    x"3330F16",
    x"3330C52",
    x"333098F",
    x"33306CD",
    x"333040C",
    x"333014B",
    x"332FE8B",
    x"332FBCC",
    x"332F90D",
    x"332F650",
    x"332F392",
    x"332F0D6",
    x"332EE1A",
    x"332EB5F",
    x"332E8A4",
    x"332E5EA",
    x"332E331",
    x"332E079",
    x"332DDC1",
    x"332DB0A",
    x"332D853",
    x"332D59E",
    x"332D2E9",
    x"332D034",
    x"332CD81",
    x"332CACE",
    x"332C81B",
    x"332C569",
    x"332C2B8",
    x"332C008",
    x"332BD58",
    x"332BAA9",
    x"332B7FB",
    x"332B54D",
    x"332B2A0",
    x"332AFF4",
    x"332AD48",
    x"332AA9D",
    x"332A7F3",
    x"332A54A",
    x"332A2A1",
    x"3329FF8",
    x"3329D51",
    x"3329AAA",
    x"3329803",
    x"332955E",
    x"33292B9",
    x"3329014",
    x"3328D70",
    x"3328ACD",
    x"332882B",
    x"3328589",
    x"33282E8",
    x"3328048",
    x"3327DA8",
    x"3327B09",
    x"332786B",
    x"33275CD",
    x"3327330",
    x"3327093",
    x"3326DF7",
    x"3326B5C",
    x"33268C2",
    x"3326628",
    x"332638F",
    x"33260F6",
    x"3325E5E",
    x"3325BC7",
    x"3325930",
    x"332569A",
    x"3325405",
    x"3325170",
    x"3324EDC",
    x"3324C49",
    x"33249B6",
    x"3324724",
    x"3324493",
    x"3324202",
    x"3323F72",
    x"3323CE2",
    x"3323A53",
    x"33237C5",
    x"3323537",
    x"33232AA",
    x"332301E",
    x"3322D92",
    x"3322B07",
    x"332287D",
    x"33225F3",
    x"332236A",
    x"33220E1",
    x"3321E59",
    x"3321BD2",
    x"332194B",
    x"33216C5",
    x"3321440",
    x"33211BB",
    x"3320F37",
    x"3320CB4",
    x"3320A31",
    x"33207AF",
    x"332052D",
    x"33202AC",
    x"332002C",
    x"331FDAC",
    x"331FB2D",
    x"331F8AE",
    x"331F630",
    x"331F3B3",
    x"331F137",
    x"331EEBB",
    x"331EC3F",
    x"331E9C4",
    x"331E74A",
    x"331E4D1",
    x"331E258",
    x"331DFE0",
    x"331DD68",
    x"331DAF1",
    x"331D87A",
    x"331D605",
    x"331D38F",
    x"331D11B",
    x"331CEA7",
    x"331CC34",
    x"331C9C1",
    x"331C74F",
    x"331C4DD",
    x"331C26C",
    x"331BFFC",
    x"331BD8C",
    x"331BB1D",
    x"331B8AF",
    x"331B641",
    x"331B3D4",
    x"331B167",
    x"331AEFB",
    x"331AC8F",
    x"331AA25",
    x"331A7BA",
    x"331A551",
    x"331A2E8",
    x"331A07F",
    x"3319E17",
    x"3319BB0",
    x"331994A",
    x"33196E4",
    x"331947E",
    x"3319219",
    x"3318FB5",
    x"3318D51",
    x"3318AEE",
    x"331888C",
    x"331862A",
    x"33183C9",
    x"3318168",
    x"3317F08",
    x"3317CA9",
    x"3317A4A",
    x"33177EC",
    x"331758E",
    x"3317331",
    x"33170D4",
    x"3316E78",
    x"3316C1D",
    x"33169C2",
    x"3316768",
    x"331650F",
    x"33162B6",
    x"331605D",
    x"3315E06",
    x"3315BAE",
    x"3315958",
    x"3315702",
    x"33154AC",
    x"3315257",
    x"3315003",
    x"3314DAF",
    x"3314B5C",
    x"331490A",
    x"33146B8",
    x"3314466",
    x"3314215",
    x"3313FC5",
    x"3313D76",
    x"3313B26",
    x"33138D8",
    x"331368A",
    x"331343D",
    x"33131F0",
    x"3312FA4",
    x"3312D58",
    x"3312B0D",
    x"33128C3",
    x"3312679",
    x"331242F",
    x"33121E7",
    x"3311F9E",
    x"3311D57",
    x"3311B10",
    x"33118C9",
    x"3311683",
    x"331143E",
    x"33111F9",
    x"3310FB5",
    x"3310D71",
    x"3310B2E",
    x"33108EC",
    x"33106AA",
    x"3310468",
    x"3310228",
    x"330FFE7",
    x"330FDA8",
    x"330FB69",
    x"330F92A",
    x"330F6EC",
    x"330F4AE",
    x"330F272",
    x"330F035",
    x"330EDF9",
    x"330EBBE",
    x"330E984",
    x"330E74A",
    x"330E510",
    x"330E2D7",
    x"330E09F",
    x"330DE67",
    x"330DC2F",
    x"330D9F9",
    x"330D7C2",
    x"330D58D",
    x"330D358",
    x"330D123",
    x"330CEEF",
    x"330CCBC",
    x"330CA89",
    x"330C856",
    x"330C624",
    x"330C3F3",
    x"330C1C2",
    x"330BF92",
    x"330BD63",
    x"330BB34",
    x"330B905",
    x"330B6D7",
    x"330B4AA",
    x"330B27D",
    x"330B050",
    x"330AE25",
    x"330ABF9",
    x"330A9CF",
    x"330A7A4",
    x"330A57B",
    x"330A352",
    x"330A129",
    x"3309F01",
    x"3309CDA",
    x"3309AB3",
    x"330988C",
    x"3309666",
    x"3309441",
    x"330921C",
    x"3308FF8",
    x"3308DD4",
    x"3308BB1",
    x"330898E",
    x"330876C",
    x"330854B",
    x"330832A",
    x"3308109",
    x"3307EE9",
    x"3307CCA",
    x"3307AAB",
    x"330788C",
    x"330766F",
    x"3307451",
    x"3307234",
    x"3307018",
    x"3306DFC",
    x"3306BE1",
    x"33069C6",
    x"33067AC",
    x"3306593",
    x"3306379",
    x"3306161",
    x"3305F49",
    x"3305D31",
    x"3305B1A",
    x"3305904",
    x"33056EE",
    x"33054D8",
    x"33052C3",
    x"33050AF",
    x"3304E9B",
    x"3304C87",
    x"3304A75",
    x"3304862",
    x"3304650",
    x"330443F",
    x"330422E",
    x"330401E",
    x"3303E0E",
    x"3303BFF",
    x"33039F0",
    x"33037E2",
    x"33035D4",
    x"33033C7",
    x"33031BA",
    x"3302FAE",
    x"3302DA3",
    x"3302B97",
    x"330298D",
    x"3302783",
    x"3302579",
    x"3302370",
    x"3302167",
    x"3301F5F",
    x"3301D58",
    x"3301B50",
    x"330194A",
    x"3301744",
    x"330153E",
    x"3301339",
    x"3301135",
    x"3300F31",
    x"3300D2D",
    x"3300B2A",
    x"3300927",
    x"3300725",
    x"3300524",
    x"3300323",
    x"3300122",
    x"32FFE45",
    x"32FFA46",
    x"32FF648",
    x"32FF24B",
    x"32FEE4F",
    x"32FEA54",
    x"32FE65A",
    x"32FE261",
    x"32FDE68",
    x"32FDA71",
    x"32FD67B",
    x"32FD286",
    x"32FCE92",
    x"32FCA9F",
    x"32FC6AD",
    x"32FC2BB",
    x"32FBECB",
    x"32FBADC",
    x"32FB6EE",
    x"32FB301",
    x"32FAF14",
    x"32FAB29",
    x"32FA73F",
    x"32FA355",
    x"32F9F6D",
    x"32F9B86",
    x"32F979F",
    x"32F93BA",
    x"32F8FD5",
    x"32F8BF2",
    x"32F880F",
    x"32F842E",
    x"32F804D",
    x"32F7C6E",
    x"32F788F",
    x"32F74B2",
    x"32F70D5",
    x"32F6CF9",
    x"32F691E",
    x"32F6545",
    x"32F616C",
    x"32F5D94",
    x"32F59BD",
    x"32F55E7",
    x"32F5212",
    x"32F4E3E",
    x"32F4A6B",
    x"32F4699",
    x"32F42C8",
    x"32F3EF7",
    x"32F3B28",
    x"32F375A",
    x"32F338C",
    x"32F2FC0",
    x"32F2BF5",
    x"32F282A",
    x"32F2460",
    x"32F2098",
    x"32F1CD0",
    x"32F1909",
    x"32F1544",
    x"32F117F",
    x"32F0DBB",
    x"32F09F8",
    x"32F0636",
    x"32F0275",
    x"32EFEB5",
    x"32EFAF5",
    x"32EF737",
    x"32EF37A",
    x"32EEFBD",
    x"32EEC02",
    x"32EE847",
    x"32EE48E",
    x"32EE0D5",
    x"32EDD1D",
    x"32ED967",
    x"32ED5B1",
    x"32ED1FC",
    x"32ECE48",
    x"32ECA95",
    x"32EC6E2",
    x"32EC331",
    x"32EBF81",
    x"32EBBD1",
    x"32EB823",
    x"32EB475",
    x"32EB0C9",
    x"32EAD1D",
    x"32EA972",
    x"32EA5C8",
    x"32EA21F",
    x"32E9E77",
    x"32E9AD0",
    x"32E972A",
    x"32E9384",
    x"32E8FE0",
    x"32E8C3C",
    x"32E889A",
    x"32E84F8",
    x"32E8157",
    x"32E7DB7",
    x"32E7A19",
    x"32E767A",
    x"32E72DD",
    x"32E6F41",
    x"32E6BA6",
    x"32E680B",
    x"32E6472",
    x"32E60D9",
    x"32E5D41",
    x"32E59AA",
    x"32E5614",
    x"32E527F",
    x"32E4EEB",
    x"32E4B58",
    x"32E47C5",
    x"32E4434",
    x"32E40A3",
    x"32E3D14",
    x"32E3985",
    x"32E35F7",
    x"32E326A",
    x"32E2EDE",
    x"32E2B52",
    x"32E27C8",
    x"32E243E",
    x"32E20B6",
    x"32E1D2E",
    x"32E19A7",
    x"32E1621",
    x"32E129C",
    x"32E0F18",
    x"32E0B95",
    x"32E0812",
    x"32E0491",
    x"32E0110",
    x"32DFD90",
    x"32DFA11",
    x"32DF693",
    x"32DF316",
    x"32DEF9A",
    x"32DEC1E",
    x"32DE8A3",
    x"32DE52A",
    x"32DE1B1",
    x"32DDE39",
    x"32DDAC2",
    x"32DD74C",
    x"32DD3D6",
    x"32DD062",
    x"32DCCEE",
    x"32DC97B",
    x"32DC609",
    x"32DC298",
    x"32DBF28",
    x"32DBBB9",
    x"32DB84A",
    x"32DB4DC",
    x"32DB170",
    x"32DAE04",
    x"32DAA99",
    x"32DA72E",
    x"32DA3C5",
    x"32DA05C",
    x"32D9CF5",
    x"32D998E",
    x"32D9628",
    x"32D92C3",
    x"32D8F5F",
    x"32D8BFB",
    x"32D8899",
    x"32D8537",
    x"32D81D6",
    x"32D7E76",
    x"32D7B17",
    x"32D77B8",
    x"32D745B",
    x"32D70FE",
    x"32D6DA2",
    x"32D6A47",
    x"32D66ED",
    x"32D6394",
    x"32D603C",
    x"32D5CE4",
    x"32D598D",
    x"32D5637",
    x"32D52E2",
    x"32D4F8E",
    x"32D4C3A",
    x"32D48E8",
    x"32D4596",
    x"32D4245",
    x"32D3EF5",
    x"32D3BA5",
    x"32D3857",
    x"32D3509",
    x"32D31BC",
    x"32D2E70",
    x"32D2B25",
    x"32D27DB",
    x"32D2491",
    x"32D2148",
    x"32D1E00",
    x"32D1AB9",
    x"32D1773",
    x"32D142E",
    x"32D10E9",
    x"32D0DA5",
    x"32D0A62",
    x"32D0720",
    x"32D03DF",
    x"32D009E",
    x"32CFD5E",
    x"32CFA1F",
    x"32CF6E1",
    x"32CF3A4",
    x"32CF067",
    x"32CED2C",
    x"32CE9F1",
    x"32CE6B7",
    x"32CE37D",
    x"32CE045",
    x"32CDD0D",
    x"32CD9D6",
    x"32CD6A0",
    x"32CD36B",
    x"32CD037",
    x"32CCD03",
    x"32CC9D0",
    x"32CC69E",
    x"32CC36D",
    x"32CC03C",
    x"32CBD0D",
    x"32CB9DE",
    x"32CB6B0",
    x"32CB383",
    x"32CB056",
    x"32CAD2A",
    x"32CAA00",
    x"32CA6D5",
    x"32CA3AC",
    x"32CA084",
    x"32C9D5C",
    x"32C9A35",
    x"32C970F",
    x"32C93E9",
    x"32C90C5",
    x"32C8DA1",
    x"32C8A7E",
    x"32C875C",
    x"32C843A",
    x"32C811A",
    x"32C7DFA",
    x"32C7ADB",
    x"32C77BC",
    x"32C749F",
    x"32C7182",
    x"32C6E66",
    x"32C6B4B",
    x"32C6830",
    x"32C6517",
    x"32C61FE",
    x"32C5EE6",
    x"32C5BCE",
    x"32C58B8",
    x"32C55A2",
    x"32C528D",
    x"32C4F79",
    x"32C4C65",
    x"32C4953",
    x"32C4641",
    x"32C432F",
    x"32C401F",
    x"32C3D0F",
    x"32C3A00",
    x"32C36F2",
    x"32C33E5",
    x"32C30D8",
    x"32C2DCD",
    x"32C2AC1",
    x"32C27B7",
    x"32C24AE",
    x"32C21A5",
    x"32C1E9D",
    x"32C1B96",
    x"32C188F",
    x"32C1589",
    x"32C1284",
    x"32C0F80",
    x"32C0C7C",
    x"32C097A",
    x"32C0678",
    x"32C0377",
    x"32C0076",
    x"32BFD76",
    x"32BFA77",
    x"32BF779",
    x"32BF47C",
    x"32BF17F",
    x"32BEE83",
    x"32BEB88",
    x"32BE88D",
    x"32BE593",
    x"32BE29A",
    x"32BDFA2",
    x"32BDCAA",
    x"32BD9B4",
    x"32BD6BE",
    x"32BD3C8",
    x"32BD0D4",
    x"32BCDE0",
    x"32BCAED",
    x"32BC7FA",
    x"32BC509",
    x"32BC218",
    x"32BBF28",
    x"32BBC38",
    x"32BB94A",
    x"32BB65C",
    x"32BB36E",
    x"32BB082",
    x"32BAD96",
    x"32BAAAB",
    x"32BA7C1",
    x"32BA4D7",
    x"32BA1EE",
    x"32B9F06",
    x"32B9C1F",
    x"32B9938",
    x"32B9652",
    x"32B936D",
    x"32B9089",
    x"32B8DA5",
    x"32B8AC2",
    x"32B87DF",
    x"32B84FE",
    x"32B821D",
    x"32B7F3D",
    x"32B7C5D",
    x"32B797F",
    x"32B76A1",
    x"32B73C3",
    x"32B70E7",
    x"32B6E0B",
    x"32B6B30",
    x"32B6855",
    x"32B657B",
    x"32B62A2",
    x"32B5FCA",
    x"32B5CF3",
    x"32B5A1C",
    x"32B5746",
    x"32B5470",
    x"32B519B",
    x"32B4EC7",
    x"32B4BF4",
    x"32B4921",
    x"32B464F",
    x"32B437E",
    x"32B40AE",
    x"32B3DDE",
    x"32B3B0F",
    x"32B3840",
    x"32B3573",
    x"32B32A6",
    x"32B2FD9",
    x"32B2D0E",
    x"32B2A43",
    x"32B2778",
    x"32B24AF",
    x"32B21E6",
    x"32B1F1E",
    x"32B1C57",
    x"32B1990",
    x"32B16CA",
    x"32B1404",
    x"32B1140",
    x"32B0E7C",
    x"32B0BB9",
    x"32B08F6",
    x"32B0634",
    x"32B0373",
    x"32B00B2",
    x"32AFDF2",
    x"32AFB33",
    x"32AF875",
    x"32AF5B7",
    x"32AF2FA",
    x"32AF03E",
    x"32AED82",
    x"32AEAC7",
    x"32AE80D",
    x"32AE553",
    x"32AE29A",
    x"32ADFE2",
    x"32ADD2A",
    x"32ADA73",
    x"32AD7BD",
    x"32AD507",
    x"32AD252",
    x"32ACF9E",
    x"32ACCEA",
    x"32ACA37",
    x"32AC785",
    x"32AC4D4",
    x"32AC223",
    x"32ABF73",
    x"32ABCC3",
    x"32ABA14",
    x"32AB766",
    x"32AB4B9",
    x"32AB20C",
    x"32AAF60",
    x"32AACB4",
    x"32AAA09",
    x"32AA75F",
    x"32AA4B5",
    x"32AA20D",
    x"32A9F64",
    x"32A9CBD",
    x"32A9A16",
    x"32A9770",
    x"32A94CA",
    x"32A9226",
    x"32A8F81",
    x"32A8CDE",
    x"32A8A3B",
    x"32A8799",
    x"32A84F7",
    x"32A8256",
    x"32A7FB6",
    x"32A7D16",
    x"32A7A77",
    x"32A77D9",
    x"32A753B",
    x"32A729E",
    x"32A7002",
    x"32A6D66",
    x"32A6ACB",
    x"32A6831",
    x"32A6597",
    x"32A62FE",
    x"32A6066",
    x"32A5DCE",
    x"32A5B37",
    x"32A58A0",
    x"32A560B",
    x"32A5375",
    x"32A50E1",
    x"32A4E4D",
    x"32A4BBA",
    x"32A4927",
    x"32A4695",
    x"32A4404",
    x"32A4173",
    x"32A3EE3",
    x"32A3C54",
    x"32A39C5",
    x"32A3737",
    x"32A34A9",
    x"32A321C",
    x"32A2F90",
    x"32A2D05",
    x"32A2A7A",
    x"32A27EF",
    x"32A2566",
    x"32A22DD",
    x"32A2054",
    x"32A1DCD",
    x"32A1B45",
    x"32A18BF",
    x"32A1639",
    x"32A13B4",
    x"32A112F",
    x"32A0EAB",
    x"32A0C28",
    x"32A09A5",
    x"32A0723",
    x"32A04A2",
    x"32A0221",
    x"329FFA1",
    x"329FD21",
    x"329FAA2",
    x"329F824",
    x"329F5A6",
    x"329F329",
    x"329F0AC",
    x"329EE30",
    x"329EBB5",
    x"329E93B",
    x"329E6C1",
    x"329E447",
    x"329E1CE",
    x"329DF56",
    x"329DCDF",
    x"329DA68",
    x"329D7F2",
    x"329D57C",
    x"329D307",
    x"329D092",
    x"329CE1F",
    x"329CBAB",
    x"329C939",
    x"329C6C7",
    x"329C455",
    x"329C1E5",
    x"329BF74",
    x"329BD05",
    x"329BA96",
    x"329B828",
    x"329B5BA",
    x"329B34D",
    x"329B0E0",
    x"329AE74",
    x"329AC09",
    x"329A99E",
    x"329A734",
    x"329A4CB",
    x"329A262",
    x"3299FF9",
    x"3299D92",
    x"3299B2B",
    x"32998C4",
    x"329965E",
    x"32993F9",
    x"3299194",
    x"3298F30",
    x"3298CCD",
    x"3298A6A",
    x"3298807",
    x"32985A6",
    x"3298345",
    x"32980E4",
    x"3297E84",
    x"3297C25",
    x"32979C6",
    x"3297768",
    x"329750A",
    x"32972AD",
    x"3297051",
    x"3296DF5",
    x"3296B9A",
    x"329693F",
    x"32966E5",
    x"329648C",
    x"3296233",
    x"3295FDB",
    x"3295D83",
    x"3295B2C",
    x"32958D6",
    x"3295680",
    x"329542A",
    x"32951D6",
    x"3294F81",
    x"3294D2E",
    x"3294ADB",
    x"3294888",
    x"3294637",
    x"32943E5",
    x"3294195",
    x"3293F45",
    x"3293CF5",
    x"3293AA6",
    x"3293858",
    x"329360A",
    x"32933BD",
    x"3293170",
    x"3292F24",
    x"3292CD8",
    x"3292A8E",
    x"3292843",
    x"32925F9",
    x"32923B0",
    x"3292168",
    x"3291F20",
    x"3291CD8",
    x"3291A91",
    x"329184B",
    x"3291605",
    x"32913C0",
    x"329117B",
    x"3290F37",
    x"3290CF3",
    x"3290AB1",
    x"329086E",
    x"329062C",
    x"32903EB",
    x"32901AA",
    x"328FF6A",
    x"328FD2B",
    x"328FAEC",
    x"328F8AD",
    x"328F66F",
    x"328F432",
    x"328F1F5",
    x"328EFB9",
    x"328ED7D",
    x"328EB42",
    x"328E908",
    x"328E6CE",
    x"328E494",
    x"328E25B",
    x"328E023",
    x"328DDEB",
    x"328DBB4",
    x"328D97D",
    x"328D747",
    x"328D512",
    x"328D2DD",
    x"328D0A8",
    x"328CE75",
    x"328CC41",
    x"328CA0E",
    x"328C7DC",
    x"328C5AA",
    x"328C379",
    x"328C149",
    x"328BF19",
    x"328BCE9",
    x"328BABA",
    x"328B88C",
    x"328B65E",
    x"328B431",
    x"328B204",
    x"328AFD8",
    x"328ADAC",
    x"328AB81",
    x"328A956",
    x"328A72C",
    x"328A503",
    x"328A2DA",
    x"328A0B1",
    x"3289E89",
    x"3289C62",
    x"3289A3B",
    x"3289815",
    x"32895EF",
    x"32893CA",
    x"32891A5",
    x"3288F81",
    x"3288D5D",
    x"3288B3A",
    x"3288918",
    x"32886F6",
    x"32884D4",
    x"32882B3",
    x"3288093",
    x"3287E73",
    x"3287C54",
    x"3287A35",
    x"3287817",
    x"32875F9",
    x"32873DC",
    x"32871BF",
    x"3286FA3",
    x"3286D87",
    x"3286B6C",
    x"3286951",
    x"3286737",
    x"328651E",
    x"3286305",
    x"32860EC",
    x"3285ED4",
    x"3285CBD",
    x"3285AA6",
    x"3285890",
    x"328567A",
    x"3285464",
    x"328524F",
    x"328503B",
    x"3284E27",
    x"3284C14",
    x"3284A01",
    x"32847EF",
    x"32845DD",
    x"32843CC",
    x"32841BB",
    x"3283FAB",
    x"3283D9C",
    x"3283B8C",
    x"328397E",
    x"3283770",
    x"3283562",
    x"3283355",
    x"3283148",
    x"3282F3C",
    x"3282D31",
    x"3282B26",
    x"328291B",
    x"3282711",
    x"3282508",
    x"32822FF",
    x"32820F6",
    x"3281EEE",
    x"3281CE7",
    x"3281AE0",
    x"32818D9",
    x"32816D3",
    x"32814CE",
    x"32812C9",
    x"32810C4",
    x"3280EC1",
    x"3280CBD",
    x"3280ABA",
    x"32808B8",
    x"32806B6",
    x"32804B4",
    x"32802B3",
    x"32800B3",
    x"327FD67",
    x"327F968",
    x"327F56A",
    x"327F16D",
    x"327ED71",
    x"327E976",
    x"327E57D",
    x"327E184",
    x"327DD8C",
    x"327D995",
    x"327D59F",
    x"327D1AA",
    x"327CDB6",
    x"327C9C3",
    x"327C5D1",
    x"327C1E0",
    x"327BDF0",
    x"327BA01",
    x"327B613",
    x"327B226",
    x"327AE3A",
    x"327AA4F",
    x"327A665",
    x"327A27C",
    x"3279E94",
    x"3279AAD",
    x"32796C7",
    x"32792E1",
    x"3278EFD",
    x"3278B1A",
    x"3278738",
    x"3278356",
    x"3277F76",
    x"3277B96",
    x"32777B8",
    x"32773DB",
    x"3276FFE",
    x"3276C23",
    x"3276848",
    x"327646E",
    x"3276096",
    x"3275CBE",
    x"32758E7",
    x"3275512",
    x"327513D",
    x"3274D69",
    x"3274996",
    x"32745C4",
    x"32741F3",
    x"3273E23",
    x"3273A54",
    x"3273686",
    x"32732B9",
    x"3272EED",
    x"3272B22",
    x"3272757",
    x"327238E",
    x"3271FC5",
    x"3271BFE",
    x"3271837",
    x"3271472",
    x"32710AD",
    x"3270CEA",
    x"3270927",
    x"3270565",
    x"32701A4",
    x"326FDE4",
    x"326FA25",
    x"326F667",
    x"326F2AA",
    x"326EEEE",
    x"326EB32",
    x"326E778",
    x"326E3BF",
    x"326E006",
    x"326DC4F",
    x"326D898",
    x"326D4E2",
    x"326D12E",
    x"326CD7A",
    x"326C9C7",
    x"326C615",
    x"326C264",
    x"326BEB4",
    x"326BB05",
    x"326B756",
    x"326B3A9",
    x"326AFFC",
    x"326AC51",
    x"326A8A6",
    x"326A4FD",
    x"326A154",
    x"3269DAC",
    x"3269A05",
    x"326965F",
    x"32692BA",
    x"3268F15",
    x"3268B72",
    x"32687D0",
    x"326842E",
    x"326808E",
    x"3267CEE",
    x"326794F",
    x"32675B1",
    x"3267214",
    x"3266E78",
    x"3266ADD",
    x"3266743",
    x"32663AA",
    x"3266011",
    x"3265C79",
    x"32658E3",
    x"326554D",
    x"32651B8",
    x"3264E24",
    x"3264A91",
    x"32646FF",
    x"326436E",
    x"3263FDD",
    x"3263C4E",
    x"32638BF",
    x"3263531",
    x"32631A4",
    x"3262E18",
    x"3262A8D",
    x"3262703",
    x"326237A",
    x"3261FF1",
    x"3261C6A",
    x"32618E3",
    x"326155D",
    x"32611D9",
    x"3260E55",
    x"3260AD1",
    x"326074F",
    x"32603CE",
    x"326004D",
    x"325FCCE",
    x"325F94F",
    x"325F5D1",
    x"325F254",
    x"325EED8",
    x"325EB5C",
    x"325E7E2",
    x"325E469",
    x"325E0F0",
    x"325DD78",
    x"325DA01",
    x"325D68B",
    x"325D316",
    x"325CFA2",
    x"325CC2E",
    x"325C8BB",
    x"325C54A",
    x"325C1D9",
    x"325BE69",
    x"325BAFA",
    x"325B78B",
    x"325B41E",
    x"325B0B1",
    x"325AD45",
    x"325A9DB",
    x"325A671",
    x"325A307",
    x"3259F9F",
    x"3259C38",
    x"32598D1",
    x"325956B",
    x"3259206",
    x"3258EA2",
    x"3258B3F",
    x"32587DC",
    x"325847B",
    x"325811A",
    x"3257DBA",
    x"3257A5B",
    x"32576FD",
    x"32573A0",
    x"3257043",
    x"3256CE8",
    x"325698D",
    x"3256633",
    x"32562DA",
    x"3255F82",
    x"3255C2A",
    x"32558D3",
    x"325557E",
    x"3255229",
    x"3254ED5",
    x"3254B81",
    x"325482F",
    x"32544DD",
    x"325418C",
    x"3253E3C",
    x"3253AED",
    x"325379F",
    x"3253451",
    x"3253105",
    x"3252DB9",
    x"3252A6E",
    x"3252724",
    x"32523DA",
    x"3252092",
    x"3251D4A",
    x"3251A03",
    x"32516BD",
    x"3251378",
    x"3251033",
    x"3250CF0",
    x"32509AD",
    x"325066B",
    x"325032A",
    x"324FFE9",
    x"324FCAA",
    x"324F96B",
    x"324F62D",
    x"324F2F0",
    x"324EFB4",
    x"324EC78",
    x"324E93D",
    x"324E603",
    x"324E2CA",
    x"324DF92",
    x"324DC5A",
    x"324D924",
    x"324D5EE",
    x"324D2B9",
    x"324CF85",
    x"324CC51",
    x"324C91E",
    x"324C5ED",
    x"324C2BB",
    x"324BF8B",
    x"324BC5C",
    x"324B92D",
    x"324B5FF",
    x"324B2D2",
    x"324AFA6",
    x"324AC7A",
    x"324A94F",
    x"324A625",
    x"324A2FC",
    x"3249FD4",
    x"3249CAC",
    x"3249986",
    x"3249660",
    x"324933A",
    x"3249016",
    x"3248CF2",
    x"32489D0",
    x"32486AE",
    x"324838C",
    x"324806C",
    x"3247D4C",
    x"3247A2D",
    x"324770F",
    x"32473F2",
    x"32470D5",
    x"3246DB9",
    x"3246A9E",
    x"3246784",
    x"324646A",
    x"3246152",
    x"3245E3A",
    x"3245B23",
    x"324580C",
    x"32454F6",
    x"32451E2",
    x"3244ECE",
    x"3244BBA",
    x"32448A8",
    x"3244596",
    x"3244285",
    x"3243F75",
    x"3243C65",
    x"3243956",
    x"3243648",
    x"324333B",
    x"324302F",
    x"3242D23",
    x"3242A18",
    x"324270E",
    x"3242405",
    x"32420FC",
    x"3241DF4",
    x"3241AED",
    x"32417E7",
    x"32414E1",
    x"32411DC",
    x"3240ED8",
    x"3240BD5",
    x"32408D2",
    x"32405D1",
    x"32402CF",
    x"323FFCF",
    x"323FCD0",
    x"323F9D1",
    x"323F6D3",
    x"323F3D5",
    x"323F0D9",
    x"323EDDD",
    x"323EAE2",
    x"323E7E7",
    x"323E4EE",
    x"323E1F5",
    x"323DEFD",
    x"323DC05",
    x"323D90F",
    x"323D619",
    x"323D324",
    x"323D02F",
    x"323CD3C",
    x"323CA49",
    x"323C757",
    x"323C465",
    x"323C174",
    x"323BE84",
    x"323BB95",
    x"323B8A7",
    x"323B5B9",
    x"323B2CC",
    x"323AFDF",
    x"323ACF4",
    x"323AA09",
    x"323A71F",
    x"323A435",
    x"323A14D",
    x"3239E65",
    x"3239B7D",
    x"3239897",
    x"32395B1",
    x"32392CC",
    x"3238FE8",
    x"3238D04",
    x"3238A21",
    x"323873F",
    x"323845E",
    x"323817D",
    x"3237E9D",
    x"3237BBE",
    x"32378DF",
    x"3237601",
    x"3237324",
    x"3237048",
    x"3236D6C",
    x"3236A91",
    x"32367B7",
    x"32364DD",
    x"3236204",
    x"3235F2C",
    x"3235C55",
    x"323597E",
    x"32356A8",
    x"32353D3",
    x"32350FE",
    x"3234E2A",
    x"3234B57",
    x"3234884",
    x"32345B3",
    x"32342E1",
    x"3234011",
    x"3233D41",
    x"3233A72",
    x"32337A4",
    x"32334D7",
    x"323320A",
    x"3232F3E",
    x"3232C72",
    x"32329A7",
    x"32326DD",
    x"3232414",
    x"323214B",
    x"3231E83",
    x"3231BBC",
    x"32318F5",
    x"3231630",
    x"323136A",
    x"32310A6",
    x"3230DE2",
    x"3230B1F",
    x"323085C",
    x"323059B",
    x"32302DA",
    x"3230019",
    x"322FD5A",
    x"322FA9B",
    x"322F7DC",
    x"322F51F",
    x"322F262",
    x"322EFA6",
    x"322ECEA",
    x"322EA2F",
    x"322E775",
    x"322E4BB",
    x"322E202",
    x"322DF4A",
    x"322DC93",
    x"322D9DC",
    x"322D726",
    x"322D470",
    x"322D1BC",
    x"322CF08",
    x"322CC54",
    x"322C9A1",
    x"322C6EF",
    x"322C43E",
    x"322C18D",
    x"322BEDD",
    x"322BC2E",
    x"322B97F",
    x"322B6D1",
    x"322B424",
    x"322B177",
    x"322AECB",
    x"322AC20",
    x"322A975",
    x"322A6CB",
    x"322A421",
    x"322A179",
    x"3229ED1",
    x"3229C29",
    x"3229983",
    x"32296DD",
    x"3229437",
    x"3229193",
    x"3228EEE",
    x"3228C4B",
    x"32289A8",
    x"3228706",
    x"3228465",
    x"32281C4",
    x"3227F24",
    x"3227C84",
    x"32279E6",
    x"3227747",
    x"32274AA",
    x"322720D",
    x"3226F71",
    x"3226CD5",
    x"3226A3B",
    x"32267A0",
    x"3226507",
    x"322626E",
    x"3225FD6",
    x"3225D3E",
    x"3225AA7",
    x"3225811",
    x"322557B",
    x"32252E6",
    x"3225051",
    x"3224DBE",
    x"3224B2B",
    x"3224898",
    x"3224606",
    x"3224375",
    x"32240E5",
    x"3223E55",
    x"3223BC5",
    x"3223937",
    x"32236A9",
    x"322341B",
    x"322318F",
    x"3222F03",
    x"3222C77",
    x"32229EC",
    x"3222762",
    x"32224D9",
    x"3222250",
    x"3221FC8",
    x"3221D40",
    x"3221AB9",
    x"3221833",
    x"32215AD",
    x"3221328",
    x"32210A3",
    x"3220E1F",
    x"3220B9C",
    x"322091A",
    x"3220698",
    x"3220416",
    x"3220196",
    x"321FF15",
    x"321FC96",
    x"321FA17",
    x"321F799",
    x"321F51B",
    x"321F29E",
    x"321F022",
    x"321EDA6",
    x"321EB2B",
    x"321E8B1",
    x"321E637",
    x"321E3BE",
    x"321E145",
    x"321DECD",
    x"321DC56",
    x"321D9DF",
    x"321D769",
    x"321D4F3",
    x"321D27E",
    x"321D00A",
    x"321CD96",
    x"321CB23",
    x"321C8B1",
    x"321C63F",
    x"321C3CE",
    x"321C15D",
    x"321BEED",
    x"321BC7D",
    x"321BA0F",
    x"321B7A0",
    x"321B533",
    x"321B2C6",
    x"321B059",
    x"321ADEE",
    x"321AB82",
    x"321A918",
    x"321A6AE",
    x"321A445",
    x"321A1DC",
    x"3219F74",
    x"3219D0C",
    x"3219AA5",
    x"321983F",
    x"32195D9",
    x"3219374",
    x"321910F",
    x"3218EAB",
    x"3218C48",
    x"32189E5",
    x"3218783",
    x"3218521",
    x"32182C0",
    x"3218060",
    x"3217E00",
    x"3217BA1",
    x"3217942",
    x"32176E4",
    x"3217487",
    x"321722A",
    x"3216FCE",
    x"3216D72",
    x"3216B17",
    x"32168BD",
    x"3216663",
    x"3216409",
    x"32161B1",
    x"3215F59",
    x"3215D01",
    x"3215AAA",
    x"3215854",
    x"32155FE",
    x"32153A9",
    x"3215154",
    x"3214F00",
    x"3214CAD",
    x"3214A5A",
    x"3214807",
    x"32145B6",
    x"3214365",
    x"3214114",
    x"3213EC4",
    x"3213C75",
    x"3213A26",
    x"32137D8",
    x"321358A",
    x"321333D",
    x"32130F0",
    x"3212EA4",
    x"3212C59",
    x"3212A0E",
    x"32127C4",
    x"321257A",
    x"3212331",
    x"32120E9",
    x"3211EA1",
    x"3211C59",
    x"3211A13",
    x"32117CC",
    x"3211587",
    x"3211342",
    x"32110FD",
    x"3210EB9",
    x"3210C76",
    x"3210A33",
    x"32107F1",
    x"32105AF",
    x"321036E",
    x"321012D",
    x"320FEED",
    x"320FCAE",
    x"320FA6F",
    x"320F830",
    x"320F5F3",
    x"320F3B5",
    x"320F179",
    x"320EF3D",
    x"320ED01",
    x"320EAC6",
    x"320E88C",
    x"320E652",
    x"320E419",
    x"320E1E0",
    x"320DFA8",
    x"320DD70",
    x"320DB39",
    x"320D902",
    x"320D6CC",
    x"320D497",
    x"320D262",
    x"320D02E",
    x"320CDFA",
    x"320CBC7",
    x"320C994",
    x"320C762",
    x"320C530",
    x"320C2FF",
    x"320C0CF",
    x"320BE9F",
    x"320BC70",
    x"320BA41",
    x"320B813",
    x"320B5E5",
    x"320B3B8",
    x"320B18B",
    x"320AF5F",
    x"320AD33",
    x"320AB08",
    x"320A8DE",
    x"320A6B4",
    x"320A48A",
    x"320A262",
    x"320A039",
    x"3209E11",
    x"3209BEA",
    x"32099C3",
    x"320979D",
    x"3209578",
    x"3209353",
    x"320912E",
    x"3208F0A",
    x"3208CE6",
    x"3208AC4",
    x"32088A1",
    x"320867F",
    x"320845E",
    x"320823D",
    x"320801D",
    x"3207DFD",
    x"3207BDE",
    x"32079BF",
    x"32077A1",
    x"3207583",
    x"3207366",
    x"3207149",
    x"3206F2D",
    x"3206D12",
    x"3206AF7",
    x"32068DC",
    x"32066C2",
    x"32064A9",
    x"3206290",
    x"3206078",
    x"3205E60",
    x"3205C49",
    x"3205A32",
    x"320581B",
    x"3205606",
    x"32053F0",
    x"32051DC",
    x"3204FC8",
    x"3204DB4",
    x"3204BA1",
    x"320498E",
    x"320477C",
    x"320456A",
    x"3204359",
    x"3204149",
    x"3203F39",
    x"3203D29",
    x"3203B1A",
    x"320390B",
    x"32036FD",
    x"32034F0",
    x"32032E3",
    x"32030D7",
    x"3202ECB",
    x"3202CBF",
    x"3202AB4",
    x"32028AA",
    x"32026A0",
    x"3202496",
    x"320228E",
    x"3202085",
    x"3201E7D",
    x"3201C76",
    x"3201A6F",
    x"3201869",
    x"3201663",
    x"320145E",
    x"3201259",
    x"3201054",
    x"3200E51",
    x"3200C4D",
    x"3200A4A",
    x"3200848",
    x"3200646",
    x"3200445",
    x"3200244",
    x"3200044",
    x"31FFC88",
    x"31FF88A",
    x"31FF48C",
    x"31FF08F",
    x"31FEC94",
    x"31FE899",
    x"31FE4A0",
    x"31FE0A7",
    x"31FDCAF",
    x"31FD8B8",
    x"31FD4C3",
    x"31FD0CE",
    x"31FCCDA",
    x"31FC8E8",
    x"31FC4F6",
    x"31FC105",
    x"31FBD15",
    x"31FB927",
    x"31FB539",
    x"31FB14C",
    x"31FAD60",
    x"31FA975",
    x"31FA58B",
    x"31FA1A3",
    x"31F9DBB",
    x"31F99D4",
    x"31F95EE",
    x"31F9209",
    x"31F8E25",
    x"31F8A42",
    x"31F8660",
    x"31F827E",
    x"31F7E9E",
    x"31F7ABF",
    x"31F76E1",
    x"31F7304",
    x"31F6F27",
    x"31F6B4C",
    x"31F6772",
    x"31F6398",
    x"31F5FC0",
    x"31F5BE9",
    x"31F5812",
    x"31F543D",
    x"31F5068",
    x"31F4C94",
    x"31F48C2",
    x"31F44F0",
    x"31F411F",
    x"31F3D4F",
    x"31F3981",
    x"31F35B3",
    x"31F31E6",
    x"31F2E1A",
    x"31F2A4F",
    x"31F2685",
    x"31F22BB",
    x"31F1EF3",
    x"31F1B2C",
    x"31F1766",
    x"31F13A0",
    x"31F0FDC",
    x"31F0C18",
    x"31F0856",
    x"31F0494",
    x"31F00D3",
    x"31EFD14",
    x"31EF955",
    x"31EF597",
    x"31EF1DA",
    x"31EEE1E",
    x"31EEA63",
    x"31EE6A9",
    x"31EE2F0",
    x"31EDF37",
    x"31EDB80",
    x"31ED7CA",
    x"31ED414",
    x"31ED060",
    x"31ECCAC",
    x"31EC8F9",
    x"31EC548",
    x"31EC197",
    x"31EBDE7",
    x"31EBA38",
    x"31EB68A",
    x"31EB2DC",
    x"31EAF30",
    x"31EAB85",
    x"31EA7DA",
    x"31EA431",
    x"31EA088",
    x"31E9CE1",
    x"31E993A",
    x"31E9594",
    x"31E91EF",
    x"31E8E4B",
    x"31E8AA8",
    x"31E8706",
    x"31E8364",
    x"31E7FC4",
    x"31E7C25",
    x"31E7886",
    x"31E74E8",
    x"31E714C",
    x"31E6DB0",
    x"31E6A15",
    x"31E667B",
    x"31E62E1",
    x"31E5F49",
    x"31E5BB2",
    x"31E581B",
    x"31E5486",
    x"31E50F1",
    x"31E4D5D",
    x"31E49CA",
    x"31E4638",
    x"31E42A7",
    x"31E3F17",
    x"31E3B88",
    x"31E37F9",
    x"31E346C",
    x"31E30DF",
    x"31E2D53",
    x"31E29C8",
    x"31E263E",
    x"31E22B5",
    x"31E1F2D",
    x"31E1BA6",
    x"31E181F",
    x"31E149A",
    x"31E1115",
    x"31E0D91",
    x"31E0A0E",
    x"31E068C",
    x"31E030B",
    x"31DFF8B",
    x"31DFC0B",
    x"31DF88C",
    x"31DF50F",
    x"31DF192",
    x"31DEE16",
    x"31DEA9B",
    x"31DE721",
    x"31DE3A7",
    x"31DE02F",
    x"31DDCB7",
    x"31DD941",
    x"31DD5CB",
    x"31DD256",
    x"31DCEE1",
    x"31DCB6E",
    x"31DC7FC",
    x"31DC48A",
    x"31DC119",
    x"31DBDAA",
    x"31DBA3B",
    x"31DB6CD",
    x"31DB35F",
    x"31DAFF3",
    x"31DAC87",
    x"31DA91D",
    x"31DA5B3",
    x"31DA24A",
    x"31D9EE2",
    x"31D9B7A",
    x"31D9814",
    x"31D94AE",
    x"31D9149",
    x"31D8DE6",
    x"31D8A83",
    x"31D8720",
    x"31D83BF",
    x"31D805E",
    x"31D7CFF",
    x"31D79A0",
    x"31D7642",
    x"31D72E5",
    x"31D6F89",
    x"31D6C2D",
    x"31D68D2",
    x"31D6579",
    x"31D6220",
    x"31D5EC8",
    x"31D5B70",
    x"31D581A",
    x"31D54C4",
    x"31D516F",
    x"31D4E1C",
    x"31D4AC8",
    x"31D4776",
    x"31D4425",
    x"31D40D4",
    x"31D3D84",
    x"31D3A35",
    x"31D36E7",
    x"31D339A",
    x"31D304D",
    x"31D2D02",
    x"31D29B7",
    x"31D266D",
    x"31D2324",
    x"31D1FDB",
    x"31D1C94",
    x"31D194D",
    x"31D1607",
    x"31D12C2",
    x"31D0F7E",
    x"31D0C3A",
    x"31D08F8",
    x"31D05B6",
    x"31D0275",
    x"31CFF35",
    x"31CFBF5",
    x"31CF8B7",
    x"31CF579",
    x"31CF23C",
    x"31CEF00",
    x"31CEBC4",
    x"31CE88A",
    x"31CE550",
    x"31CE217",
    x"31CDEDF",
    x"31CDBA8",
    x"31CD871",
    x"31CD53B",
    x"31CD207",
    x"31CCED2",
    x"31CCB9F",
    x"31CC86D",
    x"31CC53B",
    x"31CC20A",
    x"31CBEDA",
    x"31CBBAB",
    x"31CB87C",
    x"31CB54E",
    x"31CB221",
    x"31CAEF5",
    x"31CABCA",
    x"31CA89F",
    x"31CA576",
    x"31CA24D",
    x"31C9F24",
    x"31C9BFD",
    x"31C98D6",
    x"31C95B1",
    x"31C928C",
    x"31C8F67",
    x"31C8C44",
    x"31C8921",
    x"31C85FF",
    x"31C82DE",
    x"31C7FBE",
    x"31C7C9E",
    x"31C7980",
    x"31C7662",
    x"31C7344",
    x"31C7028",
    x"31C6D0C",
    x"31C69F1",
    x"31C66D7",
    x"31C63BE",
    x"31C60A5",
    x"31C5D8E",
    x"31C5A77",
    x"31C5760",
    x"31C544B",
    x"31C5136",
    x"31C4E22",
    x"31C4B0F",
    x"31C47FD",
    x"31C44EB",
    x"31C41DA",
    x"31C3ECA",
    x"31C3BBB",
    x"31C38AC",
    x"31C359F",
    x"31C3292",
    x"31C2F85",
    x"31C2C7A",
    x"31C296F",
    x"31C2665",
    x"31C235C",
    x"31C2053",
    x"31C1D4C",
    x"31C1A45",
    x"31C173F",
    x"31C1439",
    x"31C1135",
    x"31C0E31",
    x"31C0B2D",
    x"31C082B",
    x"31C0529",
    x"31C0228",
    x"31BFF28",
    x"31BFC29",
    x"31BF92A",
    x"31BF62C",
    x"31BF32F",
    x"31BF033",
    x"31BED37",
    x"31BEA3C",
    x"31BE742",
    x"31BE448",
    x"31BE150",
    x"31BDE58",
    x"31BDB61",
    x"31BD86A",
    x"31BD574",
    x"31BD27F",
    x"31BCF8B",
    x"31BCC98",
    x"31BC9A5",
    x"31BC6B3",
    x"31BC3C1",
    x"31BC0D1",
    x"31BBDE1",
    x"31BBAF2",
    x"31BB804",
    x"31BB516",
    x"31BB229",
    x"31BAF3D",
    x"31BAC51",
    x"31BA967",
    x"31BA67D",
    x"31BA393",
    x"31BA0AB",
    x"31B9DC3",
    x"31B9ADC",
    x"31B97F6",
    x"31B9510",
    x"31B922B",
    x"31B8F47",
    x"31B8C64",
    x"31B8981",
    x"31B869F",
    x"31B83BD",
    x"31B80DD",
    x"31B7DFD",
    x"31B7B1E",
    x"31B783F",
    x"31B7562",
    x"31B7285",
    x"31B6FA9",
    x"31B6CCD",
    x"31B69F2",
    x"31B6718",
    x"31B643F",
    x"31B6166",
    x"31B5E8E",
    x"31B5BB7",
    x"31B58E0",
    x"31B560A",
    x"31B5335",
    x"31B5061",
    x"31B4D8D",
    x"31B4ABA",
    x"31B47E7",
    x"31B4516",
    x"31B4245",
    x"31B3F75",
    x"31B3CA5",
    x"31B39D6",
    x"31B3708",
    x"31B343B",
    x"31B316E",
    x"31B2EA2",
    x"31B2BD7",
    x"31B290C",
    x"31B2642",
    x"31B2379",
    x"31B20B1",
    x"31B1DE9",
    x"31B1B22",
    x"31B185B",
    x"31B1595",
    x"31B12D0",
    x"31B100C",
    x"31B0D48",
    x"31B0A85",
    x"31B07C3",
    x"31B0501",
    x"31B0241",
    x"31AFF80",
    x"31AFCC1",
    x"31AFA02",
    x"31AF744",
    x"31AF486",
    x"31AF1CA",
    x"31AEF0D",
    x"31AEC52",
    x"31AE997",
    x"31AE6DD",
    x"31AE424",
    x"31AE16B",
    x"31ADEB3",
    x"31ADBFC",
    x"31AD945",
    x"31AD68F",
    x"31AD3DA",
    x"31AD125",
    x"31ACE71",
    x"31ACBBE",
    x"31AC90B",
    x"31AC65A",
    x"31AC3A8",
    x"31AC0F8",
    x"31ABE48",
    x"31ABB99",
    x"31AB8EA",
    x"31AB63C",
    x"31AB38F",
    x"31AB0E2",
    x"31AAE36",
    x"31AAB8B",
    x"31AA8E1",
    x"31AA637",
    x"31AA38E",
    x"31AA0E5",
    x"31A9E3D",
    x"31A9B96",
    x"31A98EF",
    x"31A9649",
    x"31A93A4",
    x"31A9100",
    x"31A8E5C",
    x"31A8BB8",
    x"31A8916",
    x"31A8674",
    x"31A83D3",
    x"31A8132",
    x"31A7E92",
    x"31A7BF3",
    x"31A7954",
    x"31A76B6",
    x"31A7419",
    x"31A717C",
    x"31A6EE0",
    x"31A6C44",
    x"31A69AA",
    x"31A6710",
    x"31A6476",
    x"31A61DD",
    x"31A5F45",
    x"31A5CAE",
    x"31A5A17",
    x"31A5781",
    x"31A54EB",
    x"31A5256",
    x"31A4FC2",
    x"31A4D2E",
    x"31A4A9B",
    x"31A4809",
    x"31A4577",
    x"31A42E6",
    x"31A4056",
    x"31A3DC6",
    x"31A3B37",
    x"31A38A9",
    x"31A361B",
    x"31A338E",
    x"31A3101",
    x"31A2E75",
    x"31A2BEA",
    x"31A295F",
    x"31A26D5",
    x"31A244C",
    x"31A21C3",
    x"31A1F3B",
    x"31A1CB3",
    x"31A1A2C",
    x"31A17A6",
    x"31A1521",
    x"31A129C",
    x"31A1017",
    x"31A0D94",
    x"31A0B10",
    x"31A088E",
    x"31A060C",
    x"31A038B",
    x"31A010A",
    x"319FE8A",
    x"319FC0B",
    x"319F98C",
    x"319F70E",
    x"319F491",
    x"319F214",
    x"319EF98",
    x"319ED1C",
    x"319EAA1",
    x"319E827",
    x"319E5AD",
    x"319E334",
    x"319E0BC",
    x"319DE44",
    x"319DBCD",
    x"319D956",
    x"319D6E0",
    x"319D46A",
    x"319D1F6",
    x"319CF81",
    x"319CD0E",
    x"319CA9B",
    x"319C829",
    x"319C5B7",
    x"319C346",
    x"319C0D5",
    x"319BE65",
    x"319BBF6",
    x"319B987",
    x"319B719",
    x"319B4AC",
    x"319B23F",
    x"319AFD3",
    x"319AD67",
    x"319AAFC",
    x"319A892",
    x"319A628",
    x"319A3BE",
    x"319A156",
    x"3199EEE",
    x"3199C86",
    x"3199A20",
    x"31997B9",
    x"3199554",
    x"31992EF",
    x"319908A",
    x"3198E26",
    x"3198BC3",
    x"3198960",
    x"31986FE",
    x"319849D",
    x"319823C",
    x"3197FDC",
    x"3197D7C",
    x"3197B1D",
    x"31978BF",
    x"3197661",
    x"3197403",
    x"31971A7",
    x"3196F4B",
    x"3196CEF",
    x"3196A94",
    x"319683A",
    x"31965E0",
    x"3196387",
    x"319612E",
    x"3195ED6",
    x"3195C7F",
    x"3195A28",
    x"31957D2",
    x"319557C",
    x"3195327",
    x"31950D3",
    x"3194E7F",
    x"3194C2B",
    x"31949D9",
    x"3194786",
    x"3194535",
    x"31942E4",
    x"3194093",
    x"3193E43",
    x"3193BF4",
    x"31939A5",
    x"3193757",
    x"319350A",
    x"31932BD",
    x"3193070",
    x"3192E25",
    x"3192BD9",
    x"319298F",
    x"3192745",
    x"31924FB",
    x"31922B2",
    x"319206A",
    x"3191E22",
    x"3191BDB",
    x"3191994",
    x"319174E",
    x"3191508",
    x"31912C3",
    x"319107F",
    x"3190E3B",
    x"3190BF8",
    x"31909B5",
    x"3190773",
    x"3190531",
    x"31902F0",
    x"31900B0",
    x"318FE70",
    x"318FC31",
    x"318F9F2",
    x"318F7B4",
    x"318F576",
    x"318F339",
    x"318F0FC",
    x"318EEC0",
    x"318EC85",
    x"318EA4A",
    x"318E810",
    x"318E5D6",
    x"318E39D",
    x"318E164",
    x"318DF2C",
    x"318DCF5",
    x"318DABE",
    x"318D887",
    x"318D652",
    x"318D41C",
    x"318D1E7",
    x"318CFB3",
    x"318CD80",
    x"318CB4D",
    x"318C91A",
    x"318C6E8",
    x"318C4B7",
    x"318C286",
    x"318C055",
    x"318BE25",
    x"318BBF6",
    x"318B9C7",
    x"318B799",
    x"318B56C",
    x"318B33F",
    x"318B112",
    x"318AEE6",
    x"318ACBB",
    x"318AA90",
    x"318A865",
    x"318A63C",
    x"318A412",
    x"318A1E9",
    x"3189FC1",
    x"3189D9A",
    x"3189B72",
    x"318994C",
    x"3189726",
    x"3189500",
    x"31892DB",
    x"31890B7",
    x"3188E93",
    x"3188C70",
    x"3188A4D",
    x"318882A",
    x"3188609",
    x"31883E7",
    x"31881C7",
    x"3187FA7",
    x"3187D87",
    x"3187B68",
    x"3187949",
    x"318772B",
    x"318750E",
    x"31872F1",
    x"31870D4",
    x"3186EB8",
    x"3186C9D",
    x"3186A82",
    x"3186867",
    x"318664E",
    x"3186434",
    x"318621C",
    x"3186003",
    x"3185DEC",
    x"3185BD4",
    x"31859BE",
    x"31857A7",
    x"3185592",
    x"318537D",
    x"3185168",
    x"3184F54",
    x"3184D40",
    x"3184B2D",
    x"318491B",
    x"3184709",
    x"31844F7",
    x"31842E6",
    x"31840D6",
    x"3183EC6",
    x"3183CB6",
    x"3183AA8",
    x"3183899",
    x"318368B",
    x"318347E",
    x"3183271",
    x"3183065",
    x"3182E59",
    x"3182C4D",
    x"3182A43",
    x"3182838",
    x"318262F",
    x"3182425",
    x"318221C",
    x"3182014",
    x"3181E0C",
    x"3181C05",
    x"31819FE",
    x"31817F8",
    x"31815F2",
    x"31813ED",
    x"31811E8",
    x"3180FE4",
    x"3180DE0",
    x"3180BDD",
    x"31809DB",
    x"31807D8",
    x"31805D7",
    x"31803D5",
    x"31801D5",
    x"317FFA9",
    x"317FBAA",
    x"317F7AC",
    x"317F3AE",
    x"317EFB2",
    x"317EBB6",
    x"317E7BC",
    x"317E3C3",
    x"317DFCA",
    x"317DBD3",
    x"317D7DC",
    x"317D3E7",
    x"317CFF2",
    x"317CBFF",
    x"317C80C",
    x"317C41B",
    x"317C02A",
    x"317BC3B",
    x"317B84C",
    x"317B45E",
    x"317B072",
    x"317AC86",
    x"317A89C",
    x"317A4B2",
    x"317A0C9",
    x"3179CE2",
    x"31798FB",
    x"3179515",
    x"3179130",
    x"3178D4C",
    x"317896A",
    x"3178588",
    x"31781A7",
    x"3177DC7",
    x"31779E8",
    x"317760A",
    x"317722D",
    x"3176E51",
    x"3176A76",
    x"317669C",
    x"31762C2",
    x"3175EEA",
    x"3175B13",
    x"317573D",
    x"3175367",
    x"3174F93",
    x"3174BC0",
    x"31747ED",
    x"317441C",
    x"317404B",
    x"3173C7B",
    x"31738AD",
    x"31734DF",
    x"3173112",
    x"3172D47",
    x"317297C",
    x"31725B2",
    x"31721E9",
    x"3171E21",
    x"3171A5A",
    x"3171694",
    x"31712CF",
    x"3170F0A",
    x"3170B47",
    x"3170785",
    x"31703C3",
    x"3170003",
    x"316FC43",
    x"316F885",
    x"316F4C7",
    x"316F10A",
    x"316ED4E",
    x"316E994",
    x"316E5DA",
    x"316E221",
    x"316DE69",
    x"316DAB1",
    x"316D6FB",
    x"316D346",
    x"316CF92",
    x"316CBDE",
    x"316C82C",
    x"316C47A",
    x"316C0C9",
    x"316BD1A",
    x"316B96B",
    x"316B5BD",
    x"316B210",
    x"316AE64",
    x"316AAB9",
    x"316A70F",
    x"316A365",
    x"3169FBD",
    x"3169C15",
    x"316986F",
    x"31694C9",
    x"3169124",
    x"3168D81",
    x"31689DE",
    x"316863C",
    x"316829B",
    x"3167EFA",
    x"3167B5B",
    x"31677BD",
    x"316741F",
    x"3167083",
    x"3166CE7",
    x"316694C",
    x"31665B2",
    x"3166219",
    x"3165E81",
    x"3165AEA",
    x"3165754",
    x"31653BE",
    x"316502A",
    x"3164C96",
    x"3164904",
    x"3164572",
    x"31641E1",
    x"3163E51",
    x"3163AC2",
    x"3163734",
    x"31633A6",
    x"316301A",
    x"3162C8E",
    x"3162903",
    x"316257A",
    x"31621F1",
    x"3161E69",
    x"3161AE2",
    x"316175B",
    x"31613D6",
    x"3161051",
    x"3160CCE",
    x"316094B",
    x"31605C9",
    x"3160248",
    x"315FEC8",
    x"315FB49",
    x"315F7CA",
    x"315F44D",
    x"315F0D0",
    x"315ED54",
    x"315E9D9",
    x"315E65F",
    x"315E2E6",
    x"315DF6E",
    x"315DBF7",
    x"315D880",
    x"315D50A",
    x"315D195",
    x"315CE21",
    x"315CAAE",
    x"315C73C",
    x"315C3CB",
    x"315C05A",
    x"315BCEB",
    x"315B97C",
    x"315B60E",
    x"315B2A1",
    x"315AF35",
    x"315ABC9",
    x"315A85F",
    x"315A4F5",
    x"315A18C",
    x"3159E24",
    x"3159ABD",
    x"3159757",
    x"31593F1",
    x"315908D",
    x"3158D29",
    x"31589C6",
    x"3158664",
    x"3158303",
    x"3157FA3",
    x"3157C43",
    x"31578E5",
    x"3157587",
    x"315722A",
    x"3156ECE",
    x"3156B72",
    x"3156818",
    x"31564BE",
    x"3156166",
    x"3155E0E",
    x"3155AB7",
    x"3155760",
    x"315540B",
    x"31550B6",
    x"3154D63",
    x"3154A10",
    x"31546BD",
    x"315436C",
    x"315401C",
    x"3153CCC",
    x"315397D",
    x"315362F",
    x"31532E2",
    x"3152F96",
    x"3152C4A",
    x"3152900",
    x"31525B6",
    x"315226D",
    x"3151F25",
    x"3151BDD",
    x"3151897",
    x"3151551",
    x"315120C",
    x"3150EC8",
    x"3150B85",
    x"3150842",
    x"3150501",
    x"31501C0",
    x"314FE80",
    x"314FB41",
    x"314F802",
    x"314F4C5",
    x"314F188",
    x"314EE4C",
    x"314EB11",
    x"314E7D6",
    x"314E49D",
    x"314E164",
    x"314DE2C",
    x"314DAF5",
    x"314D7BF",
    x"314D489",
    x"314D154",
    x"314CE20",
    x"314CAED",
    x"314C7BB",
    x"314C489",
    x"314C159",
    x"314BE29",
    x"314BAFA",
    x"314B7CB",
    x"314B49E",
    x"314B171",
    x"314AE45",
    x"314AB1A",
    x"314A7EF",
    x"314A4C6",
    x"314A19D",
    x"3149E75",
    x"3149B4E",
    x"3149827",
    x"3149502",
    x"31491DD",
    x"3148EB9",
    x"3148B95",
    x"3148873",
    x"3148551",
    x"3148230",
    x"3147F10",
    x"3147BF1",
    x"31478D2",
    x"31475B4",
    x"3147297",
    x"3146F7B",
    x"3146C60",
    x"3146945",
    x"314662B",
    x"3146312",
    x"3145FF9",
    x"3145CE2",
    x"31459CB",
    x"31456B5",
    x"31453A0",
    x"314508B",
    x"3144D77",
    x"3144A64",
    x"3144752",
    x"3144441",
    x"3144130",
    x"3143E20",
    x"3143B11",
    x"3143803",
    x"31434F5",
    x"31431E8",
    x"3142EDC",
    x"3142BD1",
    x"31428C6",
    x"31425BC",
    x"31422B3",
    x"3141FAB",
    x"3141CA3",
    x"314199D",
    x"3141697",
    x"3141391",
    x"314108D",
    x"3140D89",
    x"3140A86",
    x"3140784",
    x"3140482",
    x"3140181",
    x"313FE81",
    x"313FB82",
    x"313F884",
    x"313F586",
    x"313F289",
    x"313EF8D",
    x"313EC91",
    x"313E996",
    x"313E69C",
    x"313E3A3",
    x"313E0AB",
    x"313DDB3",
    x"313DABC",
    x"313D7C5",
    x"313D4D0",
    x"313D1DB",
    x"313CEE7",
    x"313CBF4",
    x"313C901",
    x"313C60F",
    x"313C31E",
    x"313C02D",
    x"313BD3E",
    x"313BA4F",
    x"313B761",
    x"313B473",
    x"313B186",
    x"313AE9A",
    x"313ABAF",
    x"313A8C5",
    x"313A5DB",
    x"313A2F2",
    x"313A009",
    x"3139D22",
    x"3139A3B",
    x"3139754",
    x"313946F",
    x"313918A",
    x"3138EA6",
    x"3138BC3",
    x"31388E0",
    x"31385FF",
    x"313831D",
    x"313803D",
    x"3137D5D",
    x"3137A7E",
    x"31377A0",
    x"31374C2",
    x"31371E6",
    x"3136F0A",
    x"3136C2E",
    x"3136953",
    x"3136679",
    x"31363A0",
    x"31360C8",
    x"3135DF0",
    x"3135B19",
    x"3135842",
    x"313556D",
    x"3135298",
    x"3134FC3",
    x"3134CF0",
    x"3134A1D",
    x"313474B",
    x"3134479",
    x"31341A8",
    x"3133ED8",
    x"3133C09",
    x"313393A",
    x"313366C",
    x"313339F",
    x"31330D2",
    x"3132E07",
    x"3132B3B",
    x"3132871",
    x"31325A7",
    x"31322DE",
    x"3132016",
    x"3131D4E",
    x"3131A87",
    x"31317C1",
    x"31314FB",
    x"3131236",
    x"3130F72",
    x"3130CAF",
    x"31309EC",
    x"313072A",
    x"3130468",
    x"31301A8",
    x"312FEE7",
    x"312FC28",
    x"312F969",
    x"312F6AB",
    x"312F3EE",
    x"312F131",
    x"312EE75",
    x"312EBBA",
    x"312E900",
    x"312E646",
    x"312E38C",
    x"312E0D4",
    x"312DE1C",
    x"312DB65",
    x"312D8AE",
    x"312D5F8",
    x"312D343",
    x"312D08F",
    x"312CDDB",
    x"312CB28",
    x"312C875",
    x"312C5C4",
    x"312C313",
    x"312C062",
    x"312BDB2",
    x"312BB03",
    x"312B855",
    x"312B5A7",
    x"312B2FA",
    x"312B04E",
    x"312ADA2",
    x"312AAF7",
    x"312A84C",
    x"312A5A3",
    x"312A2FA",
    x"312A051",
    x"3129DA9",
    x"3129B02",
    x"312985C",
    x"31295B6",
    x"3129311",
    x"312906D",
    x"3128DC9",
    x"3128B26",
    x"3128883",
    x"31285E1",
    x"3128340",
    x"31280A0",
    x"3127E00",
    x"3127B61",
    x"31278C2",
    x"3127624",
    x"3127387",
    x"31270EB",
    x"3126E4F",
    x"3126BB4",
    x"3126919",
    x"312667F",
    x"31263E6",
    x"312614D",
    x"3125EB5",
    x"3125C1E",
    x"3125987",
    x"31256F1",
    x"312545C",
    x"31251C7",
    x"3124F33",
    x"3124C9F",
    x"3124A0C",
    x"312477A",
    x"31244E9",
    x"3124258",
    x"3123FC7",
    x"3123D38",
    x"3123AA9",
    x"312381A",
    x"312358D",
    x"3123300",
    x"3123073",
    x"3122DE7",
    x"3122B5C",
    x"31228D2",
    x"3122648",
    x"31223BF",
    x"3122136",
    x"3121EAE",
    x"3121C27",
    x"31219A0",
    x"312171A",
    x"3121494",
    x"3121210",
    x"3120F8B",
    x"3120D08",
    x"3120A85",
    x"3120803",
    x"3120581",
    x"3120300",
    x"312007F",
    x"311FE00",
    x"311FB80",
    x"311F902",
    x"311F684",
    x"311F407",
    x"311F18A",
    x"311EF0E",
    x"311EC92",
    x"311EA17",
    x"311E79D",
    x"311E524",
    x"311E2AB",
    x"311E032",
    x"311DDBB",
    x"311DB43",
    x"311D8CD",
    x"311D657",
    x"311D3E2",
    x"311D16D",
    x"311CEF9",
    x"311CC86",
    x"311CA13",
    x"311C7A1",
    x"311C52F",
    x"311C2BE",
    x"311C04E",
    x"311BDDE",
    x"311BB6F",
    x"311B900",
    x"311B692",
    x"311B425",
    x"311B1B8",
    x"311AF4C",
    x"311ACE0",
    x"311AA76",
    x"311A80B",
    x"311A5A2",
    x"311A338",
    x"311A0D0",
    x"3119E68",
    x"3119C01",
    x"311999A",
    x"3119734",
    x"31194CE",
    x"3119269",
    x"3119005",
    x"3118DA1",
    x"3118B3E",
    x"31188DC",
    x"311867A",
    x"3118419",
    x"31181B8",
    x"3117F58",
    x"3117CF8",
    x"3117A99",
    x"311783B",
    x"31175DD",
    x"3117380",
    x"3117123",
    x"3116EC7",
    x"3116C6C",
    x"3116A11",
    x"31167B7",
    x"311655D",
    x"3116304",
    x"31160AC",
    x"3115E54",
    x"3115BFD",
    x"31159A6",
    x"3115750",
    x"31154FA",
    x"31152A5",
    x"3115051",
    x"3114DFD",
    x"3114BAA",
    x"3114957",
    x"3114705",
    x"31144B4",
    x"3114263",
    x"3114013",
    x"3113DC3",
    x"3113B74",
    x"3113925",
    x"31136D7",
    x"311348A",
    x"311323D",
    x"3112FF1",
    x"3112DA5",
    x"3112B5A",
    x"311290F",
    x"31126C5",
    x"311247C",
    x"3112233",
    x"3111FEB",
    x"3111DA3",
    x"3111B5C",
    x"3111915",
    x"31116CF",
    x"311148A",
    x"3111245",
    x"3111001",
    x"3110DBD",
    x"3110B7A",
    x"3110937",
    x"31106F5",
    x"31104B4",
    x"3110273",
    x"3110033",
    x"310FDF3",
    x"310FBB4",
    x"310F975",
    x"310F737",
    x"310F4F9",
    x"310F2BD",
    x"310F080",
    x"310EE44",
    x"310EC09",
    x"310E9CE",
    x"310E794",
    x"310E55A",
    x"310E321",
    x"310E0E9",
    x"310DEB1",
    x"310DC7A",
    x"310DA43",
    x"310D80C",
    x"310D5D7",
    x"310D3A1",
    x"310D16D",
    x"310CF39",
    x"310CD05",
    x"310CAD2",
    x"310C8A0",
    x"310C66E",
    x"310C43D",
    x"310C20C",
    x"310BFDC",
    x"310BDAC",
    x"310BB7D",
    x"310B94E",
    x"310B720",
    x"310B4F3",
    x"310B2C6",
    x"310B099",
    x"310AE6D",
    x"310AC42",
    x"310AA17",
    x"310A7ED",
    x"310A5C3",
    x"310A39A",
    x"310A171",
    x"3109F49",
    x"3109D22",
    x"3109AFB",
    x"31098D4",
    x"31096AE",
    x"3109489",
    x"3109264",
    x"3109040",
    x"3108E1C",
    x"3108BF9",
    x"31089D6",
    x"31087B4",
    x"3108592",
    x"3108371",
    x"3108150",
    x"3107F30",
    x"3107D11",
    x"3107AF2",
    x"31078D3",
    x"31076B5",
    x"3107498",
    x"310727B",
    x"310705F",
    x"3106E43",
    x"3106C28",
    x"3106A0D",
    x"31067F3",
    x"31065D9",
    x"31063C0",
    x"31061A7",
    x"3105F8F",
    x"3105D77",
    x"3105B60",
    x"310594A",
    x"3105733",
    x"310551E",
    x"3105309",
    x"31050F4",
    x"3104EE0",
    x"3104CCD",
    x"3104ABA",
    x"31048A8",
    x"3104696",
    x"3104484",
    x"3104273",
    x"3104063",
    x"3103E53",
    x"3103C44",
    x"3103A35",
    x"3103827",
    x"3103619",
    x"310340C",
    x"31031FF",
    x"3102FF3",
    x"3102DE7",
    x"3102BDC",
    x"31029D1",
    x"31027C7",
    x"31025BD",
    x"31023B4",
    x"31021AB",
    x"3101FA3",
    x"3101D9C",
    x"3101B94",
    x"310198E",
    x"3101788",
    x"3101582",
    x"310137D",
    x"3101178",
    x"3100F74",
    x"3100D70",
    x"3100B6D",
    x"310096B",
    x"3100769",
    x"3100567",
    x"3100366",
    x"3100165",
    x"30FFECB",
    x"30FFACC",
    x"30FF6CE",
    x"30FF2D0",
    x"30FEED4",
    x"30FEAD9",
    x"30FE6DF",
    x"30FE2E6",
    x"30FDEED",
    x"30FDAF6",
    x"30FD700",
    x"30FD30B",
    x"30FCF16",
    x"30FCB23",
    x"30FC731",
    x"30FC33F",
    x"30FBF4F",
    x"30FBB60",
    x"30FB771",
    x"30FB384",
    x"30FAF98",
    x"30FABAC",
    x"30FA7C2",
    x"30FA3D8",
    x"30F9FF0",
    x"30F9C08",
    x"30F9822",
    x"30F943C",
    x"30F9058",
    x"30F8C74",
    x"30F8892",
    x"30F84B0",
    x"30F80CF",
    x"30F7CF0",
    x"30F7911",
    x"30F7533",
    x"30F7156",
    x"30F6D7A",
    x"30F699F",
    x"30F65C5",
    x"30F61ED",
    x"30F5E15",
    x"30F5A3D",
    x"30F5667",
    x"30F5292",
    x"30F4EBE",
    x"30F4AEB",
    x"30F4719",
    x"30F4347",
    x"30F3F77",
    x"30F3BA8",
    x"30F37D9",
    x"30F340C",
    x"30F303F",
    x"30F2C74",
    x"30F28A9",
    x"30F24DF",
    x"30F2116",
    x"30F1D4F",
    x"30F1988",
    x"30F15C2",
    x"30F11FD",
    x"30F0E39",
    x"30F0A76",
    x"30F06B4",
    x"30F02F2",
    x"30EFF32",
    x"30EFB73",
    x"30EF7B5",
    x"30EF3F7",
    x"30EF03B",
    x"30EEC7F",
    x"30EE8C4",
    x"30EE50B",
    x"30EE152",
    x"30EDD9A",
    x"30ED9E3",
    x"30ED62D",
    x"30ED278",
    x"30ECEC4",
    x"30ECB10",
    x"30EC75E",
    x"30EC3AD",
    x"30EBFFC",
    x"30EBC4D",
    x"30EB89E",
    x"30EB4F0",
    x"30EB144",
    x"30EAD98",
    x"30EA9ED",
    x"30EA643",
    x"30EA29A",
    x"30E9EF2",
    x"30E9B4A",
    x"30E97A4",
    x"30E93FE",
    x"30E905A",
    x"30E8CB6",
    x"30E8914",
    x"30E8572",
    x"30E81D1",
    x"30E7E31",
    x"30E7A92",
    x"30E76F4",
    x"30E7356",
    x"30E6FBA",
    x"30E6C1E",
    x"30E6884",
    x"30E64EA",
    x"30E6151",
    x"30E5DBA",
    x"30E5A23",
    x"30E568C",
    x"30E52F7",
    x"30E4F63",
    x"30E4BD0",
    x"30E483D",
    x"30E44AB",
    x"30E411B",
    x"30E3D8B",
    x"30E39FC",
    x"30E366E",
    x"30E32E1",
    x"30E2F54",
    x"30E2BC9",
    x"30E283F",
    x"30E24B5",
    x"30E212C",
    x"30E1DA4",
    x"30E1A1D",
    x"30E1697",
    x"30E1312",
    x"30E0F8E",
    x"30E0C0A",
    x"30E0888",
    x"30E0506",
    x"30E0185",
    x"30DFE05",
    x"30DFA86",
    x"30DF708",
    x"30DF38B",
    x"30DF00E",
    x"30DEC93",
    x"30DE918",
    x"30DE59E",
    x"30DE225",
    x"30DDEAD",
    x"30DDB36",
    x"30DD7BF",
    x"30DD44A",
    x"30DD0D5",
    x"30DCD62",
    x"30DC9EF",
    x"30DC67D",
    x"30DC30B",
    x"30DBF9B",
    x"30DBC2C",
    x"30DB8BD",
    x"30DB54F",
    x"30DB1E2",
    x"30DAE76",
    x"30DAB0B",
    x"30DA7A1",
    x"30DA437",
    x"30DA0CF",
    x"30D9D67",
    x"30D9A00",
    x"30D969A",
    x"30D9335",
    x"30D8FD0",
    x"30D8C6D",
    x"30D890A",
    x"30D85A8",
    x"30D8247",
    x"30D7EE7",
    x"30D7B88",
    x"30D7829",
    x"30D74CC",
    x"30D716F",
    x"30D6E13",
    x"30D6AB8",
    x"30D675E",
    x"30D6404",
    x"30D60AC",
    x"30D5D54",
    x"30D59FD",
    x"30D56A7",
    x"30D5352",
    x"30D4FFD",
    x"30D4CAA",
    x"30D4957",
    x"30D4605",
    x"30D42B4",
    x"30D3F64",
    x"30D3C14",
    x"30D38C5",
    x"30D3578",
    x"30D322B",
    x"30D2EDF",
    x"30D2B93",
    x"30D2849",
    x"30D24FF",
    x"30D21B6",
    x"30D1E6E",
    x"30D1B27",
    x"30D17E1",
    x"30D149B",
    x"30D1156",
    x"30D0E13",
    x"30D0ACF",
    x"30D078D",
    x"30D044C",
    x"30D010B",
    x"30CFDCB",
    x"30CFA8C",
    x"30CF74E",
    x"30CF410",
    x"30CF0D4",
    x"30CED98",
    x"30CEA5D",
    x"30CE723",
    x"30CE3E9",
    x"30CE0B1",
    x"30CDD79",
    x"30CDA42",
    x"30CD70C",
    x"30CD3D7",
    x"30CD0A2",
    x"30CCD6E",
    x"30CCA3B",
    x"30CC709",
    x"30CC3D8",
    x"30CC0A7",
    x"30CBD77",
    x"30CBA49",
    x"30CB71A",
    x"30CB3ED",
    x"30CB0C0",
    x"30CAD95",
    x"30CAA6A",
    x"30CA73F",
    x"30CA416",
    x"30CA0ED",
    x"30C9DC5",
    x"30C9A9E",
    x"30C9778",
    x"30C9453",
    x"30C912E",
    x"30C8E0A",
    x"30C8AE7",
    x"30C87C5",
    x"30C84A3",
    x"30C8182",
    x"30C7E62",
    x"30C7B43",
    x"30C7825",
    x"30C7507",
    x"30C71EA",
    x"30C6ECE",
    x"30C6BB3",
    x"30C6898",
    x"30C657F",
    x"30C6266",
    x"30C5F4D",
    x"30C5C36",
    x"30C591F",
    x"30C5609",
    x"30C52F4",
    x"30C4FE0",
    x"30C4CCC",
    x"30C49B9",
    x"30C46A7",
    x"30C4396",
    x"30C4086",
    x"30C3D76",
    x"30C3A67",
    x"30C3759",
    x"30C344B",
    x"30C313E",
    x"30C2E33",
    x"30C2B27",
    x"30C281D",
    x"30C2513",
    x"30C220A",
    x"30C1F02",
    x"30C1BFB",
    x"30C18F4",
    x"30C15EE",
    x"30C12E9",
    x"30C0FE5",
    x"30C0CE1",
    x"30C09DF",
    x"30C06DC",
    x"30C03DB",
    x"30C00DB",
    x"30BFDDB",
    x"30BFADC",
    x"30BF7DD",
    x"30BF4E0",
    x"30BF1E3",
    x"30BEEE7",
    x"30BEBEB",
    x"30BE8F1",
    x"30BE5F7",
    x"30BE2FE",
    x"30BE005",
    x"30BDD0E",
    x"30BDA17",
    x"30BD721",
    x"30BD42B",
    x"30BD137",
    x"30BCE43",
    x"30BCB50",
    x"30BC85D",
    x"30BC56B",
    x"30BC27A",
    x"30BBF8A",
    x"30BBC9B",
    x"30BB9AC",
    x"30BB6BE",
    x"30BB3D0",
    x"30BB0E4",
    x"30BADF8",
    x"30BAB0D",
    x"30BA822",
    x"30BA539",
    x"30BA250",
    x"30B9F68",
    x"30B9C80",
    x"30B9999",
    x"30B96B3",
    x"30B93CE",
    x"30B90E9",
    x"30B8E06",
    x"30B8B22",
    x"30B8840",
    x"30B855E",
    x"30B827D",
    x"30B7F9D",
    x"30B7CBD",
    x"30B79DF",
    x"30B7701",
    x"30B7423",
    x"30B7146",
    x"30B6E6B",
    x"30B6B8F",
    x"30B68B5",
    x"30B65DB",
    x"30B6302",
    x"30B6029",
    x"30B5D52",
    x"30B5A7B",
    x"30B57A4",
    x"30B54CF",
    x"30B51FA",
    x"30B4F26",
    x"30B4C53",
    x"30B4980",
    x"30B46AE",
    x"30B43DC",
    x"30B410C",
    x"30B3E3C",
    x"30B3B6D",
    x"30B389E",
    x"30B35D0",
    x"30B3303",
    x"30B3037",
    x"30B2D6B",
    x"30B2AA0",
    x"30B27D6",
    x"30B250C",
    x"30B2243",
    x"30B1F7B",
    x"30B1CB4",
    x"30B19ED",
    x"30B1727",
    x"30B1461",
    x"30B119C",
    x"30B0ED8",
    x"30B0C15",
    x"30B0952",
    x"30B0690",
    x"30B03CF",
    x"30B010E",
    x"30AFE4F",
    x"30AFB8F",
    x"30AF8D1",
    x"30AF613",
    x"30AF356",
    x"30AF099",
    x"30AEDDD",
    x"30AEB22",
    x"30AE868",
    x"30AE5AE",
    x"30AE2F5",
    x"30AE03D",
    x"30ADD85",
    x"30ADACE",
    x"30AD817",
    x"30AD562",
    x"30AD2AD",
    x"30ACFF8",
    x"30ACD45",
    x"30ACA92",
    x"30AC7E0",
    x"30AC52E",
    x"30AC27D",
    x"30ABFCD",
    x"30ABD1D",
    x"30ABA6E",
    x"30AB7C0",
    x"30AB512",
    x"30AB265",
    x"30AAFB9",
    x"30AAD0D",
    x"30AAA62",
    x"30AA7B8",
    x"30AA50F",
    x"30AA266",
    x"30A9FBD",
    x"30A9D16",
    x"30A9A6F",
    x"30A97C9",
    x"30A9523",
    x"30A927E",
    x"30A8FDA",
    x"30A8D36",
    x"30A8A93",
    x"30A87F1",
    x"30A854F",
    x"30A82AE",
    x"30A800E",
    x"30A7D6E",
    x"30A7ACF",
    x"30A7831",
    x"30A7593",
    x"30A72F6",
    x"30A705A",
    x"30A6DBE",
    x"30A6B23",
    x"30A6888",
    x"30A65EE",
    x"30A6355",
    x"30A60BD",
    x"30A5E25",
    x"30A5B8E",
    x"30A58F7",
    x"30A5661",
    x"30A53CC",
    x"30A5137",
    x"30A4EA3",
    x"30A4C10",
    x"30A497D",
    x"30A46EB",
    x"30A445A",
    x"30A41C9",
    x"30A3F39",
    x"30A3CA9",
    x"30A3A1B",
    x"30A378C",
    x"30A34FF",
    x"30A3272",
    x"30A2FE6",
    x"30A2D5A",
    x"30A2ACF",
    x"30A2845",
    x"30A25BB",
    x"30A2332",
    x"30A20A9",
    x"30A1E21",
    x"30A1B9A",
    x"30A1914",
    x"30A168E",
    x"30A1408",
    x"30A1184",
    x"30A0EFF",
    x"30A0C7C",
    x"30A09F9",
    x"30A0777",
    x"30A04F5",
    x"30A0275",
    x"309FFF4",
    x"309FD75",
    x"309FAF6",
    x"309F877",
    x"309F5F9",
    x"309F37C",
    x"309F100",
    x"309EE84",
    x"309EC08",
    x"309E98E",
    x"309E714",
    x"309E49A",
    x"309E221",
    x"309DFA9",
    x"309DD31",
    x"309DABA",
    x"309D844",
    x"309D5CE",
    x"309D359",
    x"309D0E5",
    x"309CE71",
    x"309CBFD",
    x"309C98B",
    x"309C719",
    x"309C4A7",
    x"309C236",
    x"309BFC6",
    x"309BD56",
    x"309BAE7",
    x"309B879",
    x"309B60B",
    x"309B39E",
    x"309B131",
    x"309AEC5",
    x"309AC5A",
    x"309A9EF",
    x"309A785",
    x"309A51B",
    x"309A2B2",
    x"309A04A",
    x"3099DE2",
    x"3099B7B",
    x"3099915",
    x"30996AF",
    x"3099449",
    x"30991E4",
    x"3098F80",
    x"3098D1D",
    x"3098ABA",
    x"3098857",
    x"30985F5",
    x"3098394",
    x"3098134",
    x"3097ED4",
    x"3097C74",
    x"3097A15",
    x"30977B7",
    x"309755A",
    x"30972FD",
    x"30970A0",
    x"3096E44",
    x"3096BE9",
    x"309698E",
    x"3096734",
    x"30964DB",
    x"3096282",
    x"3096029",
    x"3095DD2",
    x"3095B7B",
    x"3095924",
    x"30956CE",
    x"3095479",
    x"3095224",
    x"3094FCF",
    x"3094D7C",
    x"3094B29",
    x"30948D6",
    x"3094684",
    x"3094433",
    x"30941E2",
    x"3093F92",
    x"3093D42",
    x"3093AF3",
    x"30938A5",
    x"3093657",
    x"309340A",
    x"30931BD",
    x"3092F71",
    x"3092D25",
    x"3092ADA",
    x"3092890",
    x"3092646",
    x"30923FD",
    x"30921B4",
    x"3091F6C",
    x"3091D24",
    x"3091ADD",
    x"3091897",
    x"3091651",
    x"309140C",
    x"30911C7",
    x"3090F83",
    x"3090D3F",
    x"3090AFC",
    x"30908BA",
    x"3090678",
    x"3090437",
    x"30901F6",
    x"308FFB6",
    x"308FD76",
    x"308FB37",
    x"308F8F8",
    x"308F6BA",
    x"308F47D",
    x"308F240",
    x"308F004",
    x"308EDC8",
    x"308EB8D",
    x"308E952",
    x"308E718",
    x"308E4DF",
    x"308E2A6",
    x"308E06D",
    x"308DE36",
    x"308DBFE",
    x"308D9C8",
    x"308D791",
    x"308D55C",
    x"308D327",
    x"308D0F2",
    x"308CEBE",
    x"308CC8B",
    x"308CA58",
    x"308C826",
    x"308C5F4",
    x"308C3C3",
    x"308C192",
    x"308BF62",
    x"308BD32",
    x"308BB03",
    x"308B8D5",
    x"308B6A7",
    x"308B47A",
    x"308B24D",
    x"308B020",
    x"308ADF5",
    x"308ABC9",
    x"308A99F",
    x"308A775",
    x"308A54B",
    x"308A322",
    x"308A0F9",
    x"3089ED1",
    x"3089CAA",
    x"3089A83",
    x"308985D",
    x"3089637",
    x"3089412",
    x"30891ED",
    x"3088FC9",
    x"3088DA5",
    x"3088B82",
    x"308895F",
    x"308873D",
    x"308851C",
    x"30882FB",
    x"30880DA",
    x"3087EBA",
    x"3087C9B",
    x"3087A7C",
    x"308785E",
    x"3087640",
    x"3087422",
    x"3087206",
    x"3086FE9",
    x"3086DCE",
    x"3086BB2",
    x"3086998",
    x"308677E",
    x"3086564",
    x"308634B",
    x"3086132",
    x"3085F1A",
    x"3085D03",
    x"3085AEC",
    x"30858D5",
    x"30856BF",
    x"30854AA",
    x"3085295",
    x"3085081",
    x"3084E6D",
    x"3084C5A",
    x"3084A47",
    x"3084834",
    x"3084623",
    x"3084411",
    x"3084201",
    x"3083FF0",
    x"3083DE1",
    x"3083BD1",
    x"30839C3",
    x"30837B5",
    x"30835A7",
    x"308339A",
    x"308318D",
    x"3082F81",
    x"3082D75",
    x"3082B6A",
    x"3082960",
    x"3082755",
    x"308254C",
    x"3082343",
    x"308213A",
    x"3081F32",
    x"3081D2B",
    x"3081B24",
    x"308191D",
    x"3081717",
    x"3081512",
    x"308130D",
    x"3081108",
    x"3080F04",
    x"3080D01",
    x"3080AFE",
    x"30808FB",
    x"30806F9",
    x"30804F8",
    x"30802F7",
    x"30800F6",
    x"307FDED",
    x"307F9EE",
    x"307F5F0",
    x"307F1F3",
    x"307EDF7",
    x"307E9FC",
    x"307E602",
    x"307E209",
    x"307DE11",
    x"307DA1A",
    x"307D624",
    x"307D22F",
    x"307CE3B",
    x"307CA47",
    x"307C655",
    x"307C264",
    x"307BE74",
    x"307BA85",
    x"307B697",
    x"307B2AA",
    x"307AEBE",
    x"307AAD2",
    x"307A6E8",
    x"307A2FF",
    x"3079F17",
    x"3079B2F",
    x"3079749",
    x"3079364",
    x"3078F7F",
    x"3078B9C",
    x"30787BA",
    x"30783D8",
    x"3077FF8",
    x"3077C18",
    x"307783A",
    x"307745C",
    x"307707F",
    x"3076CA4",
    x"30768C9",
    x"30764EF",
    x"3076117",
    x"3075D3F",
    x"3075968",
    x"3075592",
    x"30751BD",
    x"3074DE9",
    x"3074A16",
    x"3074644",
    x"3074273",
    x"3073EA3",
    x"3073AD4",
    x"3073706",
    x"3073338",
    x"3072F6C",
    x"3072BA1",
    x"30727D6",
    x"307240D",
    x"3072044",
    x"3071C7D",
    x"30718B6",
    x"30714F0",
    x"307112B",
    x"3070D68",
    x"30709A5",
    x"30705E3",
    x"3070222",
    x"306FE62",
    x"306FAA3",
    x"306F6E4",
    x"306F327",
    x"306EF6B",
    x"306EBAF",
    x"306E7F5",
    x"306E43B",
    x"306E083",
    x"306DCCB",
    x"306D914",
    x"306D55F",
    x"306D1AA",
    x"306CDF6",
    x"306CA43",
    x"306C691",
    x"306C2DF",
    x"306BF2F",
    x"306BB80",
    x"306B7D1",
    x"306B424",
    x"306B077",
    x"306ACCC",
    x"306A921",
    x"306A577",
    x"306A1CE",
    x"3069E26",
    x"3069A7F",
    x"30696D9",
    x"3069334",
    x"3068F8F",
    x"3068BEC",
    x"3068849",
    x"30684A8",
    x"3068107",
    x"3067D67",
    x"30679C8",
    x"306762A",
    x"306728D",
    x"3066EF1",
    x"3066B56",
    x"30667BB",
    x"3066422",
    x"3066089",
    x"3065CF2",
    x"306595B",
    x"30655C5",
    x"3065230",
    x"3064E9C",
    x"3064B09",
    x"3064776",
    x"30643E5",
    x"3064055",
    x"3063CC5",
    x"3063936",
    x"30635A8",
    x"306321B",
    x"3062E8F",
    x"3062B04",
    x"306277A",
    x"30623F0",
    x"3062068",
    x"3061CE0",
    x"3061959",
    x"30615D3",
    x"306124E",
    x"3060ECA",
    x"3060B47",
    x"30607C5",
    x"3060443",
    x"30600C2",
    x"305FD43",
    x"305F9C4",
    x"305F646",
    x"305F2C9",
    x"305EF4C",
    x"305EBD1",
    x"305E857",
    x"305E4DD",
    x"305E164",
    x"305DDEC",
    x"305DA75",
    x"305D6FF",
    x"305D38A",
    x"305D015",
    x"305CCA2",
    x"305C92F",
    x"305C5BD",
    x"305C24C",
    x"305BEDC",
    x"305BB6D",
    x"305B7FE",
    x"305B491",
    x"305B124",
    x"305ADB8",
    x"305AA4D",
    x"305A6E3",
    x"305A37A",
    x"305A011",
    x"3059CAA",
    x"3059943",
    x"30595DD",
    x"3059278",
    x"3058F14",
    x"3058BB0",
    x"305884E",
    x"30584EC",
    x"305818B",
    x"3057E2B",
    x"3057ACC",
    x"305776E",
    x"3057411",
    x"30570B4",
    x"3056D58",
    x"30569FD",
    x"30566A3",
    x"305634A",
    x"3055FF2",
    x"3055C9A",
    x"3055943",
    x"30555ED",
    x"3055298",
    x"3054F44",
    x"3054BF1",
    x"305489E",
    x"305454C",
    x"30541FB",
    x"3053EAB",
    x"3053B5C",
    x"305380E",
    x"30534C0",
    x"3053173",
    x"3052E27",
    x"3052ADC",
    x"3052792",
    x"3052448",
    x"3052100",
    x"3051DB8",
    x"3051A71",
    x"305172B",
    x"30513E5",
    x"30510A1",
    x"3050D5D",
    x"3050A1A",
    x"30506D8",
    x"3050397",
    x"3050056",
    x"304FD16",
    x"304F9D8",
    x"304F69A",
    x"304F35C",
    x"304F020",
    x"304ECE4",
    x"304E9A9",
    x"304E66F",
    x"304E336",
    x"304DFFE",
    x"304DCC6",
    x"304D98F",
    x"304D659",
    x"304D324",
    x"304CFF0",
    x"304CCBC",
    x"304C989",
    x"304C657",
    x"304C326",
    x"304BFF6",
    x"304BCC6",
    x"304B998",
    x"304B66A",
    x"304B33C",
    x"304B010",
    x"304ACE4",
    x"304A9B9",
    x"304A68F",
    x"304A366",
    x"304A03E",
    x"3049D16",
    x"30499EF",
    x"30496C9",
    x"30493A4",
    x"304907F",
    x"3048D5C",
    x"3048A39",
    x"3048716",
    x"30483F5",
    x"30480D4",
    x"3047DB5",
    x"3047A96",
    x"3047777",
    x"304745A",
    x"304713D",
    x"3046E21",
    x"3046B06",
    x"30467EC",
    x"30464D2",
    x"30461B9",
    x"3045EA1",
    x"3045B8A",
    x"3045873",
    x"304555E",
    x"3045249",
    x"3044F35",
    x"3044C21",
    x"304490F",
    x"30445FD",
    x"30442EC",
    x"3043FDB",
    x"3043CCC",
    x"30439BD",
    x"30436AF",
    x"30433A1",
    x"3043095",
    x"3042D89",
    x"3042A7E",
    x"3042774",
    x"304246A",
    x"3042162",
    x"3041E5A",
    x"3041B53",
    x"304184C",
    x"3041546",
    x"3041241",
    x"3040F3D",
    x"3040C3A",
    x"3040937",
    x"3040635",
    x"3040334",
    x"3040034",
    x"303FD34",
    x"303FA35",
    x"303F737",
    x"303F439",
    x"303F13D",
    x"303EE41",
    x"303EB46",
    x"303E84B",
    x"303E551",
    x"303E258",
    x"303DF60",
    x"303DC69",
    x"303D972",
    x"303D67C",
    x"303D387",
    x"303D092",
    x"303CD9F",
    x"303CAAC",
    x"303C7B9",
    x"303C4C8",
    x"303C1D7",
    x"303BEE7",
    x"303BBF7",
    x"303B909",
    x"303B61B",
    x"303B32E",
    x"303B041",
    x"303AD56",
    x"303AA6B",
    x"303A780",
    x"303A497",
    x"303A1AE",
    x"3039EC6",
    x"3039BDF",
    x"30398F8",
    x"3039612",
    x"303932D",
    x"3039049",
    x"3038D65",
    x"3038A82",
    x"30387A0",
    x"30384BE",
    x"30381DD",
    x"3037EFD",
    x"3037C1E",
    x"303793F",
    x"3037661",
    x"3037384",
    x"30370A7",
    x"3036DCC",
    x"3036AF0",
    x"3036816",
    x"303653C",
    x"3036263",
    x"3035F8B",
    x"3035CB4",
    x"30359DD",
    x"3035707",
    x"3035431",
    x"303515D",
    x"3034E89",
    x"3034BB5",
    x"30348E3",
    x"3034611",
    x"3034340",
    x"303406F",
    x"3033DA0",
    x"3033AD1",
    x"3033802",
    x"3033535",
    x"3033268",
    x"3032F9B",
    x"3032CD0",
    x"3032A05",
    x"303273B",
    x"3032471",
    x"30321A9",
    x"3031EE0",
    x"3031C19",
    x"3031952",
    x"303168C",
    x"30313C7",
    x"3031103",
    x"3030E3F",
    x"3030B7B",
    x"30308B9",
    x"30305F7",
    x"3030336",
    x"3030075",
    x"302FDB6",
    x"302FAF7",
    x"302F838",
    x"302F57A",
    x"302F2BD",
    x"302F001",
    x"302ED45",
    x"302EA8A",
    x"302E7D0",
    x"302E517",
    x"302E25E",
    x"302DFA5",
    x"302DCEE",
    x"302DA37",
    x"302D781",
    x"302D4CB",
    x"302D216",
    x"302CF62",
    x"302CCAF",
    x"302C9FC",
    x"302C74A",
    x"302C498",
    x"302C1E7",
    x"302BF37",
    x"302BC88",
    x"302B9D9",
    x"302B72B",
    x"302B47D",
    x"302B1D1",
    x"302AF24",
    x"302AC79",
    x"302A9CE",
    x"302A724",
    x"302A47B",
    x"302A1D2",
    x"3029F2A",
    x"3029C82",
    x"30299DB",
    x"3029735",
    x"3029490",
    x"30291EB",
    x"3028F47",
    x"3028CA3",
    x"3028A01",
    x"302875E",
    x"30284BD",
    x"302821C",
    x"3027F7C",
    x"3027CDC",
    x"3027A3D",
    x"302779F",
    x"3027502",
    x"3027265",
    x"3026FC8",
    x"3026D2D",
    x"3026A92",
    x"30267F7",
    x"302655E",
    x"30262C5",
    x"302602C",
    x"3025D95",
    x"3025AFE",
    x"3025867",
    x"30255D1",
    x"302533C",
    x"30250A8",
    x"3024E14",
    x"3024B81",
    x"30248EE",
    x"302465C",
    x"30243CB",
    x"302413A",
    x"3023EAA",
    x"3023C1B",
    x"302398C",
    x"30236FE",
    x"3023471",
    x"30231E4",
    x"3022F58",
    x"3022CCC",
    x"3022A42",
    x"30227B7",
    x"302252E",
    x"30222A5",
    x"302201C",
    x"3021D95",
    x"3021B0E",
    x"3021887",
    x"3021601",
    x"302137C",
    x"30210F8",
    x"3020E74",
    x"3020BF0",
    x"302096E",
    x"30206EC",
    x"302046A",
    x"30201E9",
    x"301FF69",
    x"301FCEA",
    x"301FA6B",
    x"301F7EC",
    x"301F56F",
    x"301F2F2",
    x"301F075",
    x"301EDFA",
    x"301EB7E",
    x"301E904",
    x"301E68A",
    x"301E410",
    x"301E198",
    x"301DF20",
    x"301DCA8",
    x"301DA31",
    x"301D7BB",
    x"301D546",
    x"301D2D0",
    x"301D05C",
    x"301CDE8",
    x"301CB75",
    x"301C903",
    x"301C691",
    x"301C41F",
    x"301C1AF",
    x"301BF3E",
    x"301BCCF",
    x"301BA60",
    x"301B7F2",
    x"301B584",
    x"301B317",
    x"301B0AB",
    x"301AE3F",
    x"301ABD3",
    x"301A969",
    x"301A6FF",
    x"301A495",
    x"301A22C",
    x"3019FC4",
    x"3019D5D",
    x"3019AF5",
    x"301988F",
    x"3019629",
    x"30193C4",
    x"301915F",
    x"3018EFB",
    x"3018C98",
    x"3018A35",
    x"30187D3",
    x"3018571",
    x"3018310",
    x"30180B0",
    x"3017E50",
    x"3017BF0",
    x"3017992",
    x"3017734",
    x"30174D6",
    x"3017279",
    x"301701D",
    x"3016DC1",
    x"3016B66",
    x"301690B",
    x"30166B1",
    x"3016458",
    x"30161FF",
    x"3015FA7",
    x"3015D4F",
    x"3015AF8",
    x"30158A2",
    x"301564C",
    x"30153F7",
    x"30151A2",
    x"3014F4E",
    x"3014CFA",
    x"3014AA8",
    x"3014855",
    x"3014603",
    x"30143B2",
    x"3014161",
    x"3013F11",
    x"3013CC2",
    x"3013A73",
    x"3013825",
    x"30135D7",
    x"301338A",
    x"301313D",
    x"3012EF1",
    x"3012CA6",
    x"3012A5B",
    x"3012811",
    x"30125C7",
    x"301237E",
    x"3012135",
    x"3011EED",
    x"3011CA6",
    x"3011A5F",
    x"3011818",
    x"30115D3",
    x"301138E",
    x"3011149",
    x"3010F05",
    x"3010CC1",
    x"3010A7E",
    x"301083C",
    x"30105FA",
    x"30103B9",
    x"3010179",
    x"300FF38",
    x"300FCF9",
    x"300FABA",
    x"300F87C",
    x"300F63E",
    x"300F400",
    x"300F1C4",
    x"300EF88",
    x"300ED4C",
    x"300EB11",
    x"300E8D6",
    x"300E69C",
    x"300E463",
    x"300E22A",
    x"300DFF2",
    x"300DDBA",
    x"300DB83",
    x"300D94D",
    x"300D716",
    x"300D4E1",
    x"300D2AC",
    x"300D078",
    x"300CE44",
    x"300CC11",
    x"300C9DE",
    x"300C7AC",
    x"300C57A",
    x"300C349",
    x"300C118",
    x"300BEE8",
    x"300BCB9",
    x"300BA8A",
    x"300B85C",
    x"300B62E",
    x"300B400",
    x"300B1D4",
    x"300AFA8",
    x"300AD7C",
    x"300AB51",
    x"300A926",
    x"300A6FC",
    x"300A4D3",
    x"300A2AA",
    x"300A081",
    x"3009E5A",
    x"3009C32",
    x"3009A0B",
    x"30097E5",
    x"30095C0",
    x"300939A",
    x"3009176",
    x"3008F52",
    x"3008D2E",
    x"3008B0B",
    x"30088E9",
    x"30086C7",
    x"30084A5",
    x"3008284",
    x"3008064",
    x"3007E44",
    x"3007C25",
    x"3007A06",
    x"30077E8",
    x"30075CA",
    x"30073AD",
    x"3007190",
    x"3006F74",
    x"3006D58",
    x"3006B3D",
    x"3006923",
    x"3006709",
    x"30064EF",
    x"30062D6",
    x"30060BE",
    x"3005EA6",
    x"3005C8F",
    x"3005A78",
    x"3005861",
    x"300564C",
    x"3005436",
    x"3005221",
    x"300500D",
    x"3004DF9",
    x"3004BE6",
    x"30049D3",
    x"30047C1",
    x"30045B0",
    x"300439E",
    x"300418E",
    x"3003F7E",
    x"3003D6E",
    x"3003B5F",
    x"3003950",
    x"3003742",
    x"3003535",
    x"3003328",
    x"300311B",
    x"3002F0F",
    x"3002D04",
    x"3002AF9",
    x"30028EE",
    x"30026E4",
    x"30024DB",
    x"30022D2",
    x"30020C9",
    x"3001EC1",
    x"3001CBA",
    x"3001AB3",
    x"30018AD",
    x"30016A7",
    x"30014A1",
    x"300129C",
    x"3001098",
    x"3000E94",
    x"3000C91",
    x"3000A8E",
    x"300088B",
    x"3000689",
    x"3000488",
    x"3000287",
    x"3000087",
    x"2FFFD0E",
    x"2FFF90F",
    x"2FFF512",
    x"2FFF115",
    x"2FFED19",
    x"2FFE91E",
    x"2FFE525",
    x"2FFE12C",
    x"2FFDD34",
    x"2FFD93D",
    x"2FFD547",
    x"2FFD153",
    x"2FFCD5F",
    x"2FFC96C",
    x"2FFC57A",
    x"2FFC189",
    x"2FFBD99",
    x"2FFB9AA",
    x"2FFB5BC",
    x"2FFB1CF",
    x"2FFADE4",
    x"2FFA9F9",
    x"2FFA60F",
    x"2FFA226",
    x"2FF9E3D",
    x"2FF9A56",
    x"2FF9670",
    x"2FF928B",
    x"2FF8EA7",
    x"2FF8AC4",
    x"2FF86E2",
    x"2FF8300",
    x"2FF7F20",
    x"2FF7B41",
    x"2FF7762",
    x"2FF7385",
    x"2FF6FA9",
    x"2FF6BCD",
    x"2FF67F3",
    x"2FF6419",
    x"2FF6041",
    x"2FF5C69",
    x"2FF5893",
    x"2FF54BD",
    x"2FF50E8",
    x"2FF4D14",
    x"2FF4942",
    x"2FF4570",
    x"2FF419F",
    x"2FF3DCF",
    x"2FF3A00",
    x"2FF3632",
    x"2FF3265",
    x"2FF2E99",
    x"2FF2ACE",
    x"2FF2703",
    x"2FF233A",
    x"2FF1F72",
    x"2FF1BAA",
    x"2FF17E4",
    x"2FF141E",
    x"2FF105A",
    x"2FF0C96",
    x"2FF08D4",
    x"2FF0512",
    x"2FF0151",
    x"2FEFD91",
    x"2FEF9D2",
    x"2FEF614",
    x"2FEF257",
    x"2FEEE9B",
    x"2FEEAE0",
    x"2FEE726",
    x"2FEE36C",
    x"2FEDFB4",
    x"2FEDBFD",
    x"2FED846",
    x"2FED490",
    x"2FED0DC",
    x"2FECD28",
    x"2FEC975",
    x"2FEC5C3",
    x"2FEC212",
    x"2FEBE62",
    x"2FEBAB3",
    x"2FEB705",
    x"2FEB358",
    x"2FEAFAB",
    x"2FEAC00",
    x"2FEA855",
    x"2FEA4AC",
    x"2FEA103",
    x"2FE9D5B",
    x"2FE99B4",
    x"2FE960E",
    x"2FE9269",
    x"2FE8EC5",
    x"2FE8B22",
    x"2FE877F",
    x"2FE83DE",
    x"2FE803D",
    x"2FE7C9E",
    x"2FE78FF",
    x"2FE7561",
    x"2FE71C4",
    x"2FE6E28",
    x"2FE6A8D",
    x"2FE66F3",
    x"2FE635A",
    x"2FE5FC2",
    x"2FE5C2A",
    x"2FE5893",
    x"2FE54FE",
    x"2FE5169",
    x"2FE4DD5",
    x"2FE4A42",
    x"2FE46B0",
    x"2FE431F",
    x"2FE3F8E",
    x"2FE3BFF",
    x"2FE3870",
    x"2FE34E3",
    x"2FE3156",
    x"2FE2DCA",
    x"2FE2A3F",
    x"2FE26B5",
    x"2FE232C",
    x"2FE1FA3",
    x"2FE1C1C",
    x"2FE1895",
    x"2FE1510",
    x"2FE118B",
    x"2FE0E07",
    x"2FE0A84",
    x"2FE0702",
    x"2FE0380",
    x"2FE0000",
    x"2FDFC80",
    x"2FDF901",
    x"2FDF584",
    x"2FDF207",
    x"2FDEE8B",
    x"2FDEB0F",
    x"2FDE795",
    x"2FDE41C",
    x"2FDE0A3",
    x"2FDDD2B",
    x"2FDD9B4",
    x"2FDD63F",
    x"2FDD2C9",
    x"2FDCF55",
    x"2FDCBE2",
    x"2FDC86F",
    x"2FDC4FD",
    x"2FDC18D",
    x"2FDBE1D",
    x"2FDBAAE",
    x"2FDB73F",
    x"2FDB3D2",
    x"2FDB065",
    x"2FDACFA",
    x"2FDA98F",
    x"2FDA625",
    x"2FDA2BC",
    x"2FD9F54",
    x"2FD9BEC",
    x"2FD9886",
    x"2FD9520",
    x"2FD91BB",
    x"2FD8E57",
    x"2FD8AF4",
    x"2FD8792",
    x"2FD8430",
    x"2FD80D0",
    x"2FD7D70",
    x"2FD7A11",
    x"2FD76B3",
    x"2FD7355",
    x"2FD6FF9",
    x"2FD6C9D",
    x"2FD6943",
    x"2FD65E9",
    x"2FD6290",
    x"2FD5F38",
    x"2FD5BE0",
    x"2FD588A",
    x"2FD5534",
    x"2FD51DF",
    x"2FD4E8B",
    x"2FD4B38",
    x"2FD47E5",
    x"2FD4494",
    x"2FD4143",
    x"2FD3DF3",
    x"2FD3AA4",
    x"2FD3756",
    x"2FD3408",
    x"2FD30BC",
    x"2FD2D70",
    x"2FD2A25",
    x"2FD26DB",
    x"2FD2392",
    x"2FD2049",
    x"2FD1D02",
    x"2FD19BB",
    x"2FD1675",
    x"2FD132F",
    x"2FD0FEB",
    x"2FD0CA8",
    x"2FD0965",
    x"2FD0623",
    x"2FD02E2",
    x"2FCFFA1",
    x"2FCFC62",
    x"2FCF923",
    x"2FCF5E5",
    x"2FCF2A8",
    x"2FCEF6C",
    x"2FCEC31",
    x"2FCE8F6",
    x"2FCE5BC",
    x"2FCE283",
    x"2FCDF4B",
    x"2FCDC13",
    x"2FCD8DD",
    x"2FCD5A7",
    x"2FCD272",
    x"2FCCF3E",
    x"2FCCC0A",
    x"2FCC8D8",
    x"2FCC5A6",
    x"2FCC275",
    x"2FCBF45",
    x"2FCBC15",
    x"2FCB8E7",
    x"2FCB5B9",
    x"2FCB28C",
    x"2FCAF5F",
    x"2FCAC34",
    x"2FCA909",
    x"2FCA5E0",
    x"2FCA2B6",
    x"2FC9F8E",
    x"2FC9C67",
    x"2FC9940",
    x"2FC961A",
    x"2FC92F5",
    x"2FC8FD1",
    x"2FC8CAD",
    x"2FC898A",
    x"2FC8668",
    x"2FC8347",
    x"2FC8027",
    x"2FC7D07",
    x"2FC79E8",
    x"2FC76CA",
    x"2FC73AD",
    x"2FC7090",
    x"2FC6D74",
    x"2FC6A59",
    x"2FC673F",
    x"2FC6426",
    x"2FC610D",
    x"2FC5DF5",
    x"2FC5ADE",
    x"2FC57C8",
    x"2FC54B2",
    x"2FC519D",
    x"2FC4E89",
    x"2FC4B76",
    x"2FC4864",
    x"2FC4552",
    x"2FC4241",
    x"2FC3F31",
    x"2FC3C21",
    x"2FC3913",
    x"2FC3605",
    x"2FC32F8",
    x"2FC2FEB",
    x"2FC2CE0",
    x"2FC29D5",
    x"2FC26CB",
    x"2FC23C2",
    x"2FC20B9",
    x"2FC1DB1",
    x"2FC1AAA",
    x"2FC17A4",
    x"2FC149E",
    x"2FC119A",
    x"2FC0E96",
    x"2FC0B92",
    x"2FC0890",
    x"2FC058E",
    x"2FC028D",
    x"2FBFF8D",
    x"2FBFC8D",
    x"2FBF98E",
    x"2FBF690",
    x"2FBF393",
    x"2FBF097",
    x"2FBED9B",
    x"2FBEAA0",
    x"2FBE7A6",
    x"2FBE4AC",
    x"2FBE1B3",
    x"2FBDEBB",
    x"2FBDBC4",
    x"2FBD8CD",
    x"2FBD5D7",
    x"2FBD2E2",
    x"2FBCFEE",
    x"2FBCCFA",
    x"2FBCA08",
    x"2FBC715",
    x"2FBC424",
    x"2FBC133",
    x"2FBBE43",
    x"2FBBB54",
    x"2FBB866",
    x"2FBB578",
    x"2FBB28B",
    x"2FBAF9F",
    x"2FBACB3",
    x"2FBA9C8",
    x"2FBA6DE",
    x"2FBA3F5",
    x"2FBA10C",
    x"2FB9E24",
    x"2FB9B3D",
    x"2FB9857",
    x"2FB9571",
    x"2FB928C",
    x"2FB8FA8",
    x"2FB8CC4",
    x"2FB89E1",
    x"2FB86FF",
    x"2FB841E",
    x"2FB813D",
    x"2FB7E5D",
    x"2FB7B7E",
    x"2FB78A0",
    x"2FB75C2",
    x"2FB72E5",
    x"2FB7008",
    x"2FB6D2D",
    x"2FB6A52",
    x"2FB6777",
    x"2FB649E",
    x"2FB61C5",
    x"2FB5EED",
    x"2FB5C16",
    x"2FB593F",
    x"2FB5669",
    x"2FB5394",
    x"2FB50BF",
    x"2FB4DEB",
    x"2FB4B18",
    x"2FB4846",
    x"2FB4574",
    x"2FB42A3",
    x"2FB3FD3",
    x"2FB3D03",
    x"2FB3A34",
    x"2FB3766",
    x"2FB3499",
    x"2FB31CC",
    x"2FB2F00",
    x"2FB2C34",
    x"2FB296A",
    x"2FB26A0",
    x"2FB23D6",
    x"2FB210E",
    x"2FB1E46",
    x"2FB1B7F",
    x"2FB18B8",
    x"2FB15F2",
    x"2FB132D",
    x"2FB1069",
    x"2FB0DA5",
    x"2FB0AE2",
    x"2FB081F",
    x"2FB055E",
    x"2FB029D",
    x"2FAFFDC",
    x"2FAFD1D",
    x"2FAFA5E",
    x"2FAF7A0",
    x"2FAF4E2",
    x"2FAF225",
    x"2FAEF69",
    x"2FAECAE",
    x"2FAE9F3",
    x"2FAE739",
    x"2FAE47F",
    x"2FAE1C6",
    x"2FADF0E",
    x"2FADC57",
    x"2FAD9A0",
    x"2FAD6EA",
    x"2FAD435",
    x"2FAD180",
    x"2FACECC",
    x"2FACC18",
    x"2FAC966",
    x"2FAC6B4",
    x"2FAC402",
    x"2FAC152",
    x"2FABEA2",
    x"2FABBF2",
    x"2FAB944",
    x"2FAB696",
    x"2FAB3E8",
    x"2FAB13C",
    x"2FAAE90",
    x"2FAABE5",
    x"2FAA93A",
    x"2FAA690",
    x"2FAA3E7",
    x"2FAA13E",
    x"2FA9E96",
    x"2FA9BEF",
    x"2FA9948",
    x"2FA96A2",
    x"2FA93FD",
    x"2FA9158",
    x"2FA8EB4",
    x"2FA8C11",
    x"2FA896E",
    x"2FA86CC",
    x"2FA842B",
    x"2FA818A",
    x"2FA7EEA",
    x"2FA7C4A",
    x"2FA79AC",
    x"2FA770E",
    x"2FA7470",
    x"2FA71D3",
    x"2FA6F37",
    x"2FA6C9C",
    x"2FA6A01",
    x"2FA6767",
    x"2FA64CD",
    x"2FA6234",
    x"2FA5F9C",
    x"2FA5D05",
    x"2FA5A6E",
    x"2FA57D7",
    x"2FA5542",
    x"2FA52AD",
    x"2FA5018",
    x"2FA4D85",
    x"2FA4AF2",
    x"2FA485F",
    x"2FA45CD",
    x"2FA433C",
    x"2FA40AC",
    x"2FA3E1C",
    x"2FA3B8D",
    x"2FA38FE",
    x"2FA3670",
    x"2FA33E3",
    x"2FA3156",
    x"2FA2ECA",
    x"2FA2C3F",
    x"2FA29B4",
    x"2FA272A",
    x"2FA24A1",
    x"2FA2218",
    x"2FA1F90",
    x"2FA1D08",
    x"2FA1A81",
    x"2FA17FB",
    x"2FA1575",
    x"2FA12F0",
    x"2FA106C",
    x"2FA0DE8",
    x"2FA0B65",
    x"2FA08E2",
    x"2FA0660",
    x"2FA03DF",
    x"2FA015E",
    x"2F9FEDE",
    x"2F9FC5F",
    x"2F9F9E0",
    x"2F9F762",
    x"2F9F4E4",
    x"2F9F267",
    x"2F9EFEB",
    x"2F9ED6F",
    x"2F9EAF4",
    x"2F9E87A",
    x"2F9E600",
    x"2F9E387",
    x"2F9E10E",
    x"2F9DE96",
    x"2F9DC1F",
    x"2F9D9A8",
    x"2F9D732",
    x"2F9D4BD",
    x"2F9D248",
    x"2F9CFD4",
    x"2F9CD60",
    x"2F9CAED",
    x"2F9C87B",
    x"2F9C609",
    x"2F9C398",
    x"2F9C127",
    x"2F9BEB7",
    x"2F9BC48",
    x"2F9B9D9",
    x"2F9B76B",
    x"2F9B4FD",
    x"2F9B290",
    x"2F9B024",
    x"2F9ADB8",
    x"2F9AB4D",
    x"2F9A8E2",
    x"2F9A678",
    x"2F9A40F",
    x"2F9A1A6",
    x"2F99F3E",
    x"2F99CD7",
    x"2F99A70",
    x"2F9980A",
    x"2F995A4",
    x"2F9933F",
    x"2F990DA",
    x"2F98E76",
    x"2F98C13",
    x"2F989B0",
    x"2F9874E",
    x"2F984ED",
    x"2F9828C",
    x"2F9802B",
    x"2F97DCC",
    x"2F97B6D",
    x"2F9790E",
    x"2F976B0",
    x"2F97453",
    x"2F971F6",
    x"2F96F9A",
    x"2F96D3E",
    x"2F96AE3",
    x"2F96889",
    x"2F9662F",
    x"2F963D5",
    x"2F9617D",
    x"2F95F25",
    x"2F95CCD",
    x"2F95A76",
    x"2F95820",
    x"2F955CA",
    x"2F95375",
    x"2F95121",
    x"2F94ECD",
    x"2F94C79",
    x"2F94A26",
    x"2F947D4",
    x"2F94582",
    x"2F94331",
    x"2F940E1",
    x"2F93E91",
    x"2F93C42",
    x"2F939F3",
    x"2F937A5",
    x"2F93557",
    x"2F9330A",
    x"2F930BD",
    x"2F92E71",
    x"2F92C26",
    x"2F929DB",
    x"2F92791",
    x"2F92548",
    x"2F922FF",
    x"2F920B6",
    x"2F91E6E",
    x"2F91C27",
    x"2F919E0",
    x"2F9179A",
    x"2F91554",
    x"2F9130F",
    x"2F910CB",
    x"2F90E87",
    x"2F90C44",
    x"2F90A01",
    x"2F907BF",
    x"2F9057D",
    x"2F9033C",
    x"2F900FB",
    x"2F8FEBB",
    x"2F8FC7C",
    x"2F8FA3D",
    x"2F8F7FF",
    x"2F8F5C1",
    x"2F8F384",
    x"2F8F147",
    x"2F8EF0B",
    x"2F8ECD0",
    x"2F8EA95",
    x"2F8E85B",
    x"2F8E621",
    x"2F8E3E7",
    x"2F8E1AF",
    x"2F8DF77",
    x"2F8DD3F",
    x"2F8DB08",
    x"2F8D8D1",
    x"2F8D69C",
    x"2F8D466",
    x"2F8D231",
    x"2F8CFFD",
    x"2F8CDC9",
    x"2F8CB96",
    x"2F8C964",
    x"2F8C732",
    x"2F8C500",
    x"2F8C2CF",
    x"2F8C09F",
    x"2F8BE6F",
    x"2F8BC3F",
    x"2F8BA11",
    x"2F8B7E2",
    x"2F8B5B5",
    x"2F8B387",
    x"2F8B15B",
    x"2F8AF2F",
    x"2F8AD03",
    x"2F8AAD8",
    x"2F8A8AE",
    x"2F8A684",
    x"2F8A45B",
    x"2F8A232",
    x"2F8A009",
    x"2F89DE2",
    x"2F89BBB",
    x"2F89994",
    x"2F8976E",
    x"2F89548",
    x"2F89323",
    x"2F890FF",
    x"2F88EDB",
    x"2F88CB7",
    x"2F88A94",
    x"2F88872",
    x"2F88650",
    x"2F8842F",
    x"2F8820E",
    x"2F87FEE",
    x"2F87DCE",
    x"2F87BAF",
    x"2F87990",
    x"2F87772",
    x"2F87554",
    x"2F87337",
    x"2F8711B",
    x"2F86EFF",
    x"2F86CE3",
    x"2F86AC8",
    x"2F868AE",
    x"2F86694",
    x"2F8647B",
    x"2F86262",
    x"2F86049",
    x"2F85E32",
    x"2F85C1A",
    x"2F85A04",
    x"2F857ED",
    x"2F855D8",
    x"2F853C2",
    x"2F851AE",
    x"2F84F9A",
    x"2F84D86",
    x"2F84B73",
    x"2F84960",
    x"2F8474E",
    x"2F8453D",
    x"2F8432B",
    x"2F8411B",
    x"2F83F0B",
    x"2F83CFB",
    x"2F83AEC",
    x"2F838DE",
    x"2F836D0",
    x"2F834C3",
    x"2F832B6",
    x"2F830A9",
    x"2F82E9D",
    x"2F82C92",
    x"2F82A87",
    x"2F8287D",
    x"2F82673",
    x"2F82469",
    x"2F82261",
    x"2F82058",
    x"2F81E50",
    x"2F81C49",
    x"2F81A42",
    x"2F8183C",
    x"2F81636",
    x"2F81431",
    x"2F8122C",
    x"2F81028",
    x"2F80E24",
    x"2F80C21",
    x"2F80A1E",
    x"2F8081C",
    x"2F8061A",
    x"2F80419",
    x"2F80218",
    x"2F80017",
    x"2F7FC30",
    x"2F7F831",
    x"2F7F434",
    x"2F7F037",
    x"2F7EC3C",
    x"2F7E841",
    x"2F7E448",
    x"2F7E04F",
    x"2F7DC57",
    x"2F7D861",
    x"2F7D46B",
    x"2F7D077",
    x"2F7CC83",
    x"2F7C890",
    x"2F7C49F",
    x"2F7C0AE",
    x"2F7BCBE",
    x"2F7B8D0",
    x"2F7B4E2",
    x"2F7B0F5",
    x"2F7AD09",
    x"2F7A91F",
    x"2F7A535",
    x"2F7A14C",
    x"2F79D64",
    x"2F7997D",
    x"2F79598",
    x"2F791B3",
    x"2F78DCF",
    x"2F789EC",
    x"2F7860A",
    x"2F78229",
    x"2F77E49",
    x"2F77A6A",
    x"2F7768B",
    x"2F772AE",
    x"2F76ED2",
    x"2F76AF7",
    x"2F7671D",
    x"2F76343",
    x"2F75F6B",
    x"2F75B94",
    x"2F757BD",
    x"2F753E8",
    x"2F75013",
    x"2F74C40",
    x"2F7486D",
    x"2F7449B",
    x"2F740CB",
    x"2F73CFB",
    x"2F7392C",
    x"2F7355E",
    x"2F73192",
    x"2F72DC6",
    x"2F729FB",
    x"2F72631",
    x"2F72268",
    x"2F71EA0",
    x"2F71AD8",
    x"2F71712",
    x"2F7134D",
    x"2F70F88",
    x"2F70BC5",
    x"2F70803",
    x"2F70441",
    x"2F70080",
    x"2F6FCC1",
    x"2F6F902",
    x"2F6F544",
    x"2F6F187",
    x"2F6EDCB",
    x"2F6EA11",
    x"2F6E656",
    x"2F6E29D",
    x"2F6DEE5",
    x"2F6DB2E",
    x"2F6D778",
    x"2F6D3C2",
    x"2F6D00E",
    x"2F6CC5A",
    x"2F6C8A8",
    x"2F6C4F6",
    x"2F6C145",
    x"2F6BD95",
    x"2F6B9E6",
    x"2F6B638",
    x"2F6B28B",
    x"2F6AEDF",
    x"2F6AB34",
    x"2F6A789",
    x"2F6A3E0",
    x"2F6A037",
    x"2F69C90",
    x"2F698E9",
    x"2F69543",
    x"2F6919E",
    x"2F68DFB",
    x"2F68A58",
    x"2F686B5",
    x"2F68314",
    x"2F67F74",
    x"2F67BD4",
    x"2F67836",
    x"2F67498",
    x"2F670FC",
    x"2F66D60",
    x"2F669C5",
    x"2F6662B",
    x"2F66292",
    x"2F65EFA",
    x"2F65B62",
    x"2F657CC",
    x"2F65436",
    x"2F650A2",
    x"2F64D0E",
    x"2F6497B",
    x"2F645E9",
    x"2F64258",
    x"2F63EC8",
    x"2F63B39",
    x"2F637AB",
    x"2F6341D",
    x"2F63091",
    x"2F62D05",
    x"2F6297A",
    x"2F625F0",
    x"2F62267",
    x"2F61EDF",
    x"2F61B58",
    x"2F617D1",
    x"2F6144C",
    x"2F610C7",
    x"2F60D43",
    x"2F609C0",
    x"2F6063E",
    x"2F602BD",
    x"2F5FF3D",
    x"2F5FBBE",
    x"2F5F83F",
    x"2F5F4C2",
    x"2F5F145",
    x"2F5EDC9",
    x"2F5EA4E",
    x"2F5E6D4",
    x"2F5E35B",
    x"2F5DFE2",
    x"2F5DC6B",
    x"2F5D8F4",
    x"2F5D57E",
    x"2F5D209",
    x"2F5CE95",
    x"2F5CB22",
    x"2F5C7B0",
    x"2F5C43E",
    x"2F5C0CD",
    x"2F5BD5E",
    x"2F5B9EF",
    x"2F5B681",
    x"2F5B313",
    x"2F5AFA7",
    x"2F5AC3C",
    x"2F5A8D1",
    x"2F5A567",
    x"2F5A1FE",
    x"2F59E96",
    x"2F59B2F",
    x"2F597C9",
    x"2F59463",
    x"2F590FE",
    x"2F58D9B",
    x"2F58A38",
    x"2F586D5",
    x"2F58374",
    x"2F58014",
    x"2F57CB4",
    x"2F57955",
    x"2F575F8",
    x"2F5729A",
    x"2F56F3E",
    x"2F56BE3",
    x"2F56888",
    x"2F5652F",
    x"2F561D6",
    x"2F55E7E",
    x"2F55B26",
    x"2F557D0",
    x"2F5547B",
    x"2F55126",
    x"2F54DD2",
    x"2F54A7F",
    x"2F5472D",
    x"2F543DB",
    x"2F5408B",
    x"2F53D3B",
    x"2F539EC",
    x"2F5369E",
    x"2F53351",
    x"2F53004",
    x"2F52CB9",
    x"2F5296E",
    x"2F52624",
    x"2F522DB",
    x"2F51F93",
    x"2F51C4B",
    x"2F51905",
    x"2F515BF",
    x"2F5127A",
    x"2F50F35",
    x"2F50BF2",
    x"2F508AF",
    x"2F5056E",
    x"2F5022D",
    x"2F4FEED",
    x"2F4FBAD",
    x"2F4F86F",
    x"2F4F531",
    x"2F4F1F4",
    x"2F4EEB8",
    x"2F4EB7D",
    x"2F4E842",
    x"2F4E509",
    x"2F4E1D0",
    x"2F4DE98",
    x"2F4DB61",
    x"2F4D82A",
    x"2F4D4F4",
    x"2F4D1C0",
    x"2F4CE8C",
    x"2F4CB58",
    x"2F4C826",
    x"2F4C4F4",
    x"2F4C1C3",
    x"2F4BE93",
    x"2F4BB64",
    x"2F4B836",
    x"2F4B508",
    x"2F4B1DB",
    x"2F4AEAF",
    x"2F4AB84",
    x"2F4A859",
    x"2F4A530",
    x"2F4A207",
    x"2F49EDF",
    x"2F49BB7",
    x"2F49891",
    x"2F4956B",
    x"2F49246",
    x"2F48F22",
    x"2F48BFE",
    x"2F488DC",
    x"2F485BA",
    x"2F48299",
    x"2F47F79",
    x"2F47C59",
    x"2F4793B",
    x"2F4761D",
    x"2F47300",
    x"2F46FE3",
    x"2F46CC8",
    x"2F469AD",
    x"2F46693",
    x"2F46379",
    x"2F46061",
    x"2F45D49",
    x"2F45A32",
    x"2F4571C",
    x"2F45407",
    x"2F450F2",
    x"2F44DDE",
    x"2F44ACB",
    x"2F447B9",
    x"2F444A7",
    x"2F44197",
    x"2F43E87",
    x"2F43B77",
    x"2F43869",
    x"2F4355B",
    x"2F4324E",
    x"2F42F42",
    x"2F42C37",
    x"2F4292C",
    x"2F42622",
    x"2F42319",
    x"2F42010",
    x"2F41D09",
    x"2F41A02",
    x"2F416FC",
    x"2F413F6",
    x"2F410F2",
    x"2F40DEE",
    x"2F40AEB",
    x"2F407E8",
    x"2F404E7",
    x"2F401E6",
    x"2F3FEE6",
    x"2F3FBE7",
    x"2F3F8E8",
    x"2F3F5EA",
    x"2F3F2ED",
    x"2F3EFF1",
    x"2F3ECF5",
    x"2F3E9FA",
    x"2F3E700",
    x"2F3E407",
    x"2F3E10E",
    x"2F3DE16",
    x"2F3DB1F",
    x"2F3D829",
    x"2F3D533",
    x"2F3D23E",
    x"2F3CF4A",
    x"2F3CC56",
    x"2F3C964",
    x"2F3C672",
    x"2F3C380",
    x"2F3C090",
    x"2F3BDA0",
    x"2F3BAB1",
    x"2F3B7C3",
    x"2F3B4D5",
    x"2F3B1E8",
    x"2F3AEFC",
    x"2F3AC11",
    x"2F3A926",
    x"2F3A63C",
    x"2F3A353",
    x"2F3A06B",
    x"2F39D83",
    x"2F39A9C",
    x"2F397B6",
    x"2F394D0",
    x"2F391EB",
    x"2F38F07",
    x"2F38C24",
    x"2F38941",
    x"2F3865F",
    x"2F3837E",
    x"2F3809D",
    x"2F37DBD",
    x"2F37ADE",
    x"2F37800",
    x"2F37522",
    x"2F37245",
    x"2F36F69",
    x"2F36C8E",
    x"2F369B3",
    x"2F366D9",
    x"2F36400",
    x"2F36127",
    x"2F35E4F",
    x"2F35B78",
    x"2F358A1",
    x"2F355CB",
    x"2F352F6",
    x"2F35022",
    x"2F34D4E",
    x"2F34A7B",
    x"2F347A9",
    x"2F344D7",
    x"2F34207",
    x"2F33F36",
    x"2F33C67",
    x"2F33998",
    x"2F336CA",
    x"2F333FD",
    x"2F33130",
    x"2F32E64",
    x"2F32B99",
    x"2F328CE",
    x"2F32605",
    x"2F3233B",
    x"2F32073",
    x"2F31DAB",
    x"2F31AE4",
    x"2F3181E",
    x"2F31558",
    x"2F31293",
    x"2F30FCF",
    x"2F30D0B",
    x"2F30A48",
    x"2F30786",
    x"2F304C5",
    x"2F30204",
    x"2F2FF44",
    x"2F2FC84",
    x"2F2F9C5",
    x"2F2F707",
    x"2F2F44A",
    x"2F2F18D",
    x"2F2EED1",
    x"2F2EC16",
    x"2F2E95B",
    x"2F2E6A1",
    x"2F2E3E8",
    x"2F2E12F",
    x"2F2DE77",
    x"2F2DBC0",
    x"2F2D909",
    x"2F2D653",
    x"2F2D39E",
    x"2F2D0E9",
    x"2F2CE36",
    x"2F2CB82",
    x"2F2C8D0",
    x"2F2C61E",
    x"2F2C36D",
    x"2F2C0BC",
    x"2F2BE0C",
    x"2F2BB5D",
    x"2F2B8AF",
    x"2F2B601",
    x"2F2B354",
    x"2F2B0A7",
    x"2F2ADFB",
    x"2F2AB50",
    x"2F2A8A6",
    x"2F2A5FC",
    x"2F2A353",
    x"2F2A0AA",
    x"2F29E02",
    x"2F29B5B",
    x"2F298B5",
    x"2F2960F",
    x"2F2936A",
    x"2F290C5",
    x"2F28E21",
    x"2F28B7E",
    x"2F288DB",
    x"2F2863A",
    x"2F28398",
    x"2F280F8",
    x"2F27E58",
    x"2F27BB9",
    x"2F2791A",
    x"2F2767C",
    x"2F273DF",
    x"2F27142",
    x"2F26EA6",
    x"2F26C0B",
    x"2F26970",
    x"2F266D6",
    x"2F2643D",
    x"2F261A4",
    x"2F25F0C",
    x"2F25C74",
    x"2F259DE",
    x"2F25748",
    x"2F254B2",
    x"2F2521D",
    x"2F24F89",
    x"2F24CF5",
    x"2F24A62",
    x"2F247D0",
    x"2F2453F",
    x"2F242AE",
    x"2F2401D",
    x"2F23D8E",
    x"2F23AFE",
    x"2F23870",
    x"2F235E2",
    x"2F23355",
    x"2F230C9",
    x"2F22E3D",
    x"2F22BB1",
    x"2F22927",
    x"2F2269D",
    x"2F22414",
    x"2F2218B",
    x"2F21F03",
    x"2F21C7B",
    x"2F219F5",
    x"2F2176E",
    x"2F214E9",
    x"2F21264",
    x"2F20FE0",
    x"2F20D5C",
    x"2F20AD9",
    x"2F20857",
    x"2F205D5",
    x"2F20354",
    x"2F200D3",
    x"2F1FE53",
    x"2F1FBD4",
    x"2F1F955",
    x"2F1F6D7",
    x"2F1F45A",
    x"2F1F1DD",
    x"2F1EF61",
    x"2F1ECE5",
    x"2F1EA6A",
    x"2F1E7F0",
    x"2F1E577",
    x"2F1E2FD",
    x"2F1E085",
    x"2F1DE0D",
    x"2F1DB96",
    x"2F1D91F",
    x"2F1D6A9",
    x"2F1D434",
    x"2F1D1BF",
    x"2F1CF4B",
    x"2F1CCD8",
    x"2F1CA65",
    x"2F1C7F2",
    x"2F1C581",
    x"2F1C310",
    x"2F1C09F",
    x"2F1BE2F",
    x"2F1BBC0",
    x"2F1B952",
    x"2F1B6E4",
    x"2F1B476",
    x"2F1B209",
    x"2F1AF9D",
    x"2F1AD31",
    x"2F1AAC6",
    x"2F1A85C",
    x"2F1A5F2",
    x"2F1A389",
    x"2F1A121",
    x"2F19EB9",
    x"2F19C51",
    x"2F199EA",
    x"2F19784",
    x"2F1951F",
    x"2F192BA",
    x"2F19055",
    x"2F18DF1",
    x"2F18B8E",
    x"2F1892C",
    x"2F186CA",
    x"2F18468",
    x"2F18208",
    x"2F17FA7",
    x"2F17D48",
    x"2F17AE9",
    x"2F1788A",
    x"2F1762C",
    x"2F173CF",
    x"2F17172",
    x"2F16F16",
    x"2F16CBB",
    x"2F16A60",
    x"2F16806",
    x"2F165AC",
    x"2F16353",
    x"2F160FA",
    x"2F15EA2",
    x"2F15C4B",
    x"2F159F4",
    x"2F1579E",
    x"2F15548",
    x"2F152F3",
    x"2F1509F",
    x"2F14E4B",
    x"2F14BF8",
    x"2F149A5",
    x"2F14753",
    x"2F14501",
    x"2F142B1",
    x"2F14060",
    x"2F13E10",
    x"2F13BC1",
    x"2F13972",
    x"2F13724",
    x"2F134D7",
    x"2F1328A",
    x"2F1303E",
    x"2F12DF2",
    x"2F12BA7",
    x"2F1295C",
    x"2F12712",
    x"2F124C8",
    x"2F12280",
    x"2F12037",
    x"2F11DEF",
    x"2F11BA8",
    x"2F11962",
    x"2F1171C",
    x"2F114D6",
    x"2F11291",
    x"2F1104D",
    x"2F10E09",
    x"2F10BC6",
    x"2F10983",
    x"2F10741",
    x"2F104FF",
    x"2F102BE",
    x"2F1007E",
    x"2F0FE3E",
    x"2F0FBFF",
    x"2F0F9C0",
    x"2F0F782",
    x"2F0F544",
    x"2F0F307",
    x"2F0F0CB",
    x"2F0EE8F",
    x"2F0EC54",
    x"2F0EA19",
    x"2F0E7DF",
    x"2F0E5A5",
    x"2F0E36C",
    x"2F0E133",
    x"2F0DEFB",
    x"2F0DCC4",
    x"2F0DA8D",
    x"2F0D856",
    x"2F0D621",
    x"2F0D3EB",
    x"2F0D1B7",
    x"2F0CF83",
    x"2F0CD4F",
    x"2F0CB1C",
    x"2F0C8E9",
    x"2F0C6B7",
    x"2F0C486",
    x"2F0C255",
    x"2F0C025",
    x"2F0BDF5",
    x"2F0BBC6",
    x"2F0B997",
    x"2F0B769",
    x"2F0B53C",
    x"2F0B30E",
    x"2F0B0E2",
    x"2F0AEB6",
    x"2F0AC8B",
    x"2F0AA60",
    x"2F0A835",
    x"2F0A60C",
    x"2F0A3E2",
    x"2F0A1BA",
    x"2F09F92",
    x"2F09D6A",
    x"2F09B43",
    x"2F0991C",
    x"2F096F6",
    x"2F094D1",
    x"2F092AC",
    x"2F09087",
    x"2F08E64",
    x"2F08C40",
    x"2F08A1D",
    x"2F087FB",
    x"2F085D9",
    x"2F083B8",
    x"2F08198",
    x"2F07F78",
    x"2F07D58",
    x"2F07B39",
    x"2F0791A",
    x"2F076FC",
    x"2F074DF",
    x"2F072C2",
    x"2F070A5",
    x"2F06E8A",
    x"2F06C6E",
    x"2F06A53",
    x"2F06839",
    x"2F0661F",
    x"2F06406",
    x"2F061ED",
    x"2F05FD5",
    x"2F05DBD",
    x"2F05BA6",
    x"2F0598F",
    x"2F05779",
    x"2F05564",
    x"2F0534F",
    x"2F0513A",
    x"2F04F26",
    x"2F04D12",
    x"2F04AFF",
    x"2F048ED",
    x"2F046DB",
    x"2F044CA",
    x"2F042B9",
    x"2F040A8",
    x"2F03E98",
    x"2F03C89",
    x"2F03A7A",
    x"2F0386C",
    x"2F0365E",
    x"2F03450",
    x"2F03244",
    x"2F03037",
    x"2F02E2C",
    x"2F02C20",
    x"2F02A15",
    x"2F0280B",
    x"2F02601",
    x"2F023F8",
    x"2F021EF",
    x"2F01FE7",
    x"2F01DDF",
    x"2F01BD8",
    x"2F019D2",
    x"2F017CB",
    x"2F015C6",
    x"2F013C0",
    x"2F011BC",
    x"2F00FB8",
    x"2F00DB4",
    x"2F00BB1",
    x"2F009AE",
    x"2F007AC",
    x"2F005AA",
    x"2F003A9",
    x"2F001A8",
    x"2EFFF51",
    x"2EFFB52",
    x"2EFF753",
    x"2EFF356",
    x"2EFEF5A",
    x"2EFEB5E",
    x"2EFE764",
    x"2EFE36B",
    x"2EFDF72",
    x"2EFDB7B",
    x"2EFD785",
    x"2EFD38F",
    x"2EFCF9B",
    x"2EFCBA7",
    x"2EFC7B5",
    x"2EFC3C3",
    x"2EFBFD3",
    x"2EFBBE4",
    x"2EFB7F5",
    x"2EFB408",
    x"2EFB01B",
    x"2EFAC30",
    x"2EFA845",
    x"2EFA45B",
    x"2EFA073",
    x"2EF9C8B",
    x"2EF98A5",
    x"2EF94BF",
    x"2EF90DA",
    x"2EF8CF6",
    x"2EF8914",
    x"2EF8532",
    x"2EF8151",
    x"2EF7D71",
    x"2EF7992",
    x"2EF75B4",
    x"2EF71D7",
    x"2EF6DFC",
    x"2EF6A20",
    x"2EF6646",
    x"2EF626D",
    x"2EF5E95",
    x"2EF5ABE",
    x"2EF56E8",
    x"2EF5313",
    x"2EF4F3E",
    x"2EF4B6B",
    x"2EF4799",
    x"2EF43C7",
    x"2EF3FF7",
    x"2EF3C27",
    x"2EF3859",
    x"2EF348B",
    x"2EF30BE",
    x"2EF2CF3",
    x"2EF2928",
    x"2EF255E",
    x"2EF2195",
    x"2EF1DCD",
    x"2EF1A06",
    x"2EF1640",
    x"2EF127B",
    x"2EF0EB7",
    x"2EF0AF4",
    x"2EF0732",
    x"2EF0370",
    x"2EEFFB0",
    x"2EEFBF0",
    x"2EEF832",
    x"2EEF474",
    x"2EEF0B8",
    x"2EEECFC",
    x"2EEE941",
    x"2EEE587",
    x"2EEE1CE",
    x"2EEDE16",
    x"2EEDA5F",
    x"2EED6A9",
    x"2EED2F4",
    x"2EECF40",
    x"2EECB8C",
    x"2EEC7DA",
    x"2EEC428",
    x"2EEC078",
    x"2EEBCC8",
    x"2EEB919",
    x"2EEB56C",
    x"2EEB1BF",
    x"2EEAE13",
    x"2EEAA68",
    x"2EEA6BE",
    x"2EEA314",
    x"2EE9F6C",
    x"2EE9BC5",
    x"2EE981E",
    x"2EE9479",
    x"2EE90D4",
    x"2EE8D30",
    x"2EE898D",
    x"2EE85EB",
    x"2EE824A",
    x"2EE7EAA",
    x"2EE7B0B",
    x"2EE776D",
    x"2EE73CF",
    x"2EE7033",
    x"2EE6C97",
    x"2EE68FD",
    x"2EE6563",
    x"2EE61CA",
    x"2EE5E32",
    x"2EE5A9B",
    x"2EE5705",
    x"2EE536F",
    x"2EE4FDB",
    x"2EE4C47",
    x"2EE48B5",
    x"2EE4523",
    x"2EE4192",
    x"2EE3E02",
    x"2EE3A73",
    x"2EE36E5",
    x"2EE3358",
    x"2EE2FCB",
    x"2EE2C40",
    x"2EE28B5",
    x"2EE252B",
    x"2EE21A3",
    x"2EE1E1B",
    x"2EE1A93",
    x"2EE170D",
    x"2EE1388",
    x"2EE1004",
    x"2EE0C80",
    x"2EE08FD",
    x"2EE057B",
    x"2EE01FB",
    x"2EDFE7A",
    x"2EDFAFB",
    x"2EDF77D",
    x"2EDF400",
    x"2EDF083",
    x"2EDED07",
    x"2EDE98C",
    x"2EDE612",
    x"2EDE299",
    x"2EDDF21",
    x"2EDDBAA",
    x"2EDD833",
    x"2EDD4BE",
    x"2EDD149",
    x"2EDCDD5",
    x"2EDCA62",
    x"2EDC6F0",
    x"2EDC37F",
    x"2EDC00E",
    x"2EDBC9F",
    x"2EDB930",
    x"2EDB5C2",
    x"2EDB255",
    x"2EDAEE9",
    x"2EDAB7E",
    x"2EDA813",
    x"2EDA4A9",
    x"2EDA141",
    x"2ED9DD9",
    x"2ED9A72",
    x"2ED970C",
    x"2ED93A6",
    x"2ED9042",
    x"2ED8CDE",
    x"2ED897B",
    x"2ED8619",
    x"2ED82B8",
    x"2ED7F58",
    x"2ED7BF9",
    x"2ED789A",
    x"2ED753C",
    x"2ED71DF",
    x"2ED6E83",
    x"2ED6B28",
    x"2ED67CE",
    x"2ED6474",
    x"2ED611C",
    x"2ED5DC4",
    x"2ED5A6D",
    x"2ED5717",
    x"2ED53C1",
    x"2ED506D",
    x"2ED4D19",
    x"2ED49C6",
    x"2ED4674",
    x"2ED4323",
    x"2ED3FD2",
    x"2ED3C83",
    x"2ED3934",
    x"2ED35E6",
    x"2ED3299",
    x"2ED2F4D",
    x"2ED2C02",
    x"2ED28B7",
    x"2ED256D",
    x"2ED2224",
    x"2ED1EDC",
    x"2ED1B95",
    x"2ED184E",
    x"2ED1509",
    x"2ED11C4",
    x"2ED0E80",
    x"2ED0B3D",
    x"2ED07FA",
    x"2ED04B9",
    x"2ED0178",
    x"2ECFE38",
    x"2ECFAF9",
    x"2ECF7BA",
    x"2ECF47D",
    x"2ECF140",
    x"2ECEE04",
    x"2ECEAC9",
    x"2ECE78F",
    x"2ECE455",
    x"2ECE11D",
    x"2ECDDE5",
    x"2ECDAAE",
    x"2ECD777",
    x"2ECD442",
    x"2ECD10D",
    x"2ECCDD9",
    x"2ECCAA6",
    x"2ECC774",
    x"2ECC443",
    x"2ECC112",
    x"2ECBDE2",
    x"2ECBAB3",
    x"2ECB785",
    x"2ECB457",
    x"2ECB12B",
    x"2ECADFF",
    x"2ECAAD4",
    x"2ECA7A9",
    x"2ECA480",
    x"2ECA157",
    x"2EC9E2F",
    x"2EC9B08",
    x"2EC97E2",
    x"2EC94BC",
    x"2EC9197",
    x"2EC8E73",
    x"2EC8B50",
    x"2EC882E",
    x"2EC850C",
    x"2EC81EB",
    x"2EC7ECB",
    x"2EC7BAC",
    x"2EC788D",
    x"2EC756F",
    x"2EC7252",
    x"2EC6F36",
    x"2EC6C1B",
    x"2EC6900",
    x"2EC65E6",
    x"2EC62CD",
    x"2EC5FB5",
    x"2EC5C9D",
    x"2EC5987",
    x"2EC5671",
    x"2EC535B",
    x"2EC5047",
    x"2EC4D33",
    x"2EC4A20",
    x"2EC470E",
    x"2EC43FD",
    x"2EC40EC",
    x"2EC3DDC",
    x"2EC3ACD",
    x"2EC37BF",
    x"2EC34B1",
    x"2EC31A5",
    x"2EC2E99",
    x"2EC2B8D",
    x"2EC2883",
    x"2EC2579",
    x"2EC2270",
    x"2EC1F68",
    x"2EC1C60",
    x"2EC195A",
    x"2EC1654",
    x"2EC134E",
    x"2EC104A",
    x"2EC0D46",
    x"2EC0A43",
    x"2EC0741",
    x"2EC0440",
    x"2EC013F",
    x"2EBFE3F",
    x"2EBFB40",
    x"2EBF841",
    x"2EBF544",
    x"2EBF247",
    x"2EBEF4B",
    x"2EBEC4F",
    x"2EBE955",
    x"2EBE65B",
    x"2EBE361",
    x"2EBE069",
    x"2EBDD71",
    x"2EBDA7A",
    x"2EBD784",
    x"2EBD48E",
    x"2EBD19A",
    x"2EBCEA6",
    x"2EBCBB2",
    x"2EBC8C0",
    x"2EBC5CE",
    x"2EBC2DD",
    x"2EBBFEC",
    x"2EBBCFD",
    x"2EBBA0E",
    x"2EBB720",
    x"2EBB432",
    x"2EBB146",
    x"2EBAE5A",
    x"2EBAB6F",
    x"2EBA884",
    x"2EBA59A",
    x"2EBA2B1",
    x"2EB9FC9",
    x"2EB9CE1",
    x"2EB99FB",
    x"2EB9714",
    x"2EB942F",
    x"2EB914A",
    x"2EB8E66",
    x"2EB8B83",
    x"2EB88A1",
    x"2EB85BF",
    x"2EB82DE",
    x"2EB7FFD",
    x"2EB7D1E",
    x"2EB7A3F",
    x"2EB7761",
    x"2EB7483",
    x"2EB71A6",
    x"2EB6ECA",
    x"2EB6BEF",
    x"2EB6914",
    x"2EB663A",
    x"2EB6361",
    x"2EB6089",
    x"2EB5DB1",
    x"2EB5ADA",
    x"2EB5803",
    x"2EB552E",
    x"2EB5259",
    x"2EB4F85",
    x"2EB4CB1",
    x"2EB49DE",
    x"2EB470C",
    x"2EB443B",
    x"2EB416A",
    x"2EB3E9A",
    x"2EB3BCB",
    x"2EB38FC",
    x"2EB362E",
    x"2EB3361",
    x"2EB3095",
    x"2EB2DC9",
    x"2EB2AFE",
    x"2EB2833",
    x"2EB256A",
    x"2EB22A1",
    x"2EB1FD8",
    x"2EB1D11",
    x"2EB1A4A",
    x"2EB1784",
    x"2EB14BE",
    x"2EB11F9",
    x"2EB0F35",
    x"2EB0C72",
    x"2EB09AF",
    x"2EB06ED",
    x"2EB042B",
    x"2EB016B",
    x"2EAFEAB",
    x"2EAFBEB",
    x"2EAF92D",
    x"2EAF66F",
    x"2EAF3B1",
    x"2EAF0F5",
    x"2EAEE39",
    x"2EAEB7E",
    x"2EAE8C3",
    x"2EAE609",
    x"2EAE350",
    x"2EAE098",
    x"2EADDE0",
    x"2EADB29",
    x"2EAD872",
    x"2EAD5BD",
    x"2EAD307",
    x"2EAD053",
    x"2EACD9F",
    x"2EACAEC",
    x"2EAC83A",
    x"2EAC588",
    x"2EAC2D7",
    x"2EAC027",
    x"2EABD77",
    x"2EABAC8",
    x"2EAB81A",
    x"2EAB56C",
    x"2EAB2BF",
    x"2EAB013",
    x"2EAAD67",
    x"2EAAABC",
    x"2EAA811",
    x"2EAA568",
    x"2EAA2BF",
    x"2EAA016",
    x"2EA9D6F",
    x"2EA9AC8",
    x"2EA9821",
    x"2EA957C",
    x"2EA92D7",
    x"2EA9032",
    x"2EA8D8E",
    x"2EA8AEB",
    x"2EA8849",
    x"2EA85A7",
    x"2EA8306",
    x"2EA8066",
    x"2EA7DC6",
    x"2EA7B27",
    x"2EA7888",
    x"2EA75EB",
    x"2EA734D",
    x"2EA70B1",
    x"2EA6E15",
    x"2EA6B7A",
    x"2EA68DF",
    x"2EA6645",
    x"2EA63AC",
    x"2EA6114",
    x"2EA5E7C",
    x"2EA5BE4",
    x"2EA594E",
    x"2EA56B8",
    x"2EA5422",
    x"2EA518E",
    x"2EA4EFA",
    x"2EA4C66",
    x"2EA49D3",
    x"2EA4741",
    x"2EA44B0",
    x"2EA421F",
    x"2EA3F8F",
    x"2EA3CFF",
    x"2EA3A70",
    x"2EA37E2",
    x"2EA3554",
    x"2EA32C7",
    x"2EA303B",
    x"2EA2DAF",
    x"2EA2B24",
    x"2EA289A",
    x"2EA2610",
    x"2EA2387",
    x"2EA20FE",
    x"2EA1E76",
    x"2EA1BEF",
    x"2EA1968",
    x"2EA16E2",
    x"2EA145D",
    x"2EA11D8",
    x"2EA0F54",
    x"2EA0CD0",
    x"2EA0A4D",
    x"2EA07CB",
    x"2EA0549",
    x"2EA02C8",
    x"2EA0048",
    x"2E9FDC8",
    x"2E9FB49",
    x"2E9F8CB",
    x"2E9F64D",
    x"2E9F3CF",
    x"2E9F153",
    x"2E9EED7",
    x"2E9EC5B",
    x"2E9E9E1",
    x"2E9E766",
    x"2E9E4ED",
    x"2E9E274",
    x"2E9DFFC",
    x"2E9DD84",
    x"2E9DB0D",
    x"2E9D896",
    x"2E9D621",
    x"2E9D3AB",
    x"2E9D137",
    x"2E9CEC3",
    x"2E9CC4F",
    x"2E9C9DD",
    x"2E9C76A",
    x"2E9C4F9",
    x"2E9C288",
    x"2E9C018",
    x"2E9BDA8",
    x"2E9BB39",
    x"2E9B8CA",
    x"2E9B65C",
    x"2E9B3EF",
    x"2E9B182",
    x"2E9AF16",
    x"2E9ACAB",
    x"2E9AA40",
    x"2E9A7D6",
    x"2E9A56C",
    x"2E9A303",
    x"2E9A09B",
    x"2E99E33",
    x"2E99BCC",
    x"2E99965",
    x"2E996FF",
    x"2E99499",
    x"2E99235",
    x"2E98FD0",
    x"2E98D6D",
    x"2E98B0A",
    x"2E988A7",
    x"2E98645",
    x"2E983E4",
    x"2E98183",
    x"2E97F23",
    x"2E97CC4",
    x"2E97A65",
    x"2E97807",
    x"2E975A9",
    x"2E9734C",
    x"2E970EF",
    x"2E96E93",
    x"2E96C38",
    x"2E969DD",
    x"2E96783",
    x"2E96529",
    x"2E962D0",
    x"2E96078",
    x"2E95E20",
    x"2E95BC9",
    x"2E95972",
    x"2E9571C",
    x"2E954C7",
    x"2E95272",
    x"2E9501D",
    x"2E94DCA",
    x"2E94B77",
    x"2E94924",
    x"2E946D2",
    x"2E94481",
    x"2E94230",
    x"2E93FDF",
    x"2E93D90",
    x"2E93B41",
    x"2E938F2",
    x"2E936A4",
    x"2E93457",
    x"2E9320A",
    x"2E92FBE",
    x"2E92D72",
    x"2E92B27",
    x"2E928DD",
    x"2E92693",
    x"2E92449",
    x"2E92201",
    x"2E91FB8",
    x"2E91D71",
    x"2E91B2A",
    x"2E918E3",
    x"2E9169D",
    x"2E91458",
    x"2E91213",
    x"2E90FCF",
    x"2E90D8B",
    x"2E90B48",
    x"2E90905",
    x"2E906C3",
    x"2E90482",
    x"2E90241",
    x"2E90001",
    x"2E8FDC1",
    x"2E8FB82",
    x"2E8F943",
    x"2E8F705",
    x"2E8F4C8",
    x"2E8F28B",
    x"2E8F04F",
    x"2E8EE13",
    x"2E8EBD8",
    x"2E8E99D",
    x"2E8E763",
    x"2E8E529",
    x"2E8E2F0",
    x"2E8E0B8",
    x"2E8DE80",
    x"2E8DC49",
    x"2E8DA12",
    x"2E8D7DB",
    x"2E8D5A6",
    x"2E8D371",
    x"2E8D13C",
    x"2E8CF08",
    x"2E8CCD5",
    x"2E8CAA2",
    x"2E8C86F",
    x"2E8C63D",
    x"2E8C40C",
    x"2E8C1DB",
    x"2E8BFAB",
    x"2E8BD7C",
    x"2E8BB4C",
    x"2E8B91E",
    x"2E8B6F0",
    x"2E8B4C2",
    x"2E8B296",
    x"2E8B069",
    x"2E8AE3D",
    x"2E8AC12",
    x"2E8A9E7",
    x"2E8A7BD",
    x"2E8A593",
    x"2E8A36A",
    x"2E8A142",
    x"2E89F1A",
    x"2E89CF2",
    x"2E89ACB",
    x"2E898A5",
    x"2E8967F",
    x"2E89459",
    x"2E89235",
    x"2E89010",
    x"2E88DED",
    x"2E88BC9",
    x"2E889A7",
    x"2E88785",
    x"2E88563",
    x"2E88342",
    x"2E88121",
    x"2E87F01",
    x"2E87CE2",
    x"2E87AC3",
    x"2E878A4",
    x"2E87687",
    x"2E87469",
    x"2E8724C",
    x"2E87030",
    x"2E86E14",
    x"2E86BF9",
    x"2E869DE",
    x"2E867C4",
    x"2E865AA",
    x"2E86391",
    x"2E86179",
    x"2E85F61",
    x"2E85D49",
    x"2E85B32",
    x"2E8591B",
    x"2E85705",
    x"2E854F0",
    x"2E852DB",
    x"2E850C6",
    x"2E84EB2",
    x"2E84C9F",
    x"2E84A8C",
    x"2E8487A",
    x"2E84668",
    x"2E84457",
    x"2E84246",
    x"2E84035",
    x"2E83E26",
    x"2E83C16",
    x"2E83A08",
    x"2E837F9",
    x"2E835EC",
    x"2E833DE",
    x"2E831D2",
    x"2E82FC5",
    x"2E82DBA",
    x"2E82BAF",
    x"2E829A4",
    x"2E8279A",
    x"2E82590",
    x"2E82387",
    x"2E8217E",
    x"2E81F76",
    x"2E81D6F",
    x"2E81B68",
    x"2E81961",
    x"2E8175B",
    x"2E81555",
    x"2E81350",
    x"2E8114C",
    x"2E80F48",
    x"2E80D44",
    x"2E80B41",
    x"2E8093E",
    x"2E8073C",
    x"2E8053B",
    x"2E8033A",
    x"2E80139",
    x"2E7FE73",
    x"2E7FA73",
    x"2E7F675",
    x"2E7F278",
    x"2E7EE7C",
    x"2E7EA81",
    x"2E7E687",
    x"2E7E28E",
    x"2E7DE96",
    x"2E7DA9E",
    x"2E7D6A8",
    x"2E7D2B3",
    x"2E7CEBF",
    x"2E7CACC",
    x"2E7C6D9",
    x"2E7C2E8",
    x"2E7BEF8",
    x"2E7BB09",
    x"2E7B71B",
    x"2E7B32D",
    x"2E7AF41",
    x"2E7AB56",
    x"2E7A76B",
    x"2E7A382",
    x"2E79F99",
    x"2E79BB2",
    x"2E797CC",
    x"2E793E6",
    x"2E79002",
    x"2E78C1E",
    x"2E7883C",
    x"2E7845A",
    x"2E78079",
    x"2E77C9A",
    x"2E778BB",
    x"2E774DD",
    x"2E77101",
    x"2E76D25",
    x"2E7694A",
    x"2E76570",
    x"2E76197",
    x"2E75DC0",
    x"2E759E9",
    x"2E75613",
    x"2E7523E",
    x"2E74E69",
    x"2E74A96",
    x"2E746C4",
    x"2E742F3",
    x"2E73F23",
    x"2E73B53",
    x"2E73785",
    x"2E733B8",
    x"2E72FEB",
    x"2E72C20",
    x"2E72855",
    x"2E7248B",
    x"2E720C3",
    x"2E71CFB",
    x"2E71934",
    x"2E7156E",
    x"2E711AA",
    x"2E70DE6",
    x"2E70A23",
    x"2E70661",
    x"2E7029F",
    x"2E6FEDF",
    x"2E6FB20",
    x"2E6F762",
    x"2E6F3A4",
    x"2E6EFE8",
    x"2E6EC2C",
    x"2E6E872",
    x"2E6E4B8",
    x"2E6E0FF",
    x"2E6DD48",
    x"2E6D991",
    x"2E6D5DB",
    x"2E6D226",
    x"2E6CE72",
    x"2E6CABF",
    x"2E6C70C",
    x"2E6C35B",
    x"2E6BFAB",
    x"2E6BBFB",
    x"2E6B84D",
    x"2E6B49F",
    x"2E6B0F2",
    x"2E6AD47",
    x"2E6A99C",
    x"2E6A5F2",
    x"2E6A249",
    x"2E69EA1",
    x"2E69AFA",
    x"2E69753",
    x"2E693AE",
    x"2E69009",
    x"2E68C66",
    x"2E688C3",
    x"2E68521",
    x"2E68181",
    x"2E67DE1",
    x"2E67A42",
    x"2E676A4",
    x"2E67306",
    x"2E66F6A",
    x"2E66BCF",
    x"2E66834",
    x"2E6649B",
    x"2E66102",
    x"2E65D6A",
    x"2E659D3",
    x"2E6563D",
    x"2E652A8",
    x"2E64F14",
    x"2E64B80",
    x"2E647EE",
    x"2E6445D",
    x"2E640CC",
    x"2E63D3C",
    x"2E639AD",
    x"2E6361F",
    x"2E63292",
    x"2E62F06",
    x"2E62B7B",
    x"2E627F0",
    x"2E62467",
    x"2E620DE",
    x"2E61D56",
    x"2E619CF",
    x"2E61649",
    x"2E612C4",
    x"2E60F40",
    x"2E60BBD",
    x"2E6083A",
    x"2E604B8",
    x"2E60138",
    x"2E5FDB8",
    x"2E5FA39",
    x"2E5F6BB",
    x"2E5F33E",
    x"2E5EFC1",
    x"2E5EC46",
    x"2E5E8CB",
    x"2E5E551",
    x"2E5E1D8",
    x"2E5DE60",
    x"2E5DAE9",
    x"2E5D773",
    x"2E5D3FD",
    x"2E5D089",
    x"2E5CD15",
    x"2E5C9A2",
    x"2E5C630",
    x"2E5C2BF",
    x"2E5BF4F",
    x"2E5BBE0",
    x"2E5B871",
    x"2E5B503",
    x"2E5B197",
    x"2E5AE2B",
    x"2E5AABF",
    x"2E5A755",
    x"2E5A3EC",
    x"2E5A083",
    x"2E59D1C",
    x"2E599B5",
    x"2E5964F",
    x"2E592EA",
    x"2E58F85",
    x"2E58C22",
    x"2E588BF",
    x"2E5855D",
    x"2E581FC",
    x"2E57E9C",
    x"2E57B3D",
    x"2E577DF",
    x"2E57481",
    x"2E57124",
    x"2E56DC9",
    x"2E56A6E",
    x"2E56713",
    x"2E563BA",
    x"2E56062",
    x"2E55D0A",
    x"2E559B3",
    x"2E5565D",
    x"2E55308",
    x"2E54FB4",
    x"2E54C60",
    x"2E5490D",
    x"2E545BB",
    x"2E5426A",
    x"2E53F1A",
    x"2E53BCB",
    x"2E5387C",
    x"2E5352F",
    x"2E531E2",
    x"2E52E96",
    x"2E52B4A",
    x"2E52800",
    x"2E524B6",
    x"2E5216E",
    x"2E51E26",
    x"2E51ADF",
    x"2E51798",
    x"2E51453",
    x"2E5110E",
    x"2E50DCA",
    x"2E50A87",
    x"2E50745",
    x"2E50404",
    x"2E500C3",
    x"2E4FD83",
    x"2E4FA44",
    x"2E4F706",
    x"2E4F3C9",
    x"2E4F08C",
    x"2E4ED50",
    x"2E4EA16",
    x"2E4E6DB",
    x"2E4E3A2",
    x"2E4E06A",
    x"2E4DD32",
    x"2E4D9FB",
    x"2E4D6C5",
    x"2E4D390",
    x"2E4D05B",
    x"2E4CD27",
    x"2E4C9F5",
    x"2E4C6C2",
    x"2E4C391",
    x"2E4C061",
    x"2E4BD31",
    x"2E4BA02",
    x"2E4B6D4",
    x"2E4B3A7",
    x"2E4B07A",
    x"2E4AD4E",
    x"2E4AA24",
    x"2E4A6F9",
    x"2E4A3D0",
    x"2E4A0A7",
    x"2E49D80",
    x"2E49A59",
    x"2E49733",
    x"2E4940D",
    x"2E490E8",
    x"2E48DC5",
    x"2E48AA2",
    x"2E4877F",
    x"2E4845E",
    x"2E4813D",
    x"2E47E1D",
    x"2E47AFE",
    x"2E477E0",
    x"2E474C2",
    x"2E471A5",
    x"2E46E89",
    x"2E46B6E",
    x"2E46854",
    x"2E4653A",
    x"2E46221",
    x"2E45F09",
    x"2E45BF1",
    x"2E458DB",
    x"2E455C5",
    x"2E452B0",
    x"2E44F9C",
    x"2E44C88",
    x"2E44975",
    x"2E44663",
    x"2E44352",
    x"2E44042",
    x"2E43D32",
    x"2E43A23",
    x"2E43715",
    x"2E43408",
    x"2E430FB",
    x"2E42DEF",
    x"2E42AE4",
    x"2E427DA",
    x"2E424D0",
    x"2E421C7",
    x"2E41EBF",
    x"2E41BB8",
    x"2E418B1",
    x"2E415AC",
    x"2E412A7",
    x"2E40FA2",
    x"2E40C9F",
    x"2E4099C",
    x"2E4069A",
    x"2E40399",
    x"2E40098",
    x"2E3FD98",
    x"2E3FA99",
    x"2E3F79B",
    x"2E3F49E",
    x"2E3F1A1",
    x"2E3EEA5",
    x"2E3EBA9",
    x"2E3E8AF",
    x"2E3E5B5",
    x"2E3E2BC",
    x"2E3DFC4",
    x"2E3DCCC",
    x"2E3D9D5",
    x"2E3D6DF",
    x"2E3D3EA",
    x"2E3D0F5",
    x"2E3CE01",
    x"2E3CB0E",
    x"2E3C81C",
    x"2E3C52A",
    x"2E3C239",
    x"2E3BF49",
    x"2E3BC5A",
    x"2E3B96B",
    x"2E3B67D",
    x"2E3B390",
    x"2E3B0A3",
    x"2E3ADB7",
    x"2E3AACC",
    x"2E3A7E2",
    x"2E3A4F8",
    x"2E3A20F",
    x"2E39F27",
    x"2E39C40",
    x"2E39959",
    x"2E39673",
    x"2E3938E",
    x"2E390A9",
    x"2E38DC6",
    x"2E38AE3",
    x"2E38800",
    x"2E3851F",
    x"2E3823E",
    x"2E37F5D",
    x"2E37C7E",
    x"2E3799F",
    x"2E376C1",
    x"2E373E4",
    x"2E37107",
    x"2E36E2B",
    x"2E36B50",
    x"2E36876",
    x"2E3659C",
    x"2E362C3",
    x"2E35FEA",
    x"2E35D13",
    x"2E35A3C",
    x"2E35766",
    x"2E35490",
    x"2E351BB",
    x"2E34EE7",
    x"2E34C14",
    x"2E34941",
    x"2E3466F",
    x"2E3439E",
    x"2E340CE",
    x"2E33DFE",
    x"2E33B2F",
    x"2E33860",
    x"2E33592",
    x"2E332C5",
    x"2E32FF9",
    x"2E32D2D",
    x"2E32A62",
    x"2E32798",
    x"2E324CF",
    x"2E32206",
    x"2E31F3E",
    x"2E31C76",
    x"2E319AF",
    x"2E316E9",
    x"2E31424",
    x"2E3115F",
    x"2E30E9B",
    x"2E30BD8",
    x"2E30915",
    x"2E30653",
    x"2E30392",
    x"2E300D2",
    x"2E2FE12",
    x"2E2FB53",
    x"2E2F894",
    x"2E2F5D6",
    x"2E2F319",
    x"2E2F05D",
    x"2E2EDA1",
    x"2E2EAE6",
    x"2E2E82C",
    x"2E2E572",
    x"2E2E2B9",
    x"2E2E000",
    x"2E2DD49",
    x"2E2DA92",
    x"2E2D7DB",
    x"2E2D526",
    x"2E2D271",
    x"2E2CFBD",
    x"2E2CD09",
    x"2E2CA56",
    x"2E2C7A4",
    x"2E2C4F2",
    x"2E2C241",
    x"2E2BF91",
    x"2E2BCE2",
    x"2E2BA33",
    x"2E2B785",
    x"2E2B4D7",
    x"2E2B22A",
    x"2E2AF7E",
    x"2E2ACD2",
    x"2E2AA27",
    x"2E2A77D",
    x"2E2A4D4",
    x"2E2A22B",
    x"2E29F83",
    x"2E29CDB",
    x"2E29A34",
    x"2E2978E",
    x"2E294E8",
    x"2E29244",
    x"2E28F9F",
    x"2E28CFC",
    x"2E28A59",
    x"2E287B7",
    x"2E28515",
    x"2E28274",
    x"2E27FD4",
    x"2E27D34",
    x"2E27A95",
    x"2E277F7",
    x"2E27559",
    x"2E272BC",
    x"2E27020",
    x"2E26D84",
    x"2E26AE9",
    x"2E2684F",
    x"2E265B5",
    x"2E2631C",
    x"2E26083",
    x"2E25DEC",
    x"2E25B54",
    x"2E258BE",
    x"2E25628",
    x"2E25393",
    x"2E250FE",
    x"2E24E6A",
    x"2E24BD7",
    x"2E24944",
    x"2E246B2",
    x"2E24421",
    x"2E24190",
    x"2E23F00",
    x"2E23C71",
    x"2E239E2",
    x"2E23754",
    x"2E234C6",
    x"2E23239",
    x"2E22FAD",
    x"2E22D22",
    x"2E22A97",
    x"2E2280C",
    x"2E22583",
    x"2E222FA",
    x"2E22071",
    x"2E21DE9",
    x"2E21B62",
    x"2E218DC",
    x"2E21656",
    x"2E213D0",
    x"2E2114C",
    x"2E20EC8",
    x"2E20C44",
    x"2E209C2",
    x"2E20740",
    x"2E204BE",
    x"2E2023D",
    x"2E1FFBD",
    x"2E1FD3D",
    x"2E1FABE",
    x"2E1F840",
    x"2E1F5C2",
    x"2E1F345",
    x"2E1F0C9",
    x"2E1EE4D",
    x"2E1EBD1",
    x"2E1E957",
    x"2E1E6DD",
    x"2E1E463",
    x"2E1E1EB",
    x"2E1DF72",
    x"2E1DCFB",
    x"2E1DA84",
    x"2E1D80E",
    x"2E1D598",
    x"2E1D323",
    x"2E1D0AE",
    x"2E1CE3A",
    x"2E1CBC7",
    x"2E1C955",
    x"2E1C6E3",
    x"2E1C471",
    x"2E1C200",
    x"2E1BF90",
    x"2E1BD21",
    x"2E1BAB2",
    x"2E1B843",
    x"2E1B5D5",
    x"2E1B368",
    x"2E1B0FC",
    x"2E1AE90",
    x"2E1AC24",
    x"2E1A9BA",
    x"2E1A750",
    x"2E1A4E6",
    x"2E1A27D",
    x"2E1A015",
    x"2E19DAD",
    x"2E19B46",
    x"2E198DF",
    x"2E19679",
    x"2E19414",
    x"2E191AF",
    x"2E18F4B",
    x"2E18CE8",
    x"2E18A85",
    x"2E18823",
    x"2E185C1",
    x"2E18360",
    x"2E180FF",
    x"2E17E9F",
    x"2E17C40",
    x"2E179E1",
    x"2E17783",
    x"2E17525",
    x"2E172C8",
    x"2E1706C",
    x"2E16E10",
    x"2E16BB5",
    x"2E1695A",
    x"2E16700",
    x"2E164A7",
    x"2E1624E",
    x"2E15FF6",
    x"2E15D9E",
    x"2E15B47",
    x"2E158F0",
    x"2E1569A",
    x"2E15445",
    x"2E151F0",
    x"2E14F9C",
    x"2E14D48",
    x"2E14AF5",
    x"2E148A3",
    x"2E14651",
    x"2E14400",
    x"2E141AF",
    x"2E13F5F",
    x"2E13D0F",
    x"2E13AC0",
    x"2E13872",
    x"2E13624",
    x"2E133D7",
    x"2E1318A",
    x"2E12F3E",
    x"2E12CF3",
    x"2E12AA8",
    x"2E1285D",
    x"2E12613",
    x"2E123CA",
    x"2E12182",
    x"2E11F39",
    x"2E11CF2",
    x"2E11AAB",
    x"2E11865",
    x"2E1161F",
    x"2E113DA",
    x"2E11195",
    x"2E10F51",
    x"2E10D0D",
    x"2E10ACA",
    x"2E10888",
    x"2E10646",
    x"2E10405",
    x"2E101C4",
    x"2E0FF84",
    x"2E0FD44",
    x"2E0FB05",
    x"2E0F8C7",
    x"2E0F689",
    x"2E0F44B",
    x"2E0F20F",
    x"2E0EFD2",
    x"2E0ED97",
    x"2E0EB5C",
    x"2E0E921",
    x"2E0E6E7",
    x"2E0E4AE",
    x"2E0E275",
    x"2E0E03C",
    x"2E0DE05",
    x"2E0DBCD",
    x"2E0D997",
    x"2E0D761",
    x"2E0D52B",
    x"2E0D2F6",
    x"2E0D0C1",
    x"2E0CE8E",
    x"2E0CC5A",
    x"2E0CA27",
    x"2E0C7F5",
    x"2E0C5C3",
    x"2E0C392",
    x"2E0C162",
    x"2E0BF32",
    x"2E0BD02",
    x"2E0BAD3",
    x"2E0B8A5",
    x"2E0B677",
    x"2E0B449",
    x"2E0B21D",
    x"2E0AFF0",
    x"2E0ADC5",
    x"2E0AB99",
    x"2E0A96F",
    x"2E0A745",
    x"2E0A51B",
    x"2E0A2F2",
    x"2E0A0CA",
    x"2E09EA2",
    x"2E09C7A",
    x"2E09A54",
    x"2E0982D",
    x"2E09607",
    x"2E093E2",
    x"2E091BD",
    x"2E08F99",
    x"2E08D76",
    x"2E08B53",
    x"2E08930",
    x"2E0870E",
    x"2E084ED",
    x"2E082CC",
    x"2E080AB",
    x"2E07E8B",
    x"2E07C6C",
    x"2E07A4D",
    x"2E0782F",
    x"2E07611",
    x"2E073F4",
    x"2E071D7",
    x"2E06FBB",
    x"2E06D9F",
    x"2E06B84",
    x"2E06969",
    x"2E0674F",
    x"2E06536",
    x"2E0631D",
    x"2E06104",
    x"2E05EEC",
    x"2E05CD5",
    x"2E05ABE",
    x"2E058A7",
    x"2E05691",
    x"2E0547C",
    x"2E05267",
    x"2E05053",
    x"2E04E3F",
    x"2E04C2C",
    x"2E04A19",
    x"2E04807",
    x"2E045F5",
    x"2E043E4",
    x"2E041D3",
    x"2E03FC3",
    x"2E03DB3",
    x"2E03BA4",
    x"2E03995",
    x"2E03787",
    x"2E03579",
    x"2E0336C",
    x"2E03160",
    x"2E02F54",
    x"2E02D48",
    x"2E02B3D",
    x"2E02932",
    x"2E02728",
    x"2E0251F",
    x"2E02316",
    x"2E0210D",
    x"2E01F05",
    x"2E01CFE",
    x"2E01AF7",
    x"2E018F0",
    x"2E016EA",
    x"2E014E5",
    x"2E012E0",
    x"2E010DB",
    x"2E00ED7",
    x"2E00CD4",
    x"2E00AD1",
    x"2E008CF",
    x"2E006CD",
    x"2E004CB",
    x"2E002CA",
    x"2E000CA",
    x"2DFFD94",
    x"2DFF995",
    x"2DFF597",
    x"2DFF19A",
    x"2DFED9F",
    x"2DFE9A4",
    x"2DFE5AA",
    x"2DFE1B1",
    x"2DFDDB9",
    x"2DFD9C2",
    x"2DFD5CC",
    x"2DFD1D7",
    x"2DFCDE3",
    x"2DFC9F0",
    x"2DFC5FE",
    x"2DFC20D",
    x"2DFBE1D",
    x"2DFBA2E",
    x"2DFB640",
    x"2DFB253",
    x"2DFAE67",
    x"2DFAA7C",
    x"2DFA692",
    x"2DFA2A8",
    x"2DF9EC0",
    x"2DF9AD9",
    x"2DF96F3",
    x"2DF930E",
    x"2DF8F29",
    x"2DF8B46",
    x"2DF8764",
    x"2DF8382",
    x"2DF7FA2",
    x"2DF7BC2",
    x"2DF77E4",
    x"2DF7407",
    x"2DF702A",
    x"2DF6C4E",
    x"2DF6874",
    x"2DF649A",
    x"2DF60C2",
    x"2DF5CEA",
    x"2DF5913",
    x"2DF553D",
    x"2DF5168",
    x"2DF4D95",
    x"2DF49C2",
    x"2DF45F0",
    x"2DF421F",
    x"2DF3E4F",
    x"2DF3A80",
    x"2DF36B1",
    x"2DF32E4",
    x"2DF2F18",
    x"2DF2B4D",
    x"2DF2782",
    x"2DF23B9",
    x"2DF1FF0",
    x"2DF1C29",
    x"2DF1862",
    x"2DF149D",
    x"2DF10D8",
    x"2DF0D14",
    x"2DF0952",
    x"2DF0590",
    x"2DF01CF",
    x"2DEFE0F",
    x"2DEFA50",
    x"2DEF692",
    x"2DEF2D4",
    x"2DEEF18",
    x"2DEEB5D",
    x"2DEE7A3",
    x"2DEE3E9",
    x"2DEE031",
    x"2DEDC79",
    x"2DED8C2",
    x"2DED50D",
    x"2DED158",
    x"2DECDA4",
    x"2DEC9F1",
    x"2DEC63F",
    x"2DEC28E",
    x"2DEBEDE",
    x"2DEBB2E",
    x"2DEB780",
    x"2DEB3D3",
    x"2DEB026",
    x"2DEAC7B",
    x"2DEA8D0",
    x"2DEA526",
    x"2DEA17D",
    x"2DE9DD5",
    x"2DE9A2E",
    x"2DE9688",
    x"2DE92E3",
    x"2DE8F3F",
    x"2DE8B9C",
    x"2DE87F9",
    x"2DE8458",
    x"2DE80B7",
    x"2DE7D17",
    x"2DE7978",
    x"2DE75DA",
    x"2DE723D",
    x"2DE6EA1",
    x"2DE6B06",
    x"2DE676C",
    x"2DE63D2",
    x"2DE603A",
    x"2DE5CA2",
    x"2DE590C",
    x"2DE5576",
    x"2DE51E1",
    x"2DE4E4D",
    x"2DE4ABA",
    x"2DE4727",
    x"2DE4396",
    x"2DE4006",
    x"2DE3C76",
    x"2DE38E7",
    x"2DE355A",
    x"2DE31CD",
    x"2DE2E41",
    x"2DE2AB6",
    x"2DE272B",
    x"2DE23A2",
    x"2DE201A",
    x"2DE1C92",
    x"2DE190B",
    x"2DE1585",
    x"2DE1201",
    x"2DE0E7C",
    x"2DE0AF9",
    x"2DE0777",
    x"2DE03F6",
    x"2DE0075",
    x"2DDFCF5",
    x"2DDF977",
    x"2DDF5F9",
    x"2DDF27C",
    x"2DDEEFF",
    x"2DDEB84",
    x"2DDE80A",
    x"2DDE490",
    x"2DDE117",
    x"2DDDD9F",
    x"2DDDA28",
    x"2DDD6B2",
    x"2DDD33D",
    x"2DDCFC9",
    x"2DDCC55",
    x"2DDC8E3",
    x"2DDC571",
    x"2DDC200",
    x"2DDBE90",
    x"2DDBB21",
    x"2DDB7B2",
    x"2DDB445",
    x"2DDB0D8",
    x"2DDAD6C",
    x"2DDAA01",
    x"2DDA697",
    x"2DDA32E",
    x"2DD9FC6",
    x"2DD9C5E",
    x"2DD98F8",
    x"2DD9592",
    x"2DD922D",
    x"2DD8EC9",
    x"2DD8B65",
    x"2DD8803",
    x"2DD84A1",
    x"2DD8141",
    x"2DD7DE1",
    x"2DD7A82",
    x"2DD7723",
    x"2DD73C6",
    x"2DD706A",
    x"2DD6D0E",
    x"2DD69B3",
    x"2DD6659",
    x"2DD6300",
    x"2DD5FA8",
    x"2DD5C50",
    x"2DD58F9",
    x"2DD55A4",
    x"2DD524F",
    x"2DD4EFA",
    x"2DD4BA7",
    x"2DD4855",
    x"2DD4503",
    x"2DD41B2",
    x"2DD3E62",
    x"2DD3B13",
    x"2DD37C5",
    x"2DD3477",
    x"2DD312A",
    x"2DD2DDE",
    x"2DD2A93",
    x"2DD2749",
    x"2DD2400",
    x"2DD20B7",
    x"2DD1D6F",
    x"2DD1A28",
    x"2DD16E2",
    x"2DD139D",
    x"2DD1058",
    x"2DD0D15",
    x"2DD09D2",
    x"2DD0690",
    x"2DD034F",
    x"2DD000E",
    x"2DCFCCF",
    x"2DCF990",
    x"2DCF652",
    x"2DCF315",
    x"2DCEFD8",
    x"2DCEC9D",
    x"2DCE962",
    x"2DCE628",
    x"2DCE2EF",
    x"2DCDFB7",
    x"2DCDC7F",
    x"2DCD948",
    x"2DCD612",
    x"2DCD2DD",
    x"2DCCFA9",
    x"2DCCC75",
    x"2DCC943",
    x"2DCC611",
    x"2DCC2E0",
    x"2DCBFAF",
    x"2DCBC80",
    x"2DCB951",
    x"2DCB623",
    x"2DCB2F6",
    x"2DCAFCA",
    x"2DCAC9E",
    x"2DCA973",
    x"2DCA649",
    x"2DCA320",
    x"2DC9FF8",
    x"2DC9CD0",
    x"2DC99A9",
    x"2DC9683",
    x"2DC935E",
    x"2DC903A",
    x"2DC8D16",
    x"2DC89F3",
    x"2DC86D1",
    x"2DC83B0",
    x"2DC808F",
    x"2DC7D70",
    x"2DC7A51",
    x"2DC7732",
    x"2DC7415",
    x"2DC70F8",
    x"2DC6DDC",
    x"2DC6AC1",
    x"2DC67A7",
    x"2DC648E",
    x"2DC6175",
    x"2DC5E5D",
    x"2DC5B46",
    x"2DC582F",
    x"2DC551A",
    x"2DC5205",
    x"2DC4EF1",
    x"2DC4BDD",
    x"2DC48CB",
    x"2DC45B9",
    x"2DC42A8",
    x"2DC3F97",
    x"2DC3C88",
    x"2DC3979",
    x"2DC366B",
    x"2DC335E",
    x"2DC3052",
    x"2DC2D46",
    x"2DC2A3B",
    x"2DC2731",
    x"2DC2427",
    x"2DC211F",
    x"2DC1E17",
    x"2DC1B10",
    x"2DC1809",
    x"2DC1504",
    x"2DC11FF",
    x"2DC0EFB",
    x"2DC0BF7",
    x"2DC08F5",
    x"2DC05F3",
    x"2DC02F2",
    x"2DBFFF1",
    x"2DBFCF2",
    x"2DBF9F3",
    x"2DBF6F5",
    x"2DBF3F7",
    x"2DBF0FB",
    x"2DBEDFF",
    x"2DBEB04",
    x"2DBE809",
    x"2DBE510",
    x"2DBE217",
    x"2DBDF1F",
    x"2DBDC27",
    x"2DBD931",
    x"2DBD63B",
    x"2DBD345",
    x"2DBD051",
    x"2DBCD5D",
    x"2DBCA6A",
    x"2DBC778",
    x"2DBC487",
    x"2DBC196",
    x"2DBBEA6",
    x"2DBBBB6",
    x"2DBB8C8",
    x"2DBB5DA",
    x"2DBB2ED",
    x"2DBB001",
    x"2DBAD15",
    x"2DBAA2A",
    x"2DBA740",
    x"2DBA456",
    x"2DBA16E",
    x"2DB9E86",
    x"2DB9B9E",
    x"2DB98B8",
    x"2DB95D2",
    x"2DB92ED",
    x"2DB9009",
    x"2DB8D25",
    x"2DB8A42",
    x"2DB8760",
    x"2DB847E",
    x"2DB819E",
    x"2DB7EBE",
    x"2DB7BDE",
    x"2DB7900",
    x"2DB7622",
    x"2DB7345",
    x"2DB7068",
    x"2DB6D8C",
    x"2DB6AB1",
    x"2DB67D7",
    x"2DB64FD",
    x"2DB6225",
    x"2DB5F4C",
    x"2DB5C75",
    x"2DB599E",
    x"2DB56C8",
    x"2DB53F3",
    x"2DB511E",
    x"2DB4E4A",
    x"2DB4B77",
    x"2DB48A4",
    x"2DB45D3",
    x"2DB4301",
    x"2DB4031",
    x"2DB3D61",
    x"2DB3A92",
    x"2DB37C4",
    x"2DB34F7",
    x"2DB322A",
    x"2DB2F5D",
    x"2DB2C92",
    x"2DB29C7",
    x"2DB26FD",
    x"2DB2434",
    x"2DB216B",
    x"2DB1EA3",
    x"2DB1BDC",
    x"2DB1915",
    x"2DB164F",
    x"2DB138A",
    x"2DB10C5",
    x"2DB0E01",
    x"2DB0B3E",
    x"2DB087C",
    x"2DB05BA",
    x"2DB02F9",
    x"2DB0039",
    x"2DAFD79",
    x"2DAFABA",
    x"2DAF7FC",
    x"2DAF53E",
    x"2DAF281",
    x"2DAEFC5",
    x"2DAED09",
    x"2DAEA4E",
    x"2DAE794",
    x"2DAE4DA",
    x"2DAE221",
    x"2DADF69",
    x"2DADCB2",
    x"2DAD9FB",
    x"2DAD745",
    x"2DAD48F",
    x"2DAD1DA",
    x"2DACF26",
    x"2DACC73",
    x"2DAC9C0",
    x"2DAC70E",
    x"2DAC45D",
    x"2DAC1AC",
    x"2DABEFC",
    x"2DABC4C",
    x"2DAB99E",
    x"2DAB6F0",
    x"2DAB442",
    x"2DAB195",
    x"2DAAEE9",
    x"2DAAC3E",
    x"2DAA993",
    x"2DAA6E9",
    x"2DAA440",
    x"2DAA197",
    x"2DA9EEF",
    x"2DA9C48",
    x"2DA99A1",
    x"2DA96FB",
    x"2DA9455",
    x"2DA91B1",
    x"2DA8F0C",
    x"2DA8C69",
    x"2DA89C6",
    x"2DA8724",
    x"2DA8483",
    x"2DA81E2",
    x"2DA7F42",
    x"2DA7CA2",
    x"2DA7A03",
    x"2DA7765",
    x"2DA74C8",
    x"2DA722B",
    x"2DA6F8F",
    x"2DA6CF3",
    x"2DA6A58",
    x"2DA67BE",
    x"2DA6524",
    x"2DA628B",
    x"2DA5FF3",
    x"2DA5D5B",
    x"2DA5AC4",
    x"2DA582E",
    x"2DA5598",
    x"2DA5303",
    x"2DA506F",
    x"2DA4DDB",
    x"2DA4B48",
    x"2DA48B5",
    x"2DA4623",
    x"2DA4392",
    x"2DA4102",
    x"2DA3E72",
    x"2DA3BE2",
    x"2DA3954",
    x"2DA36C6",
    x"2DA3438",
    x"2DA31AC",
    x"2DA2F20",
    x"2DA2C94",
    x"2DA2A09",
    x"2DA277F",
    x"2DA24F6",
    x"2DA226D",
    x"2DA1FE4",
    x"2DA1D5D",
    x"2DA1AD6",
    x"2DA184F",
    x"2DA15C9",
    x"2DA1344",
    x"2DA10C0",
    x"2DA0E3C",
    x"2DA0BB9",
    x"2DA0936",
    x"2DA06B4",
    x"2DA0433",
    x"2DA01B2",
    x"2D9FF32",
    x"2D9FCB2",
    x"2D9FA34",
    x"2D9F7B5",
    x"2D9F538",
    x"2D9F2BB",
    x"2D9F03E",
    x"2D9EDC3",
    x"2D9EB47",
    x"2D9E8CD",
    x"2D9E653",
    x"2D9E3DA",
    x"2D9E161",
    x"2D9DEE9",
    x"2D9DC72",
    x"2D9D9FB",
    x"2D9D785",
    x"2D9D50F",
    x"2D9D29A",
    x"2D9D026",
    x"2D9CDB2",
    x"2D9CB3F",
    x"2D9C8CC",
    x"2D9C65B",
    x"2D9C3E9",
    x"2D9C179",
    x"2D9BF09",
    x"2D9BC99",
    x"2D9BA2A",
    x"2D9B7BC",
    x"2D9B54E",
    x"2D9B2E1",
    x"2D9B075",
    x"2D9AE09",
    x"2D9AB9E",
    x"2D9A933",
    x"2D9A6C9",
    x"2D9A460",
    x"2D9A1F7",
    x"2D99F8F",
    x"2D99D27",
    x"2D99AC0",
    x"2D9985A",
    x"2D995F4",
    x"2D9938F",
    x"2D9912A",
    x"2D98EC6",
    x"2D98C63",
    x"2D98A00",
    x"2D9879E",
    x"2D9853C",
    x"2D982DB",
    x"2D9807B",
    x"2D97E1B",
    x"2D97BBC",
    x"2D9795D",
    x"2D976FF",
    x"2D974A2",
    x"2D97245",
    x"2D96FE9",
    x"2D96D8D",
    x"2D96B32",
    x"2D968D7",
    x"2D9667D",
    x"2D96424",
    x"2D961CB",
    x"2D95F73",
    x"2D95D1C",
    x"2D95AC5",
    x"2D9586E",
    x"2D95618",
    x"2D953C3",
    x"2D9516F",
    x"2D94F1A",
    x"2D94CC7",
    x"2D94A74",
    x"2D94822",
    x"2D945D0",
    x"2D9437F",
    x"2D9412E",
    x"2D93EDE",
    x"2D93C8F",
    x"2D93A40",
    x"2D937F2",
    x"2D935A4",
    x"2D93357",
    x"2D9310A",
    x"2D92EBE",
    x"2D92C73",
    x"2D92A28",
    x"2D927DE",
    x"2D92594",
    x"2D9234B",
    x"2D92103",
    x"2D91EBB",
    x"2D91C73",
    x"2D91A2C",
    x"2D917E6",
    x"2D915A0",
    x"2D9135B",
    x"2D91117",
    x"2D90ED3",
    x"2D90C8F",
    x"2D90A4C",
    x"2D9080A",
    x"2D905C8",
    x"2D90387",
    x"2D90147",
    x"2D8FF07",
    x"2D8FCC7",
    x"2D8FA88",
    x"2D8F84A",
    x"2D8F60C",
    x"2D8F3CF",
    x"2D8F192",
    x"2D8EF56",
    x"2D8ED1B",
    x"2D8EAE0",
    x"2D8E8A5",
    x"2D8E66B",
    x"2D8E432",
    x"2D8E1F9",
    x"2D8DFC1",
    x"2D8DD89",
    x"2D8DB52",
    x"2D8D91C",
    x"2D8D6E6",
    x"2D8D4B0",
    x"2D8D27B",
    x"2D8D047",
    x"2D8CE13",
    x"2D8CBE0",
    x"2D8C9AD",
    x"2D8C77B",
    x"2D8C549",
    x"2D8C318",
    x"2D8C0E8",
    x"2D8BEB8",
    x"2D8BC89",
    x"2D8BA5A",
    x"2D8B82B",
    x"2D8B5FE",
    x"2D8B3D0",
    x"2D8B1A4",
    x"2D8AF78",
    x"2D8AD4C",
    x"2D8AB21",
    x"2D8A8F6",
    x"2D8A6CC",
    x"2D8A4A3",
    x"2D8A27A",
    x"2D8A052",
    x"2D89E2A",
    x"2D89C03",
    x"2D899DC",
    x"2D897B6",
    x"2D89590",
    x"2D8936B",
    x"2D89146",
    x"2D88F22",
    x"2D88CFF",
    x"2D88ADC",
    x"2D888B9",
    x"2D88697",
    x"2D88476",
    x"2D88255",
    x"2D88035",
    x"2D87E15",
    x"2D87BF6",
    x"2D879D7",
    x"2D877B9",
    x"2D8759B",
    x"2D8737E",
    x"2D87161",
    x"2D86F45",
    x"2D86D2A",
    x"2D86B0F",
    x"2D868F4",
    x"2D866DA",
    x"2D864C1",
    x"2D862A8",
    x"2D86090",
    x"2D85E78",
    x"2D85C60",
    x"2D85A4A",
    x"2D85833",
    x"2D8561D",
    x"2D85408",
    x"2D851F3",
    x"2D84FDF",
    x"2D84DCB",
    x"2D84BB8",
    x"2D849A6",
    x"2D84793",
    x"2D84582",
    x"2D84371",
    x"2D84160",
    x"2D83F50",
    x"2D83D40",
    x"2D83B31",
    x"2D83923",
    x"2D83715",
    x"2D83507",
    x"2D832FA",
    x"2D830EE",
    x"2D82EE2",
    x"2D82CD6",
    x"2D82ACB",
    x"2D828C1",
    x"2D826B7",
    x"2D824AE",
    x"2D822A5",
    x"2D8209C",
    x"2D81E94",
    x"2D81C8D",
    x"2D81A86",
    x"2D81880",
    x"2D8167A",
    x"2D81474",
    x"2D81270",
    x"2D8106B",
    x"2D80E67",
    x"2D80C64",
    x"2D80A61",
    x"2D8085F",
    x"2D8065D",
    x"2D8045C",
    x"2D8025B",
    x"2D8005B",
    x"2D7FCB6",
    x"2D7F8B7",
    x"2D7F4B9",
    x"2D7F0BD",
    x"2D7ECC1",
    x"2D7E8C6",
    x"2D7E4CD",
    x"2D7E0D4",
    x"2D7DCDC",
    x"2D7D8E6",
    x"2D7D4F0",
    x"2D7D0FB",
    x"2D7CD07",
    x"2D7C915",
    x"2D7C523",
    x"2D7C132",
    x"2D7BD42",
    x"2D7B953",
    x"2D7B566",
    x"2D7B179",
    x"2D7AD8D",
    x"2D7A9A2",
    x"2D7A5B8",
    x"2D7A1CF",
    x"2D79DE7",
    x"2D79A00",
    x"2D7961A",
    x"2D79235",
    x"2D78E51",
    x"2D78A6E",
    x"2D7868C",
    x"2D782AB",
    x"2D77ECA",
    x"2D77AEB",
    x"2D7770D",
    x"2D77330",
    x"2D76F53",
    x"2D76B78",
    x"2D7679E",
    x"2D763C4",
    x"2D75FEC",
    x"2D75C14",
    x"2D7583E",
    x"2D75468",
    x"2D75093",
    x"2D74CC0",
    x"2D748ED",
    x"2D7451B",
    x"2D7414B",
    x"2D73D7B",
    x"2D739AC",
    x"2D735DE",
    x"2D73211",
    x"2D72E45",
    x"2D72A7A",
    x"2D726B0",
    x"2D722E6",
    x"2D71F1E",
    x"2D71B57",
    x"2D71790",
    x"2D713CB",
    x"2D71007",
    x"2D70C43",
    x"2D70880",
    x"2D704BF",
    x"2D700FE",
    x"2D6FD3E",
    x"2D6F97F",
    x"2D6F5C2",
    x"2D6F205",
    x"2D6EE49",
    x"2D6EA8D",
    x"2D6E6D3",
    x"2D6E31A",
    x"2D6DF62",
    x"2D6DBAA",
    x"2D6D7F4",
    x"2D6D43E",
    x"2D6D08A",
    x"2D6CCD6",
    x"2D6C923",
    x"2D6C572",
    x"2D6C1C1",
    x"2D6BE11",
    x"2D6BA62",
    x"2D6B6B3",
    x"2D6B306",
    x"2D6AF5A",
    x"2D6ABAF",
    x"2D6A804",
    x"2D6A45B",
    x"2D6A0B2",
    x"2D69D0A",
    x"2D69963",
    x"2D695BD",
    x"2D69219",
    x"2D68E74",
    x"2D68AD1",
    x"2D6872F",
    x"2D6838E",
    x"2D67FED",
    x"2D67C4E",
    x"2D678AF",
    x"2D67511",
    x"2D67175",
    x"2D66DD9",
    x"2D66A3E",
    x"2D666A4",
    x"2D6630A",
    x"2D65F72",
    x"2D65BDB",
    x"2D65844",
    x"2D654AE",
    x"2D6511A",
    x"2D64D86",
    x"2D649F3",
    x"2D64661",
    x"2D642D0",
    x"2D63F40",
    x"2D63BB0",
    x"2D63822",
    x"2D63494",
    x"2D63107",
    x"2D62D7C",
    x"2D629F1",
    x"2D62667",
    x"2D622DD",
    x"2D61F55",
    x"2D61BCE",
    x"2D61847",
    x"2D614C2",
    x"2D6113D",
    x"2D60DB9",
    x"2D60A36",
    x"2D606B4",
    x"2D60333",
    x"2D5FFB2",
    x"2D5FC33",
    x"2D5F8B4",
    x"2D5F536",
    x"2D5F1BA",
    x"2D5EE3E",
    x"2D5EAC2",
    x"2D5E748",
    x"2D5E3CF",
    x"2D5E056",
    x"2D5DCDF",
    x"2D5D968",
    x"2D5D5F2",
    x"2D5D27D",
    x"2D5CF09",
    x"2D5CB95",
    x"2D5C823",
    x"2D5C4B1",
    x"2D5C141",
    x"2D5BDD1",
    x"2D5BA62",
    x"2D5B6F4",
    x"2D5B386",
    x"2D5B01A",
    x"2D5ACAE",
    x"2D5A943",
    x"2D5A5DA",
    x"2D5A270",
    x"2D59F08",
    x"2D59BA1",
    x"2D5983A",
    x"2D594D5",
    x"2D59170",
    x"2D58E0C",
    x"2D58AA9",
    x"2D58747",
    x"2D583E5",
    x"2D58085",
    x"2D57D25",
    x"2D579C6",
    x"2D57668",
    x"2D5730B",
    x"2D56FAF",
    x"2D56C53",
    x"2D568F9",
    x"2D5659F",
    x"2D56246",
    x"2D55EEE",
    x"2D55B96",
    x"2D55840",
    x"2D554EA",
    x"2D55195",
    x"2D54E41",
    x"2D54AEE",
    x"2D5479C",
    x"2D5444A",
    x"2D540FA",
    x"2D53DAA",
    x"2D53A5B",
    x"2D5370D",
    x"2D533BF",
    x"2D53073",
    x"2D52D27",
    x"2D529DC",
    x"2D52692",
    x"2D52349",
    x"2D52001",
    x"2D51CB9",
    x"2D51972",
    x"2D5162C",
    x"2D512E7",
    x"2D50FA3",
    x"2D50C5F",
    x"2D5091D",
    x"2D505DB",
    x"2D5029A",
    x"2D4FF59",
    x"2D4FC1A",
    x"2D4F8DB",
    x"2D4F59E",
    x"2D4F261",
    x"2D4EF24",
    x"2D4EBE9",
    x"2D4E8AE",
    x"2D4E575",
    x"2D4E23C",
    x"2D4DF04",
    x"2D4DBCC",
    x"2D4D896",
    x"2D4D560",
    x"2D4D22B",
    x"2D4CEF7",
    x"2D4CBC3",
    x"2D4C891",
    x"2D4C55F",
    x"2D4C22E",
    x"2D4BEFE",
    x"2D4BBCF",
    x"2D4B8A0",
    x"2D4B572",
    x"2D4B245",
    x"2D4AF19",
    x"2D4ABEE",
    x"2D4A8C3",
    x"2D4A59A",
    x"2D4A271",
    x"2D49F48",
    x"2D49C21",
    x"2D498FA",
    x"2D495D4",
    x"2D492AF",
    x"2D48F8B",
    x"2D48C68",
    x"2D48945",
    x"2D48623",
    x"2D48302",
    x"2D47FE1",
    x"2D47CC2",
    x"2D479A3",
    x"2D47685",
    x"2D47368",
    x"2D4704B",
    x"2D46D30",
    x"2D46A15",
    x"2D466FB",
    x"2D463E1",
    x"2D460C9",
    x"2D45DB1",
    x"2D45A9A",
    x"2D45784",
    x"2D4546E",
    x"2D45159",
    x"2D44E45",
    x"2D44B32",
    x"2D44820",
    x"2D4450E",
    x"2D441FD",
    x"2D43EED",
    x"2D43BDE",
    x"2D438CF",
    x"2D435C1",
    x"2D432B4",
    x"2D42FA8",
    x"2D42C9D",
    x"2D42992",
    x"2D42688",
    x"2D4237E",
    x"2D42076",
    x"2D41D6E",
    x"2D41A67",
    x"2D41761",
    x"2D4145C",
    x"2D41157",
    x"2D40E53",
    x"2D40B50",
    x"2D4084D",
    x"2D4054C",
    x"2D4024B",
    x"2D3FF4A",
    x"2D3FC4B",
    x"2D3F94C",
    x"2D3F64E",
    x"2D3F351",
    x"2D3F055",
    x"2D3ED59",
    x"2D3EA5E",
    x"2D3E764",
    x"2D3E46A",
    x"2D3E172",
    x"2D3DE7A",
    x"2D3DB82",
    x"2D3D88C",
    x"2D3D596",
    x"2D3D2A1",
    x"2D3CFAD",
    x"2D3CCB9",
    x"2D3C9C6",
    x"2D3C6D4",
    x"2D3C3E3",
    x"2D3C0F2",
    x"2D3BE02",
    x"2D3BB13",
    x"2D3B825",
    x"2D3B537",
    x"2D3B24A",
    x"2D3AF5E",
    x"2D3AC73",
    x"2D3A988",
    x"2D3A69E",
    x"2D3A3B5",
    x"2D3A0CC",
    x"2D39DE4",
    x"2D39AFD",
    x"2D39817",
    x"2D39531",
    x"2D3924C",
    x"2D38F68",
    x"2D38C84",
    x"2D389A2",
    x"2D386C0",
    x"2D383DE",
    x"2D380FE",
    x"2D37E1E",
    x"2D37B3F",
    x"2D37860",
    x"2D37582",
    x"2D372A5",
    x"2D36FC9",
    x"2D36CED",
    x"2D36A13",
    x"2D36738",
    x"2D3645F",
    x"2D36186",
    x"2D35EAE",
    x"2D35BD7",
    x"2D35900",
    x"2D3562A",
    x"2D35355",
    x"2D35081",
    x"2D34DAD",
    x"2D34ADA",
    x"2D34808",
    x"2D34536",
    x"2D34265",
    x"2D33F95",
    x"2D33CC5",
    x"2D339F6",
    x"2D33728",
    x"2D3345B",
    x"2D3318E",
    x"2D32EC2",
    x"2D32BF7",
    x"2D3292C",
    x"2D32662",
    x"2D32399",
    x"2D320D0",
    x"2D31E08",
    x"2D31B41",
    x"2D3187B",
    x"2D315B5",
    x"2D312F0",
    x"2D3102B",
    x"2D30D68",
    x"2D30AA5",
    x"2D307E2",
    x"2D30521",
    x"2D30260",
    x"2D2FFA0",
    x"2D2FCE0",
    x"2D2FA21",
    x"2D2F763",
    x"2D2F4A5",
    x"2D2F1E9",
    x"2D2EF2D",
    x"2D2EC71",
    x"2D2E9B6",
    x"2D2E6FC",
    x"2D2E443",
    x"2D2E18A",
    x"2D2DED2",
    x"2D2DC1B",
    x"2D2D964",
    x"2D2D6AE",
    x"2D2D3F9",
    x"2D2D144",
    x"2D2CE90",
    x"2D2CBDD",
    x"2D2C92A",
    x"2D2C678",
    x"2D2C3C7",
    x"2D2C116",
    x"2D2BE66",
    x"2D2BBB7",
    x"2D2B908",
    x"2D2B65B",
    x"2D2B3AD",
    x"2D2B101",
    x"2D2AE55",
    x"2D2ABAA",
    x"2D2A8FF",
    x"2D2A655",
    x"2D2A3AC",
    x"2D2A103",
    x"2D29E5B",
    x"2D29BB4",
    x"2D2990D",
    x"2D29667",
    x"2D293C2",
    x"2D2911E",
    x"2D28E7A",
    x"2D28BD6",
    x"2D28934",
    x"2D28692",
    x"2D283F0",
    x"2D28150",
    x"2D27EB0",
    x"2D27C10",
    x"2D27972",
    x"2D276D4",
    x"2D27436",
    x"2D2719A",
    x"2D26EFE",
    x"2D26C62",
    x"2D269C7",
    x"2D2672D",
    x"2D26494",
    x"2D261FB",
    x"2D25F63",
    x"2D25CCB",
    x"2D25A34",
    x"2D2579E",
    x"2D25509",
    x"2D25274",
    x"2D24FDF",
    x"2D24D4C",
    x"2D24AB9",
    x"2D24826",
    x"2D24595",
    x"2D24304",
    x"2D24073",
    x"2D23DE3",
    x"2D23B54",
    x"2D238C6",
    x"2D23638",
    x"2D233AB",
    x"2D2311E",
    x"2D22E92",
    x"2D22C07",
    x"2D2297C",
    x"2D226F2",
    x"2D22468",
    x"2D221E0",
    x"2D21F58",
    x"2D21CD0",
    x"2D21A49",
    x"2D217C3",
    x"2D2153D",
    x"2D212B8",
    x"2D21034",
    x"2D20DB0",
    x"2D20B2D",
    x"2D208AB",
    x"2D20629",
    x"2D203A7",
    x"2D20127",
    x"2D1FEA7",
    x"2D1FC28",
    x"2D1F9A9",
    x"2D1F72B",
    x"2D1F4AD",
    x"2D1F230",
    x"2D1EFB4",
    x"2D1ED39",
    x"2D1EABE",
    x"2D1E843",
    x"2D1E5C9",
    x"2D1E350",
    x"2D1E0D8",
    x"2D1DE60",
    x"2D1DBE9",
    x"2D1D972",
    x"2D1D6FC",
    x"2D1D486",
    x"2D1D212",
    x"2D1CF9D",
    x"2D1CD2A",
    x"2D1CAB7",
    x"2D1C844",
    x"2D1C5D3",
    x"2D1C361",
    x"2D1C0F1",
    x"2D1BE81",
    x"2D1BC12",
    x"2D1B9A3",
    x"2D1B735",
    x"2D1B4C7",
    x"2D1B25A",
    x"2D1AFEE",
    x"2D1AD83",
    x"2D1AB17",
    x"2D1A8AD",
    x"2D1A643",
    x"2D1A3DA",
    x"2D1A171",
    x"2D19F09",
    x"2D19CA2",
    x"2D19A3B",
    x"2D197D5",
    x"2D1956F",
    x"2D1930A",
    x"2D190A5",
    x"2D18E42",
    x"2D18BDE",
    x"2D1897C",
    x"2D18719",
    x"2D184B8",
    x"2D18257",
    x"2D17FF7",
    x"2D17D97",
    x"2D17B38",
    x"2D178DA",
    x"2D1767C",
    x"2D1741E",
    x"2D171C2",
    x"2D16F65",
    x"2D16D0A",
    x"2D16AAF",
    x"2D16855",
    x"2D165FB",
    x"2D163A2",
    x"2D16149",
    x"2D15EF1",
    x"2D15C99",
    x"2D15A43",
    x"2D157EC",
    x"2D15597",
    x"2D15342",
    x"2D150ED",
    x"2D14E99",
    x"2D14C46",
    x"2D149F3",
    x"2D147A1",
    x"2D1454F",
    x"2D142FE",
    x"2D140AE",
    x"2D13E5E",
    x"2D13C0E",
    x"2D139C0",
    x"2D13772",
    x"2D13524",
    x"2D132D7",
    x"2D1308B",
    x"2D12E3F",
    x"2D12BF3",
    x"2D129A9",
    x"2D1275F",
    x"2D12515",
    x"2D122CC",
    x"2D12084",
    x"2D11E3C",
    x"2D11BF5",
    x"2D119AE",
    x"2D11768",
    x"2D11522",
    x"2D112DD",
    x"2D11099",
    x"2D10E55",
    x"2D10C12",
    x"2D109CF",
    x"2D1078D",
    x"2D1054B",
    x"2D1030A",
    x"2D100C9",
    x"2D0FE8A",
    x"2D0FC4A",
    x"2D0FA0B",
    x"2D0F7CD",
    x"2D0F590",
    x"2D0F352",
    x"2D0F116",
    x"2D0EEDA",
    x"2D0EC9E",
    x"2D0EA64",
    x"2D0E829",
    x"2D0E5EF",
    x"2D0E3B6",
    x"2D0E17E",
    x"2D0DF46",
    x"2D0DD0E",
    x"2D0DAD7",
    x"2D0D8A1",
    x"2D0D66B",
    x"2D0D435",
    x"2D0D201",
    x"2D0CFCC",
    x"2D0CD99",
    x"2D0CB66",
    x"2D0C933",
    x"2D0C701",
    x"2D0C4CF",
    x"2D0C29F",
    x"2D0C06E",
    x"2D0BE3E",
    x"2D0BC0F",
    x"2D0B9E0",
    x"2D0B7B2",
    x"2D0B584",
    x"2D0B357",
    x"2D0B12B",
    x"2D0AEFF",
    x"2D0ACD3",
    x"2D0AAA8",
    x"2D0A87E",
    x"2D0A654",
    x"2D0A42B",
    x"2D0A202",
    x"2D09FDA",
    x"2D09DB2",
    x"2D09B8B",
    x"2D09964",
    x"2D0973E",
    x"2D09519",
    x"2D092F4",
    x"2D090CF",
    x"2D08EAB",
    x"2D08C88",
    x"2D08A65",
    x"2D08843",
    x"2D08621",
    x"2D08400",
    x"2D081DF",
    x"2D07FBF",
    x"2D07D9F",
    x"2D07B80",
    x"2D07961",
    x"2D07743",
    x"2D07526",
    x"2D07309",
    x"2D070EC",
    x"2D06ED0",
    x"2D06CB5",
    x"2D06A9A",
    x"2D0687F",
    x"2D06666",
    x"2D0644C",
    x"2D06233",
    x"2D0601B",
    x"2D05E03",
    x"2D05BEC",
    x"2D059D5",
    x"2D057BF",
    x"2D055A9",
    x"2D05394",
    x"2D05180",
    x"2D04F6C",
    x"2D04D58",
    x"2D04B45",
    x"2D04932",
    x"2D04720",
    x"2D0450F",
    x"2D042FE",
    x"2D040ED",
    x"2D03EDD",
    x"2D03CCE",
    x"2D03ABF",
    x"2D038B0",
    x"2D036A3",
    x"2D03495",
    x"2D03288",
    x"2D0307C",
    x"2D02E70",
    x"2D02C65",
    x"2D02A5A",
    x"2D0284F",
    x"2D02646",
    x"2D0243C",
    x"2D02234",
    x"2D0202B",
    x"2D01E23",
    x"2D01C1C",
    x"2D01A15",
    x"2D0180F",
    x"2D01609",
    x"2D01404",
    x"2D011FF",
    x"2D00FFB",
    x"2D00DF7",
    x"2D00BF4",
    x"2D009F1",
    x"2D007EF",
    x"2D005ED",
    x"2D003EC",
    x"2D001EB",
    x"2CFFFD7",
    x"2CFFBD7",
    x"2CFF7D9",
    x"2CFF3DC",
    x"2CFEFDF",
    x"2CFEBE4",
    x"2CFE7E9",
    x"2CFE3F0",
    x"2CFDFF7",
    x"2CFDC00",
    x"2CFD809",
    x"2CFD414",
    x"2CFD01F",
    x"2CFCC2C",
    x"2CFC839",
    x"2CFC448",
    x"2CFC057",
    x"2CFBC67",
    x"2CFB879",
    x"2CFB48B",
    x"2CFB09E",
    x"2CFACB3",
    x"2CFA8C8",
    x"2CFA4DE",
    x"2CFA0F6",
    x"2CF9D0E",
    x"2CF9927",
    x"2CF9541",
    x"2CF915D",
    x"2CF8D79",
    x"2CF8996",
    x"2CF85B4",
    x"2CF81D3",
    x"2CF7DF3",
    x"2CF7A14",
    x"2CF7636",
    x"2CF7259",
    x"2CF6E7D",
    x"2CF6AA2",
    x"2CF66C7",
    x"2CF62EE",
    x"2CF5F16",
    x"2CF5B3F",
    x"2CF5768",
    x"2CF5393",
    x"2CF4FBF",
    x"2CF4BEB",
    x"2CF4819",
    x"2CF4447",
    x"2CF4076",
    x"2CF3CA7",
    x"2CF38D8",
    x"2CF350A",
    x"2CF313E",
    x"2CF2D72",
    x"2CF29A7",
    x"2CF25DD",
    x"2CF2214",
    x"2CF1E4C",
    x"2CF1A85",
    x"2CF16BF",
    x"2CF12F9",
    x"2CF0F35",
    x"2CF0B72",
    x"2CF07AF",
    x"2CF03EE",
    x"2CF002D",
    x"2CEFC6E",
    x"2CEF8AF",
    x"2CEF4F2",
    x"2CEF135",
    x"2CEED79",
    x"2CEE9BE",
    x"2CEE604",
    x"2CEE24B",
    x"2CEDE93",
    x"2CEDADC",
    x"2CED725",
    x"2CED370",
    x"2CECFBC",
    x"2CECC08",
    x"2CEC856",
    x"2CEC4A4",
    x"2CEC0F3",
    x"2CEBD44",
    x"2CEB995",
    x"2CEB5E7",
    x"2CEB23A",
    x"2CEAE8E",
    x"2CEAAE3",
    x"2CEA738",
    x"2CEA38F",
    x"2CE9FE7",
    x"2CE9C3F",
    x"2CE9898",
    x"2CE94F3",
    x"2CE914E",
    x"2CE8DAA",
    x"2CE8A07",
    x"2CE8665",
    x"2CE82C4",
    x"2CE7F24",
    x"2CE7B84",
    x"2CE77E6",
    x"2CE7448",
    x"2CE70AC",
    x"2CE6D10",
    x"2CE6975",
    x"2CE65DB",
    x"2CE6242",
    x"2CE5EAA",
    x"2CE5B13",
    x"2CE577D",
    x"2CE53E7",
    x"2CE5053",
    x"2CE4CBF",
    x"2CE492C",
    x"2CE459A",
    x"2CE4209",
    x"2CE3E79",
    x"2CE3AEA",
    x"2CE375C",
    x"2CE33CF",
    x"2CE3042",
    x"2CE2CB6",
    x"2CE292C",
    x"2CE25A2",
    x"2CE2219",
    x"2CE1E91",
    x"2CE1B0A",
    x"2CE1783",
    x"2CE13FE",
    x"2CE1079",
    x"2CE0CF6",
    x"2CE0973",
    x"2CE05F1",
    x"2CE0270",
    x"2CDFEF0",
    x"2CDFB70",
    x"2CDF7F2",
    x"2CDF474",
    x"2CDF0F8",
    x"2CDED7C",
    x"2CDEA01",
    x"2CDE687",
    x"2CDE30E",
    x"2CDDF95",
    x"2CDDC1E",
    x"2CDD8A7",
    x"2CDD532",
    x"2CDD1BD",
    x"2CDCE49",
    x"2CDCAD6",
    x"2CDC763",
    x"2CDC3F2",
    x"2CDC081",
    x"2CDBD12",
    x"2CDB9A3",
    x"2CDB635",
    x"2CDB2C8",
    x"2CDAF5B",
    x"2CDABF0",
    x"2CDA885",
    x"2CDA51C",
    x"2CDA1B3",
    x"2CD9E4B",
    x"2CD9AE4",
    x"2CD977D",
    x"2CD9418",
    x"2CD90B3",
    x"2CD8D50",
    x"2CD89ED",
    x"2CD868B",
    x"2CD8329",
    x"2CD7FC9",
    x"2CD7C6A",
    x"2CD790B",
    x"2CD75AD",
    x"2CD7250",
    x"2CD6EF4",
    x"2CD6B99",
    x"2CD683E",
    x"2CD64E4",
    x"2CD618C",
    x"2CD5E34",
    x"2CD5ADD",
    x"2CD5786",
    x"2CD5431",
    x"2CD50DC",
    x"2CD4D88",
    x"2CD4A35",
    x"2CD46E3",
    x"2CD4392",
    x"2CD4041",
    x"2CD3CF2",
    x"2CD39A3",
    x"2CD3655",
    x"2CD3308",
    x"2CD2FBB",
    x"2CD2C70",
    x"2CD2925",
    x"2CD25DB",
    x"2CD2292",
    x"2CD1F4A",
    x"2CD1C03",
    x"2CD18BC",
    x"2CD1576",
    x"2CD1231",
    x"2CD0EED",
    x"2CD0BAA",
    x"2CD0867",
    x"2CD0526",
    x"2CD01E5",
    x"2CCFEA5",
    x"2CCFB65",
    x"2CCF827",
    x"2CCF4E9",
    x"2CCF1AD",
    x"2CCEE71",
    x"2CCEB35",
    x"2CCE7FB",
    x"2CCE4C1",
    x"2CCE189",
    x"2CCDE51",
    x"2CCDB19",
    x"2CCD7E3",
    x"2CCD4AD",
    x"2CCD179",
    x"2CCCE45",
    x"2CCCB12",
    x"2CCC7DF",
    x"2CCC4AE",
    x"2CCC17D",
    x"2CCBE4D",
    x"2CCBB1E",
    x"2CCB7EF",
    x"2CCB4C2",
    x"2CCB195",
    x"2CCAE69",
    x"2CCAB3E",
    x"2CCA813",
    x"2CCA4EA",
    x"2CCA1C1",
    x"2CC9E99",
    x"2CC9B72",
    x"2CC984B",
    x"2CC9525",
    x"2CC9201",
    x"2CC8EDC",
    x"2CC8BB9",
    x"2CC8897",
    x"2CC8575",
    x"2CC8254",
    x"2CC7F34",
    x"2CC7C14",
    x"2CC78F6",
    x"2CC75D8",
    x"2CC72BB",
    x"2CC6F9E",
    x"2CC6C83",
    x"2CC6968",
    x"2CC664E",
    x"2CC6335",
    x"2CC601D",
    x"2CC5D05",
    x"2CC59EE",
    x"2CC56D8",
    x"2CC53C3",
    x"2CC50AE",
    x"2CC4D9A",
    x"2CC4A87",
    x"2CC4775",
    x"2CC4464",
    x"2CC4153",
    x"2CC3E43",
    x"2CC3B34",
    x"2CC3825",
    x"2CC3518",
    x"2CC320B",
    x"2CC2EFF",
    x"2CC2BF3",
    x"2CC28E9",
    x"2CC25DF",
    x"2CC22D6",
    x"2CC1FCD",
    x"2CC1CC6",
    x"2CC19BF",
    x"2CC16B9",
    x"2CC13B4",
    x"2CC10AF",
    x"2CC0DAB",
    x"2CC0AA8",
    x"2CC07A6",
    x"2CC04A4",
    x"2CC01A4",
    x"2CBFEA4",
    x"2CBFBA4",
    x"2CBF8A6",
    x"2CBF5A8",
    x"2CBF2AB",
    x"2CBEFAF",
    x"2CBECB3",
    x"2CBE9B8",
    x"2CBE6BE",
    x"2CBE3C5",
    x"2CBE0CC",
    x"2CBDDD4",
    x"2CBDADD",
    x"2CBD7E7",
    x"2CBD4F1",
    x"2CBD1FD",
    x"2CBCF08",
    x"2CBCC15",
    x"2CBC922",
    x"2CBC631",
    x"2CBC33F",
    x"2CBC04F",
    x"2CBBD5F",
    x"2CBBA70",
    x"2CBB782",
    x"2CBB494",
    x"2CBB1A8",
    x"2CBAEBC",
    x"2CBABD0",
    x"2CBA8E6",
    x"2CBA5FC",
    x"2CBA313",
    x"2CBA02A",
    x"2CB9D43",
    x"2CB9A5C",
    x"2CB9775",
    x"2CB9490",
    x"2CB91AB",
    x"2CB8EC7",
    x"2CB8BE4",
    x"2CB8901",
    x"2CB861F",
    x"2CB833E",
    x"2CB805E",
    x"2CB7D7E",
    x"2CB7A9F",
    x"2CB77C1",
    x"2CB74E3",
    x"2CB7206",
    x"2CB6F2A",
    x"2CB6C4F",
    x"2CB6974",
    x"2CB669A",
    x"2CB63C1",
    x"2CB60E8",
    x"2CB5E10",
    x"2CB5B39",
    x"2CB5862",
    x"2CB558D",
    x"2CB52B8",
    x"2CB4FE3",
    x"2CB4D10",
    x"2CB4A3D",
    x"2CB476B",
    x"2CB4499",
    x"2CB41C8",
    x"2CB3EF8",
    x"2CB3C29",
    x"2CB395A",
    x"2CB368C",
    x"2CB33BF",
    x"2CB30F2",
    x"2CB2E26",
    x"2CB2B5B",
    x"2CB2891",
    x"2CB25C7",
    x"2CB22FE",
    x"2CB2035",
    x"2CB1D6E",
    x"2CB1AA7",
    x"2CB17E0",
    x"2CB151B",
    x"2CB1256",
    x"2CB0F92",
    x"2CB0CCE",
    x"2CB0A0B",
    x"2CB0749",
    x"2CB0488",
    x"2CB01C7",
    x"2CAFF07",
    x"2CAFC47",
    x"2CAF989",
    x"2CAF6CB",
    x"2CAF40D",
    x"2CAF150",
    x"2CAEE94",
    x"2CAEBD9",
    x"2CAE91F",
    x"2CAE665",
    x"2CAE3AB",
    x"2CAE0F3",
    x"2CADE3B",
    x"2CADB84",
    x"2CAD8CD",
    x"2CAD617",
    x"2CAD362",
    x"2CAD0AE",
    x"2CACDFA",
    x"2CACB47",
    x"2CAC894",
    x"2CAC5E2",
    x"2CAC331",
    x"2CAC081",
    x"2CABDD1",
    x"2CABB22",
    x"2CAB873",
    x"2CAB5C6",
    x"2CAB318",
    x"2CAB06C",
    x"2CAADC0",
    x"2CAAB15",
    x"2CAA86B",
    x"2CAA5C1",
    x"2CAA318",
    x"2CAA06F",
    x"2CA9DC8",
    x"2CA9B20",
    x"2CA987A",
    x"2CA95D4",
    x"2CA932F",
    x"2CA908B",
    x"2CA8DE7",
    x"2CA8B44",
    x"2CA88A1",
    x"2CA85FF",
    x"2CA835E",
    x"2CA80BE",
    x"2CA7E1E",
    x"2CA7B7F",
    x"2CA78E0",
    x"2CA7642",
    x"2CA73A5",
    x"2CA7108",
    x"2CA6E6C",
    x"2CA6BD1",
    x"2CA6937",
    x"2CA669D",
    x"2CA6403",
    x"2CA616B",
    x"2CA5ED3",
    x"2CA5C3B",
    x"2CA59A4",
    x"2CA570E",
    x"2CA5479",
    x"2CA51E4",
    x"2CA4F50",
    x"2CA4CBC",
    x"2CA4A2A",
    x"2CA4797",
    x"2CA4506",
    x"2CA4275",
    x"2CA3FE5",
    x"2CA3D55",
    x"2CA3AC6",
    x"2CA3838",
    x"2CA35AA",
    x"2CA331D",
    x"2CA3090",
    x"2CA2E04",
    x"2CA2B79",
    x"2CA28EF",
    x"2CA2665",
    x"2CA23DB",
    x"2CA2153",
    x"2CA1ECB",
    x"2CA1C43",
    x"2CA19BD",
    x"2CA1737",
    x"2CA14B1",
    x"2CA122C",
    x"2CA0FA8",
    x"2CA0D24",
    x"2CA0AA1",
    x"2CA081F",
    x"2CA059D",
    x"2CA031C",
    x"2CA009C",
    x"2C9FE1C",
    x"2C9FB9D",
    x"2C9F91E",
    x"2C9F6A0",
    x"2C9F423",
    x"2C9F1A6",
    x"2C9EF2A",
    x"2C9ECAF",
    x"2C9EA34",
    x"2C9E7B9",
    x"2C9E540",
    x"2C9E2C7",
    x"2C9E04E",
    x"2C9DDD7",
    x"2C9DB5F",
    x"2C9D8E9",
    x"2C9D673",
    x"2C9D3FE",
    x"2C9D189",
    x"2C9CF15",
    x"2C9CCA1",
    x"2C9CA2F",
    x"2C9C7BC",
    x"2C9C54B",
    x"2C9C2DA",
    x"2C9C069",
    x"2C9BDFA",
    x"2C9BB8A",
    x"2C9B91C",
    x"2C9B6AE",
    x"2C9B440",
    x"2C9B1D4",
    x"2C9AF68",
    x"2C9ACFC",
    x"2C9AA91",
    x"2C9A827",
    x"2C9A5BD",
    x"2C9A354",
    x"2C9A0EB",
    x"2C99E83",
    x"2C99C1C",
    x"2C999B5",
    x"2C9974F",
    x"2C994EA",
    x"2C99285",
    x"2C99020",
    x"2C98DBD",
    x"2C98B59",
    x"2C988F7",
    x"2C98695",
    x"2C98434",
    x"2C981D3",
    x"2C97F73",
    x"2C97D13",
    x"2C97AB4",
    x"2C97856",
    x"2C975F8",
    x"2C9739B",
    x"2C9713E",
    x"2C96EE2",
    x"2C96C87",
    x"2C96A2C",
    x"2C967D2",
    x"2C96578",
    x"2C9631F",
    x"2C960C6",
    x"2C95E6F",
    x"2C95C17",
    x"2C959C1",
    x"2C9576A",
    x"2C95515",
    x"2C952C0",
    x"2C9506B",
    x"2C94E18",
    x"2C94BC4",
    x"2C94972",
    x"2C94720",
    x"2C944CE",
    x"2C9427D",
    x"2C9402D",
    x"2C93DDD",
    x"2C93B8E",
    x"2C9393F",
    x"2C936F1",
    x"2C934A4",
    x"2C93257",
    x"2C9300B",
    x"2C92DBF",
    x"2C92B74",
    x"2C92929",
    x"2C926DF",
    x"2C92496",
    x"2C9224D",
    x"2C92005",
    x"2C91DBD",
    x"2C91B76",
    x"2C9192F",
    x"2C916E9",
    x"2C914A4",
    x"2C9125F",
    x"2C9101B",
    x"2C90DD7",
    x"2C90B94",
    x"2C90951",
    x"2C9070F",
    x"2C904CE",
    x"2C9028D",
    x"2C9004C",
    x"2C8FE0D",
    x"2C8FBCD",
    x"2C8F98F",
    x"2C8F750",
    x"2C8F513",
    x"2C8F2D6",
    x"2C8F09A",
    x"2C8EE5E",
    x"2C8EC22",
    x"2C8E9E8",
    x"2C8E7AD",
    x"2C8E574",
    x"2C8E33B",
    x"2C8E102",
    x"2C8DECA",
    x"2C8DC93",
    x"2C8DA5C",
    x"2C8D826",
    x"2C8D5F0",
    x"2C8D3BB",
    x"2C8D186",
    x"2C8CF52",
    x"2C8CD1E",
    x"2C8CAEB",
    x"2C8C8B9",
    x"2C8C687",
    x"2C8C456",
    x"2C8C225",
    x"2C8BFF4",
    x"2C8BDC5",
    x"2C8BB96",
    x"2C8B967",
    x"2C8B739",
    x"2C8B50B",
    x"2C8B2DE",
    x"2C8B0B2",
    x"2C8AE86",
    x"2C8AC5B",
    x"2C8AA30",
    x"2C8A806",
    x"2C8A5DC",
    x"2C8A3B3",
    x"2C8A18A",
    x"2C89F62",
    x"2C89D3A",
    x"2C89B13",
    x"2C898ED",
    x"2C896C7",
    x"2C894A1",
    x"2C8927C",
    x"2C89058",
    x"2C88E34",
    x"2C88C11",
    x"2C889EE",
    x"2C887CC",
    x"2C885AA",
    x"2C88389",
    x"2C88169",
    x"2C87F48",
    x"2C87D29",
    x"2C87B0A",
    x"2C878EB",
    x"2C876CD",
    x"2C874B0",
    x"2C87293",
    x"2C87077",
    x"2C86E5B",
    x"2C86C40",
    x"2C86A25",
    x"2C8680A",
    x"2C865F1",
    x"2C863D8",
    x"2C861BF",
    x"2C85FA7",
    x"2C85D8F",
    x"2C85B78",
    x"2C85961",
    x"2C8574B",
    x"2C85536",
    x"2C85321",
    x"2C8510C",
    x"2C84EF8",
    x"2C84CE5",
    x"2C84AD2",
    x"2C848BF",
    x"2C846AD",
    x"2C8449C",
    x"2C8428B",
    x"2C8407B",
    x"2C83E6B",
    x"2C83C5B",
    x"2C83A4C",
    x"2C8383E",
    x"2C83630",
    x"2C83423",
    x"2C83216",
    x"2C8300A",
    x"2C82DFE",
    x"2C82BF3",
    x"2C829E8",
    x"2C827DE",
    x"2C825D4",
    x"2C823CB",
    x"2C821C2",
    x"2C81FBA",
    x"2C81DB3",
    x"2C81BAB",
    x"2C819A5",
    x"2C8179F",
    x"2C81599",
    x"2C81394",
    x"2C8118F",
    x"2C80F8B",
    x"2C80D87",
    x"2C80B84",
    x"2C80982",
    x"2C80780",
    x"2C8057E",
    x"2C8037D",
    x"2C8017C",
    x"2C7FEF8",
    x"2C7FAF9",
    x"2C7F6FB",
    x"2C7F2FE",
    x"2C7EF02",
    x"2C7EB06",
    x"2C7E70C",
    x"2C7E313",
    x"2C7DF1A",
    x"2C7DB23",
    x"2C7D72D",
    x"2C7D338",
    x"2C7CF43",
    x"2C7CB50",
    x"2C7C75E",
    x"2C7C36C",
    x"2C7BF7C",
    x"2C7BB8D",
    x"2C7B79E",
    x"2C7B3B1",
    x"2C7AFC4",
    x"2C7ABD9",
    x"2C7A7EE",
    x"2C7A405",
    x"2C7A01C",
    x"2C79C35",
    x"2C7984E",
    x"2C79469",
    x"2C79084",
    x"2C78CA0",
    x"2C788BE",
    x"2C784DC",
    x"2C780FB",
    x"2C77D1C",
    x"2C7793D",
    x"2C7755F",
    x"2C77182",
    x"2C76DA6",
    x"2C769CB",
    x"2C765F1",
    x"2C76218",
    x"2C75E40",
    x"2C75A69",
    x"2C75693",
    x"2C752BE",
    x"2C74EEA",
    x"2C74B16",
    x"2C74744",
    x"2C74373",
    x"2C73FA2",
    x"2C73BD3",
    x"2C73804",
    x"2C73437",
    x"2C7306A",
    x"2C72C9F",
    x"2C728D4",
    x"2C7250A",
    x"2C72142",
    x"2C71D7A",
    x"2C719B3",
    x"2C715ED",
    x"2C71228",
    x"2C70E64",
    x"2C70AA1",
    x"2C706DE",
    x"2C7031D",
    x"2C6FF5D",
    x"2C6FB9D",
    x"2C6F7DF",
    x"2C6F422",
    x"2C6F065",
    x"2C6ECA9",
    x"2C6E8EF",
    x"2C6E535",
    x"2C6E17C",
    x"2C6DDC4",
    x"2C6DA0D",
    x"2C6D657",
    x"2C6D2A2",
    x"2C6CEEE",
    x"2C6CB3B",
    x"2C6C788",
    x"2C6C3D7",
    x"2C6C026",
    x"2C6BC77",
    x"2C6B8C8",
    x"2C6B51A",
    x"2C6B16D",
    x"2C6ADC2",
    x"2C6AA17",
    x"2C6A66D",
    x"2C6A2C3",
    x"2C69F1B",
    x"2C69B74",
    x"2C697CD",
    x"2C69428",
    x"2C69083",
    x"2C68CE0",
    x"2C6893D",
    x"2C6859B",
    x"2C681FA",
    x"2C67E5A",
    x"2C67ABB",
    x"2C6771D",
    x"2C6737F",
    x"2C66FE3",
    x"2C66C47",
    x"2C668AD",
    x"2C66513",
    x"2C6617A",
    x"2C65DE2",
    x"2C65A4B",
    x"2C656B5",
    x"2C65320",
    x"2C64F8C",
    x"2C64BF8",
    x"2C64866",
    x"2C644D4",
    x"2C64143",
    x"2C63DB3",
    x"2C63A24",
    x"2C63696",
    x"2C63309",
    x"2C62F7D",
    x"2C62BF1",
    x"2C62867",
    x"2C624DD",
    x"2C62154",
    x"2C61DCC",
    x"2C61A45",
    x"2C616BF",
    x"2C6133A",
    x"2C60FB6",
    x"2C60C32",
    x"2C608B0",
    x"2C6052E",
    x"2C601AD",
    x"2C5FE2D",
    x"2C5FAAE",
    x"2C5F730",
    x"2C5F3B2",
    x"2C5F036",
    x"2C5ECBA",
    x"2C5E93F",
    x"2C5E5C6",
    x"2C5E24D",
    x"2C5DED4",
    x"2C5DB5D",
    x"2C5D7E7",
    x"2C5D471",
    x"2C5D0FD",
    x"2C5CD89",
    x"2C5CA16",
    x"2C5C6A4",
    x"2C5C332",
    x"2C5BFC2",
    x"2C5BC53",
    x"2C5B8E4",
    x"2C5B576",
    x"2C5B209",
    x"2C5AE9D",
    x"2C5AB32",
    x"2C5A7C8",
    x"2C5A45E",
    x"2C5A0F5",
    x"2C59D8E",
    x"2C59A27",
    x"2C596C0",
    x"2C5935B",
    x"2C58FF7",
    x"2C58C93",
    x"2C58930",
    x"2C585CF",
    x"2C5826E",
    x"2C57F0D",
    x"2C57BAE",
    x"2C57850",
    x"2C574F2",
    x"2C57195",
    x"2C56E39",
    x"2C56ADE",
    x"2C56784",
    x"2C5642A",
    x"2C560D2",
    x"2C55D7A",
    x"2C55A23",
    x"2C556CD",
    x"2C55377",
    x"2C55023",
    x"2C54CCF",
    x"2C5497D",
    x"2C5462B",
    x"2C542D9",
    x"2C53F89",
    x"2C53C3A",
    x"2C538EB",
    x"2C5359D",
    x"2C53250",
    x"2C52F04",
    x"2C52BB9",
    x"2C5286E",
    x"2C52525",
    x"2C521DC",
    x"2C51E94",
    x"2C51B4C",
    x"2C51806",
    x"2C514C0",
    x"2C5117C",
    x"2C50E38",
    x"2C50AF4",
    x"2C507B2",
    x"2C50471",
    x"2C50130",
    x"2C4FDF0",
    x"2C4FAB1",
    x"2C4F773",
    x"2C4F435",
    x"2C4F0F9",
    x"2C4EDBD",
    x"2C4EA82",
    x"2C4E747",
    x"2C4E40E",
    x"2C4E0D5",
    x"2C4DD9E",
    x"2C4DA67",
    x"2C4D730",
    x"2C4D3FB",
    x"2C4D0C6",
    x"2C4CD93",
    x"2C4CA60",
    x"2C4C72D",
    x"2C4C3FC",
    x"2C4C0CB",
    x"2C4BD9C",
    x"2C4BA6D",
    x"2C4B73E",
    x"2C4B411",
    x"2C4B0E4",
    x"2C4ADB9",
    x"2C4AA8E",
    x"2C4A763",
    x"2C4A43A",
    x"2C4A111",
    x"2C49DE9",
    x"2C49AC2",
    x"2C4979C",
    x"2C49476",
    x"2C49152",
    x"2C48E2E",
    x"2C48B0B",
    x"2C487E8",
    x"2C484C7",
    x"2C481A6",
    x"2C47E86",
    x"2C47B67",
    x"2C47848",
    x"2C4752A",
    x"2C4720E",
    x"2C46EF1",
    x"2C46BD6",
    x"2C468BC",
    x"2C465A2",
    x"2C46289",
    x"2C45F70",
    x"2C45C59",
    x"2C45942",
    x"2C4562C",
    x"2C45317",
    x"2C45003",
    x"2C44CEF",
    x"2C449DC",
    x"2C446CA",
    x"2C443B9",
    x"2C440A8",
    x"2C43D99",
    x"2C43A8A",
    x"2C4377B",
    x"2C4346E",
    x"2C43161",
    x"2C42E55",
    x"2C42B4A",
    x"2C42840",
    x"2C42536",
    x"2C4222D",
    x"2C41F25",
    x"2C41C1D",
    x"2C41917",
    x"2C41611",
    x"2C4130C",
    x"2C41007",
    x"2C40D04",
    x"2C40A01",
    x"2C406FF",
    x"2C403FD",
    x"2C400FD",
    x"2C3FDFD",
    x"2C3FAFE",
    x"2C3F7FF",
    x"2C3F502",
    x"2C3F205",
    x"2C3EF09",
    x"2C3EC0D",
    x"2C3E913",
    x"2C3E619",
    x"2C3E320",
    x"2C3E027",
    x"2C3DD2F",
    x"2C3DA39",
    x"2C3D742",
    x"2C3D44D",
    x"2C3D158",
    x"2C3CE64",
    x"2C3CB71",
    x"2C3C87F",
    x"2C3C58D",
    x"2C3C29C",
    x"2C3BFAB",
    x"2C3BCBC",
    x"2C3B9CD",
    x"2C3B6DF",
    x"2C3B3F2",
    x"2C3B105",
    x"2C3AE19",
    x"2C3AB2E",
    x"2C3A844",
    x"2C3A55A",
    x"2C3A271",
    x"2C39F89",
    x"2C39CA1",
    x"2C399BA",
    x"2C396D4",
    x"2C393EF",
    x"2C3910A",
    x"2C38E26",
    x"2C38B43",
    x"2C38861",
    x"2C3857F",
    x"2C3829E",
    x"2C37FBE",
    x"2C37CDE",
    x"2C379FF",
    x"2C37721",
    x"2C37444",
    x"2C37167",
    x"2C36E8B",
    x"2C36BB0",
    x"2C368D5",
    x"2C365FB",
    x"2C36322",
    x"2C3604A",
    x"2C35D72",
    x"2C35A9B",
    x"2C357C5",
    x"2C354EF",
    x"2C3521A",
    x"2C34F46",
    x"2C34C73",
    x"2C349A0",
    x"2C346CE",
    x"2C343FC",
    x"2C3412C",
    x"2C33E5C",
    x"2C33B8D",
    x"2C338BE",
    x"2C335F0",
    x"2C33323",
    x"2C33057",
    x"2C32D8B",
    x"2C32AC0",
    x"2C327F6",
    x"2C3252C",
    x"2C32263",
    x"2C31F9B",
    x"2C31CD3",
    x"2C31A0C",
    x"2C31746",
    x"2C31481",
    x"2C311BC",
    x"2C30EF8",
    x"2C30C34",
    x"2C30972",
    x"2C306B0",
    x"2C303EE",
    x"2C3012E",
    x"2C2FE6E",
    x"2C2FBAF",
    x"2C2F8F0",
    x"2C2F632",
    x"2C2F375",
    x"2C2F0B8",
    x"2C2EDFC",
    x"2C2EB41",
    x"2C2E887",
    x"2C2E5CD",
    x"2C2E314",
    x"2C2E05C",
    x"2C2DDA4",
    x"2C2DAED",
    x"2C2D836",
    x"2C2D581",
    x"2C2D2CC",
    x"2C2D017",
    x"2C2CD64",
    x"2C2CAB1",
    x"2C2C7FE",
    x"2C2C54D",
    x"2C2C29C",
    x"2C2BFEB",
    x"2C2BD3C",
    x"2C2BA8D",
    x"2C2B7DE",
    x"2C2B531",
    x"2C2B284",
    x"2C2AFD7",
    x"2C2AD2C",
    x"2C2AA81",
    x"2C2A7D7",
    x"2C2A52D",
    x"2C2A284",
    x"2C29FDC",
    x"2C29D34",
    x"2C29A8D",
    x"2C297E7",
    x"2C29541",
    x"2C2929C",
    x"2C28FF8",
    x"2C28D54",
    x"2C28AB1",
    x"2C2880F",
    x"2C2856D",
    x"2C282CC",
    x"2C2802C",
    x"2C27D8C",
    x"2C27AED",
    x"2C2784E",
    x"2C275B1",
    x"2C27314",
    x"2C27077",
    x"2C26DDB",
    x"2C26B40",
    x"2C268A6",
    x"2C2660C",
    x"2C26373",
    x"2C260DA",
    x"2C25E42",
    x"2C25BAB",
    x"2C25914",
    x"2C2567F",
    x"2C253E9",
    x"2C25155",
    x"2C24EC1",
    x"2C24C2D",
    x"2C2499A",
    x"2C24708",
    x"2C24477",
    x"2C241E6",
    x"2C23F56",
    x"2C23CC7",
    x"2C23A38",
    x"2C237A9",
    x"2C2351C",
    x"2C2328F",
    x"2C23003",
    x"2C22D77",
    x"2C22AEC",
    x"2C22861",
    x"2C225D8",
    x"2C2234E",
    x"2C220C6",
    x"2C21E3E",
    x"2C21BB7",
    x"2C21930",
    x"2C216AA",
    x"2C21425",
    x"2C211A0",
    x"2C20F1C",
    x"2C20C99",
    x"2C20A16",
    x"2C20794",
    x"2C20512",
    x"2C20291",
    x"2C20011",
    x"2C1FD91",
    x"2C1FB12",
    x"2C1F893",
    x"2C1F616",
    x"2C1F398",
    x"2C1F11C",
    x"2C1EEA0",
    x"2C1EC25",
    x"2C1E9AA",
    x"2C1E730",
    x"2C1E4B6",
    x"2C1E23D",
    x"2C1DFC5",
    x"2C1DD4D",
    x"2C1DAD6",
    x"2C1D860",
    x"2C1D5EA",
    x"2C1D375",
    x"2C1D100",
    x"2C1CE8D",
    x"2C1CC19",
    x"2C1C9A6",
    x"2C1C734",
    x"2C1C4C3",
    x"2C1C252",
    x"2C1BFE2",
    x"2C1BD72",
    x"2C1BB03",
    x"2C1B895",
    x"2C1B627",
    x"2C1B3B9",
    x"2C1B14D",
    x"2C1AEE1",
    x"2C1AC75",
    x"2C1AA0B",
    x"2C1A7A0",
    x"2C1A537",
    x"2C1A2CE",
    x"2C1A065",
    x"2C19DFE",
    x"2C19B96",
    x"2C19930",
    x"2C196CA",
    x"2C19464",
    x"2C19200",
    x"2C18F9B",
    x"2C18D38",
    x"2C18AD5",
    x"2C18872",
    x"2C18611",
    x"2C183AF",
    x"2C1814F",
    x"2C17EEF",
    x"2C17C8F",
    x"2C17A30",
    x"2C177D2",
    x"2C17574",
    x"2C17317",
    x"2C170BB",
    x"2C16E5F",
    x"2C16C04",
    x"2C169A9",
    x"2C1674F",
    x"2C164F5",
    x"2C1629C",
    x"2C16044",
    x"2C15DEC",
    x"2C15B95",
    x"2C1593F",
    x"2C156E9",
    x"2C15493",
    x"2C1523E",
    x"2C14FEA",
    x"2C14D96",
    x"2C14B43",
    x"2C148F1",
    x"2C1469F",
    x"2C1444D",
    x"2C141FD",
    x"2C13FAC",
    x"2C13D5D",
    x"2C13B0E",
    x"2C138BF",
    x"2C13671",
    x"2C13424",
    x"2C131D7",
    x"2C12F8B",
    x"2C12D3F",
    x"2C12AF4",
    x"2C128AA",
    x"2C12660",
    x"2C12417",
    x"2C121CE",
    x"2C11F86",
    x"2C11D3E",
    x"2C11AF7",
    x"2C118B1",
    x"2C1166B",
    x"2C11426",
    x"2C111E1",
    x"2C10F9D",
    x"2C10D59",
    x"2C10B16",
    x"2C108D3",
    x"2C10692",
    x"2C10450",
    x"2C1020F",
    x"2C0FFCF",
    x"2C0FD8F",
    x"2C0FB50",
    x"2C0F912",
    x"2C0F6D4",
    x"2C0F496",
    x"2C0F25A",
    x"2C0F01D",
    x"2C0EDE1",
    x"2C0EBA6",
    x"2C0E96C",
    x"2C0E732",
    x"2C0E4F8",
    x"2C0E2BF",
    x"2C0E087",
    x"2C0DE4F",
    x"2C0DC18",
    x"2C0D9E1",
    x"2C0D7AB",
    x"2C0D575",
    x"2C0D340",
    x"2C0D10B",
    x"2C0CED7",
    x"2C0CCA4",
    x"2C0CA71",
    x"2C0C83F",
    x"2C0C60D",
    x"2C0C3DC",
    x"2C0C1AB",
    x"2C0BF7B",
    x"2C0BD4B",
    x"2C0BB1C",
    x"2C0B8EE",
    x"2C0B6C0",
    x"2C0B492",
    x"2C0B265",
    x"2C0B039",
    x"2C0AE0D",
    x"2C0ABE2",
    x"2C0A9B7",
    x"2C0A78D",
    x"2C0A564",
    x"2C0A33A",
    x"2C0A112",
    x"2C09EEA",
    x"2C09CC2",
    x"2C09A9C",
    x"2C09875",
    x"2C0964F",
    x"2C0942A",
    x"2C09205",
    x"2C08FE1",
    x"2C08DBD",
    x"2C08B9A",
    x"2C08978",
    x"2C08755",
    x"2C08534",
    x"2C08313",
    x"2C080F2",
    x"2C07ED2",
    x"2C07CB3",
    x"2C07A94",
    x"2C07876",
    x"2C07658",
    x"2C0743A",
    x"2C0721E",
    x"2C07001",
    x"2C06DE6",
    x"2C06BCA",
    x"2C069B0",
    x"2C06796",
    x"2C0657C",
    x"2C06363",
    x"2C0614A",
    x"2C05F32",
    x"2C05D1B",
    x"2C05B04",
    x"2C058ED",
    x"2C056D7",
    x"2C054C2",
    x"2C052AD",
    x"2C05098",
    x"2C04E84",
    x"2C04C71",
    x"2C04A5E",
    x"2C0484C",
    x"2C0463A",
    x"2C04429",
    x"2C04218",
    x"2C04008",
    x"2C03DF8",
    x"2C03BE9",
    x"2C039DA",
    x"2C037CC",
    x"2C035BE",
    x"2C033B1",
    x"2C031A4",
    x"2C02F98",
    x"2C02D8D",
    x"2C02B81",
    x"2C02977",
    x"2C0276D",
    x"2C02563",
    x"2C0235A",
    x"2C02151",
    x"2C01F49",
    x"2C01D42",
    x"2C01B3B",
    x"2C01934",
    x"2C0172E",
    x"2C01529",
    x"2C01323",
    x"2C0111F",
    x"2C00F1B",
    x"2C00D17",
    x"2C00B14",
    x"2C00912",
    x"2C00710",
    x"2C0050E",
    x"2C0030D",
    x"2C0010D",
    x"2BFFE1A",
    x"2BFFA1B",
    x"2BFF61D",
    x"2BFF220",
    x"2BFEE24",
    x"2BFEA29",
    x"2BFE62F",
    x"2BFE236",
    x"2BFDE3E",
    x"2BFDA47",
    x"2BFD651",
    x"2BFD25C",
    x"2BFCE67",
    x"2BFCA74",
    x"2BFC682",
    x"2BFC291",
    x"2BFBEA1",
    x"2BFBAB2",
    x"2BFB6C4",
    x"2BFB2D6",
    x"2BFAEEA",
    x"2BFAAFF",
    x"2BFA715",
    x"2BFA32B",
    x"2BF9F43",
    x"2BF9B5C",
    x"2BF9775",
    x"2BF9390",
    x"2BF8FAC",
    x"2BF8BC8",
    x"2BF87E6",
    x"2BF8404",
    x"2BF8024",
    x"2BF7C44",
    x"2BF7866",
    x"2BF7488",
    x"2BF70AB",
    x"2BF6CD0",
    x"2BF68F5",
    x"2BF651B",
    x"2BF6142",
    x"2BF5D6B",
    x"2BF5994",
    x"2BF55BE",
    x"2BF51E9",
    x"2BF4E15",
    x"2BF4A42",
    x"2BF4670",
    x"2BF429F",
    x"2BF3ECE",
    x"2BF3AFF",
    x"2BF3731",
    x"2BF3364",
    x"2BF2F97",
    x"2BF2BCC",
    x"2BF2801",
    x"2BF2438",
    x"2BF206F",
    x"2BF1CA7",
    x"2BF18E1",
    x"2BF151B",
    x"2BF1156",
    x"2BF0D92",
    x"2BF09CF",
    x"2BF060D",
    x"2BF024C",
    x"2BEFE8C",
    x"2BEFACD",
    x"2BEF70F",
    x"2BEF352",
    x"2BEEF95",
    x"2BEEBDA",
    x"2BEE81F",
    x"2BEE466",
    x"2BEE0AD",
    x"2BEDCF5",
    x"2BED93F",
    x"2BED589",
    x"2BED1D4",
    x"2BECE20",
    x"2BECA6D",
    x"2BEC6BB",
    x"2BEC309",
    x"2BEBF59",
    x"2BEBBAA",
    x"2BEB7FB",
    x"2BEB44E",
    x"2BEB0A1",
    x"2BEACF5",
    x"2BEA94B",
    x"2BEA5A1",
    x"2BEA1F8",
    x"2BE9E50",
    x"2BE9AA9",
    x"2BE9703",
    x"2BE935D",
    x"2BE8FB9",
    x"2BE8C15",
    x"2BE8873",
    x"2BE84D1",
    x"2BE8130",
    x"2BE7D91",
    x"2BE79F2",
    x"2BE7654",
    x"2BE72B6",
    x"2BE6F1A",
    x"2BE6B7F",
    x"2BE67E4",
    x"2BE644B",
    x"2BE60B2",
    x"2BE5D1B",
    x"2BE5984",
    x"2BE55EE",
    x"2BE5259",
    x"2BE4EC5",
    x"2BE4B31",
    x"2BE479F",
    x"2BE440E",
    x"2BE407D",
    x"2BE3CED",
    x"2BE395F",
    x"2BE35D1",
    x"2BE3244",
    x"2BE2EB8",
    x"2BE2B2C",
    x"2BE27A2",
    x"2BE2418",
    x"2BE2090",
    x"2BE1D08",
    x"2BE1981",
    x"2BE15FB",
    x"2BE1276",
    x"2BE0EF2",
    x"2BE0B6F",
    x"2BE07EC",
    x"2BE046B",
    x"2BE00EA",
    x"2BDFD6A",
    x"2BDF9EC",
    x"2BDF66E",
    x"2BDF2F0",
    x"2BDEF74",
    x"2BDEBF9",
    x"2BDE87E",
    x"2BDE504",
    x"2BDE18C",
    x"2BDDE14",
    x"2BDDA9D",
    x"2BDD726",
    x"2BDD3B1",
    x"2BDD03C",
    x"2BDCCC9",
    x"2BDC956",
    x"2BDC5E4",
    x"2BDC273",
    x"2BDBF03",
    x"2BDBB94",
    x"2BDB825",
    x"2BDB4B8",
    x"2BDB14B",
    x"2BDADDF",
    x"2BDAA74",
    x"2BDA70A",
    x"2BDA3A0",
    x"2BDA038",
    x"2BD9CD0",
    x"2BD9969",
    x"2BD9603",
    x"2BD929E",
    x"2BD8F3A",
    x"2BD8BD7",
    x"2BD8874",
    x"2BD8513",
    x"2BD81B2",
    x"2BD7E52",
    x"2BD7AF3",
    x"2BD7794",
    x"2BD7437",
    x"2BD70DA",
    x"2BD6D7E",
    x"2BD6A23",
    x"2BD66C9",
    x"2BD6370",
    x"2BD6018",
    x"2BD5CC0",
    x"2BD5969",
    x"2BD5613",
    x"2BD52BE",
    x"2BD4F6A",
    x"2BD4C16",
    x"2BD48C4",
    x"2BD4572",
    x"2BD4221",
    x"2BD3ED1",
    x"2BD3B82",
    x"2BD3833",
    x"2BD34E6",
    x"2BD3199",
    x"2BD2E4D",
    x"2BD2B02",
    x"2BD27B7",
    x"2BD246E",
    x"2BD2125",
    x"2BD1DDD",
    x"2BD1A96",
    x"2BD1750",
    x"2BD140A",
    x"2BD10C6",
    x"2BD0D82",
    x"2BD0A3F",
    x"2BD06FD",
    x"2BD03BC",
    x"2BD007B",
    x"2BCFD3B",
    x"2BCF9FC",
    x"2BCF6BE",
    x"2BCF381",
    x"2BCF045",
    x"2BCED09",
    x"2BCE9CE",
    x"2BCE694",
    x"2BCE35B",
    x"2BCE022",
    x"2BCDCEB",
    x"2BCD9B4",
    x"2BCD67E",
    x"2BCD349",
    x"2BCD014",
    x"2BCCCE1",
    x"2BCC9AE",
    x"2BCC67C",
    x"2BCC34B",
    x"2BCC01A",
    x"2BCBCEB",
    x"2BCB9BC",
    x"2BCB68E",
    x"2BCB360",
    x"2BCB034",
    x"2BCAD08",
    x"2BCA9DD",
    x"2BCA6B3",
    x"2BCA38A",
    x"2BCA062",
    x"2BC9D3A",
    x"2BC9A13",
    x"2BC96ED",
    x"2BC93C8",
    x"2BC90A3",
    x"2BC8D7F",
    x"2BC8A5C",
    x"2BC873A",
    x"2BC8419",
    x"2BC80F8",
    x"2BC7DD8",
    x"2BC7AB9",
    x"2BC779B",
    x"2BC747D",
    x"2BC7161",
    x"2BC6E45",
    x"2BC6B29",
    x"2BC680F",
    x"2BC64F5",
    x"2BC61DD",
    x"2BC5EC4",
    x"2BC5BAD",
    x"2BC5897",
    x"2BC5581",
    x"2BC526C",
    x"2BC4F58",
    x"2BC4C44",
    x"2BC4931",
    x"2BC4620",
    x"2BC430E",
    x"2BC3FFE",
    x"2BC3CEE",
    x"2BC39E0",
    x"2BC36D1",
    x"2BC33C4",
    x"2BC30B8",
    x"2BC2DAC",
    x"2BC2AA1",
    x"2BC2796",
    x"2BC248D",
    x"2BC2184",
    x"2BC1E7C",
    x"2BC1B75",
    x"2BC186E",
    x"2BC1569",
    x"2BC1264",
    x"2BC0F60",
    x"2BC0C5C",
    x"2BC0959",
    x"2BC0657",
    x"2BC0356",
    x"2BC0056",
    x"2BBFD56",
    x"2BBFA57",
    x"2BBF759",
    x"2BBF45B",
    x"2BBF15F",
    x"2BBEE63",
    x"2BBEB67",
    x"2BBE86D",
    x"2BBE573",
    x"2BBE27A",
    x"2BBDF82",
    x"2BBDC8B",
    x"2BBD994",
    x"2BBD69E",
    x"2BBD3A8",
    x"2BBD0B4",
    x"2BBCDC0",
    x"2BBCACD",
    x"2BBC7DB",
    x"2BBC4E9",
    x"2BBC1F8",
    x"2BBBF08",
    x"2BBBC19",
    x"2BBB92A",
    x"2BBB63C",
    x"2BBB34F",
    x"2BBB062",
    x"2BBAD77",
    x"2BBAA8C",
    x"2BBA7A1",
    x"2BBA4B8",
    x"2BBA1CF",
    x"2BB9EE7",
    x"2BB9C00",
    x"2BB9919",
    x"2BB9633",
    x"2BB934E",
    x"2BB9069",
    x"2BB8D86",
    x"2BB8AA3",
    x"2BB87C0",
    x"2BB84DF",
    x"2BB81FE",
    x"2BB7F1E",
    x"2BB7C3E",
    x"2BB7960",
    x"2BB7682",
    x"2BB73A4",
    x"2BB70C8",
    x"2BB6DEC",
    x"2BB6B11",
    x"2BB6837",
    x"2BB655D",
    x"2BB6284",
    x"2BB5FAC",
    x"2BB5CD4",
    x"2BB59FD",
    x"2BB5727",
    x"2BB5452",
    x"2BB517D",
    x"2BB4EA9",
    x"2BB4BD6",
    x"2BB4903",
    x"2BB4631",
    x"2BB4360",
    x"2BB408F",
    x"2BB3DC0",
    x"2BB3AF0",
    x"2BB3822",
    x"2BB3554",
    x"2BB3287",
    x"2BB2FBB",
    x"2BB2CF0",
    x"2BB2A25",
    x"2BB275A",
    x"2BB2491",
    x"2BB21C8",
    x"2BB1F00",
    x"2BB1C39",
    x"2BB1972",
    x"2BB16AC",
    x"2BB13E7",
    x"2BB1122",
    x"2BB0E5E",
    x"2BB0B9B",
    x"2BB08D8",
    x"2BB0616",
    x"2BB0355",
    x"2BB0095",
    x"2BAFDD5",
    x"2BAFB16",
    x"2BAF857",
    x"2BAF59A",
    x"2BAF2DD",
    x"2BAF020",
    x"2BAED65",
    x"2BAEAAA",
    x"2BAE7EF",
    x"2BAE536",
    x"2BAE27D",
    x"2BADFC4",
    x"2BADD0D",
    x"2BADA56",
    x"2BAD7A0",
    x"2BAD4EA",
    x"2BAD235",
    x"2BACF81",
    x"2BACCCD",
    x"2BACA1A",
    x"2BAC768",
    x"2BAC4B7",
    x"2BAC206",
    x"2BABF56",
    x"2BABCA6",
    x"2BAB9F7",
    x"2BAB749",
    x"2BAB49C",
    x"2BAB1EF",
    x"2BAAF43",
    x"2BAAC97",
    x"2BAA9EC",
    x"2BAA742",
    x"2BAA499",
    x"2BAA1F0",
    x"2BA9F48",
    x"2BA9CA0",
    x"2BA99FA",
    x"2BA9753",
    x"2BA94AE",
    x"2BA9209",
    x"2BA8F65",
    x"2BA8CC1",
    x"2BA8A1F",
    x"2BA877C",
    x"2BA84DB",
    x"2BA823A",
    x"2BA7F9A",
    x"2BA7CFA",
    x"2BA7A5B",
    x"2BA77BD",
    x"2BA751F",
    x"2BA7282",
    x"2BA6FE6",
    x"2BA6D4A",
    x"2BA6AAF",
    x"2BA6815",
    x"2BA657B",
    x"2BA62E2",
    x"2BA604A",
    x"2BA5DB2",
    x"2BA5B1B",
    x"2BA5885",
    x"2BA55EF",
    x"2BA535A",
    x"2BA50C5",
    x"2BA4E31",
    x"2BA4B9E",
    x"2BA490B",
    x"2BA467A",
    x"2BA43E8",
    x"2BA4158",
    x"2BA3EC8",
    x"2BA3C38",
    x"2BA39A9",
    x"2BA371B",
    x"2BA348E",
    x"2BA3201",
    x"2BA2F75",
    x"2BA2CE9",
    x"2BA2A5E",
    x"2BA27D4",
    x"2BA254A",
    x"2BA22C1",
    x"2BA2039",
    x"2BA1DB1",
    x"2BA1B2A",
    x"2BA18A4",
    x"2BA161E",
    x"2BA1399",
    x"2BA1114",
    x"2BA0E90",
    x"2BA0C0D",
    x"2BA098A",
    x"2BA0708",
    x"2BA0487",
    x"2BA0206",
    x"2B9FF86",
    x"2B9FD06",
    x"2B9FA87",
    x"2B9F809",
    x"2B9F58B",
    x"2B9F30E",
    x"2B9F092",
    x"2B9EE16",
    x"2B9EB9B",
    x"2B9E920",
    x"2B9E6A6",
    x"2B9E42D",
    x"2B9E1B4",
    x"2B9DF3C",
    x"2B9DCC4",
    x"2B9DA4D",
    x"2B9D7D7",
    x"2B9D561",
    x"2B9D2EC",
    x"2B9D078",
    x"2B9CE04",
    x"2B9CB91",
    x"2B9C91E",
    x"2B9C6AC",
    x"2B9C43B",
    x"2B9C1CA",
    x"2B9BF5A",
    x"2B9BCEB",
    x"2B9BA7C",
    x"2B9B80D",
    x"2B9B5A0",
    x"2B9B333",
    x"2B9B0C6",
    x"2B9AE5A",
    x"2B9ABEF",
    x"2B9A984",
    x"2B9A71A",
    x"2B9A4B1",
    x"2B9A248",
    x"2B99FE0",
    x"2B99D78",
    x"2B99B11",
    x"2B998AA",
    x"2B99644",
    x"2B993DF",
    x"2B9917B",
    x"2B98F16",
    x"2B98CB3",
    x"2B98A50",
    x"2B987EE",
    x"2B9858C",
    x"2B9832B",
    x"2B980CB",
    x"2B97E6B",
    x"2B97C0B",
    x"2B979AD",
    x"2B9774E",
    x"2B974F1",
    x"2B97294",
    x"2B97038",
    x"2B96DDC",
    x"2B96B81",
    x"2B96926",
    x"2B966CC",
    x"2B96473",
    x"2B9621A",
    x"2B95FC2",
    x"2B95D6A",
    x"2B95B13",
    x"2B958BD",
    x"2B95667",
    x"2B95411",
    x"2B951BD",
    x"2B94F68",
    x"2B94D15",
    x"2B94AC2",
    x"2B94870",
    x"2B9461E",
    x"2B943CC",
    x"2B9417C",
    x"2B93F2C",
    x"2B93CDC",
    x"2B93A8D",
    x"2B9383F",
    x"2B935F1",
    x"2B933A4",
    x"2B93157",
    x"2B92F0B",
    x"2B92CC0",
    x"2B92A75",
    x"2B9282B",
    x"2B925E1",
    x"2B92398",
    x"2B9214F",
    x"2B91F07",
    x"2B91CC0",
    x"2B91A79",
    x"2B91832",
    x"2B915ED",
    x"2B913A7",
    x"2B91163",
    x"2B90F1F",
    x"2B90CDB",
    x"2B90A98",
    x"2B90856",
    x"2B90614",
    x"2B903D3",
    x"2B90192",
    x"2B8FF52",
    x"2B8FD12",
    x"2B8FAD3",
    x"2B8F895",
    x"2B8F657",
    x"2B8F41A",
    x"2B8F1DD",
    x"2B8EFA1",
    x"2B8ED65",
    x"2B8EB2A",
    x"2B8E8F0",
    x"2B8E6B6",
    x"2B8E47C",
    x"2B8E244",
    x"2B8E00B",
    x"2B8DDD3",
    x"2B8DB9C",
    x"2B8D966",
    x"2B8D730",
    x"2B8D4FA",
    x"2B8D2C5",
    x"2B8D091",
    x"2B8CE5D",
    x"2B8CC2A",
    x"2B8C9F7",
    x"2B8C7C5",
    x"2B8C593",
    x"2B8C362",
    x"2B8C131",
    x"2B8BF01",
    x"2B8BCD2",
    x"2B8BAA3",
    x"2B8B874",
    x"2B8B647",
    x"2B8B419",
    x"2B8B1EC",
    x"2B8AFC0",
    x"2B8AD95",
    x"2B8AB69",
    x"2B8A93F",
    x"2B8A715",
    x"2B8A4EB",
    x"2B8A2C2",
    x"2B8A09A",
    x"2B89E72",
    x"2B89C4B",
    x"2B89A24",
    x"2B897FE",
    x"2B895D8",
    x"2B893B3",
    x"2B8918E",
    x"2B88F6A",
    x"2B88D46",
    x"2B88B23",
    x"2B88901",
    x"2B886DF",
    x"2B884BD",
    x"2B8829C",
    x"2B8807C",
    x"2B87E5C",
    x"2B87C3D",
    x"2B87A1E",
    x"2B87800",
    x"2B875E2",
    x"2B873C5",
    x"2B871A8",
    x"2B86F8C",
    x"2B86D70",
    x"2B86B55",
    x"2B8693B",
    x"2B86721",
    x"2B86507",
    x"2B862EE",
    x"2B860D6",
    x"2B85EBE",
    x"2B85CA6",
    x"2B85A8F",
    x"2B85879",
    x"2B85663",
    x"2B8544E",
    x"2B85239",
    x"2B85025",
    x"2B84E11",
    x"2B84BFE",
    x"2B849EB",
    x"2B847D9",
    x"2B845C7",
    x"2B843B6",
    x"2B841A5",
    x"2B83F95",
    x"2B83D85",
    x"2B83B76",
    x"2B83968",
    x"2B8375A",
    x"2B8354C",
    x"2B8333F",
    x"2B83132",
    x"2B82F26",
    x"2B82D1B",
    x"2B82B10",
    x"2B82905",
    x"2B826FB",
    x"2B824F2",
    x"2B822E9",
    x"2B820E0",
    x"2B81ED8",
    x"2B81CD1",
    x"2B81ACA",
    x"2B818C4",
    x"2B816BE",
    x"2B814B8",
    x"2B812B3",
    x"2B810AF",
    x"2B80EAB",
    x"2B80CA7",
    x"2B80AA5",
    x"2B808A2",
    x"2B806A0",
    x"2B8049F",
    x"2B8029E",
    x"2B8009E",
    x"2B7FD3C",
    x"2B7F93D",
    x"2B7F53F",
    x"2B7F142",
    x"2B7ED46",
    x"2B7E94C",
    x"2B7E552",
    x"2B7E159",
    x"2B7DD61",
    x"2B7D96A",
    x"2B7D574",
    x"2B7D180",
    x"2B7CD8C",
    x"2B7C999",
    x"2B7C5A7",
    x"2B7C1B6",
    x"2B7BDC6",
    x"2B7B9D7",
    x"2B7B5E9",
    x"2B7B1FC",
    x"2B7AE10",
    x"2B7AA25",
    x"2B7A63B",
    x"2B7A252",
    x"2B79E6A",
    x"2B79A83",
    x"2B7969D",
    x"2B792B7",
    x"2B78ED3",
    x"2B78AF0",
    x"2B7870E",
    x"2B7832C",
    x"2B77F4C",
    x"2B77B6D",
    x"2B7778E",
    x"2B773B1",
    x"2B76FD5",
    x"2B76BF9",
    x"2B7681F",
    x"2B76445",
    x"2B7606C",
    x"2B75C95",
    x"2B758BE",
    x"2B754E8",
    x"2B75114",
    x"2B74D40",
    x"2B7496D",
    x"2B7459B",
    x"2B741CA",
    x"2B73DFA",
    x"2B73A2B",
    x"2B7365D",
    x"2B73290",
    x"2B72EC4",
    x"2B72AF9",
    x"2B7272E",
    x"2B72365",
    x"2B71F9D",
    x"2B71BD5",
    x"2B7180F",
    x"2B71449",
    x"2B71085",
    x"2B70CC1",
    x"2B708FE",
    x"2B7053D",
    x"2B7017C",
    x"2B6FDBC",
    x"2B6F9FD",
    x"2B6F63F",
    x"2B6F282",
    x"2B6EEC6",
    x"2B6EB0A",
    x"2B6E750",
    x"2B6E397",
    x"2B6DFDE",
    x"2B6DC27",
    x"2B6D870",
    x"2B6D4BB",
    x"2B6D106",
    x"2B6CD52",
    x"2B6C99F",
    x"2B6C5ED",
    x"2B6C23C",
    x"2B6BE8C",
    x"2B6BADD",
    x"2B6B72F",
    x"2B6B381",
    x"2B6AFD5",
    x"2B6AC29",
    x"2B6A87F",
    x"2B6A4D5",
    x"2B6A12C",
    x"2B69D85",
    x"2B699DE",
    x"2B69638",
    x"2B69293",
    x"2B68EEE",
    x"2B68B4B",
    x"2B687A9",
    x"2B68407",
    x"2B68067",
    x"2B67CC7",
    x"2B67928",
    x"2B6758A",
    x"2B671EE",
    x"2B66E51",
    x"2B66AB6",
    x"2B6671C",
    x"2B66383",
    x"2B65FEA",
    x"2B65C53",
    x"2B658BC",
    x"2B65526",
    x"2B65192",
    x"2B64DFE",
    x"2B64A6B",
    x"2B646D8",
    x"2B64347",
    x"2B63FB7",
    x"2B63C27",
    x"2B63899",
    x"2B6350B",
    x"2B6317E",
    x"2B62DF2",
    x"2B62A67",
    x"2B626DD",
    x"2B62354",
    x"2B61FCB",
    x"2B61C44",
    x"2B618BD",
    x"2B61538",
    x"2B611B3",
    x"2B60E2F",
    x"2B60AAC",
    x"2B60729",
    x"2B603A8",
    x"2B60028",
    x"2B5FCA8",
    x"2B5F929",
    x"2B5F5AB",
    x"2B5F22E",
    x"2B5EEB2",
    x"2B5EB37",
    x"2B5E7BD",
    x"2B5E443",
    x"2B5E0CB",
    x"2B5DD53",
    x"2B5D9DC",
    x"2B5D666",
    x"2B5D2F1",
    x"2B5CF7C",
    x"2B5CC09",
    x"2B5C896",
    x"2B5C525",
    x"2B5C1B4",
    x"2B5BE44",
    x"2B5BAD5",
    x"2B5B766",
    x"2B5B3F9",
    x"2B5B08C",
    x"2B5AD21",
    x"2B5A9B6",
    x"2B5A64C",
    x"2B5A2E3",
    x"2B59F7A",
    x"2B59C13",
    x"2B598AC",
    x"2B59547",
    x"2B591E2",
    x"2B58E7E",
    x"2B58B1A",
    x"2B587B8",
    x"2B58457",
    x"2B580F6",
    x"2B57D96",
    x"2B57A37",
    x"2B576D9",
    x"2B5737C",
    x"2B5701F",
    x"2B56CC4",
    x"2B56969",
    x"2B5660F",
    x"2B562B6",
    x"2B55F5E",
    x"2B55C06",
    x"2B558B0",
    x"2B5555A",
    x"2B55205",
    x"2B54EB1",
    x"2B54B5E",
    x"2B5480B",
    x"2B544BA",
    x"2B54169",
    x"2B53E19",
    x"2B53ACA",
    x"2B5377B",
    x"2B5342E",
    x"2B530E1",
    x"2B52D96",
    x"2B52A4B",
    x"2B52700",
    x"2B523B7",
    x"2B5206F",
    x"2B51D27",
    x"2B519E0",
    x"2B5169A",
    x"2B51355",
    x"2B51010",
    x"2B50CCD",
    x"2B5098A",
    x"2B50648",
    x"2B50307",
    x"2B4FFC6",
    x"2B4FC87",
    x"2B4F948",
    x"2B4F60A",
    x"2B4F2CD",
    x"2B4EF91",
    x"2B4EC55",
    x"2B4E91B",
    x"2B4E5E1",
    x"2B4E2A8",
    x"2B4DF6F",
    x"2B4DC38",
    x"2B4D901",
    x"2B4D5CB",
    x"2B4D296",
    x"2B4CF62",
    x"2B4CC2F",
    x"2B4C8FC",
    x"2B4C5CA",
    x"2B4C299",
    x"2B4BF69",
    x"2B4BC39",
    x"2B4B90B",
    x"2B4B5DD",
    x"2B4B2B0",
    x"2B4AF84",
    x"2B4AC58",
    x"2B4A92D",
    x"2B4A603",
    x"2B4A2DA",
    x"2B49FB2",
    x"2B49C8B",
    x"2B49964",
    x"2B4963E",
    x"2B49319",
    x"2B48FF4",
    x"2B48CD1",
    x"2B489AE",
    x"2B4868C",
    x"2B4836B",
    x"2B4804A",
    x"2B47D2A",
    x"2B47A0C",
    x"2B476ED",
    x"2B473D0",
    x"2B470B4",
    x"2B46D98",
    x"2B46A7D",
    x"2B46762",
    x"2B46449",
    x"2B46130",
    x"2B45E18",
    x"2B45B01",
    x"2B457EB",
    x"2B454D5",
    x"2B451C1",
    x"2B44EAC",
    x"2B44B99",
    x"2B44887",
    x"2B44575",
    x"2B44264",
    x"2B43F54",
    x"2B43C44",
    x"2B43936",
    x"2B43628",
    x"2B4331A",
    x"2B4300E",
    x"2B42D02",
    x"2B429F8",
    x"2B426ED",
    x"2B423E4",
    x"2B420DC",
    x"2B41DD4",
    x"2B41ACD",
    x"2B417C6",
    x"2B414C1",
    x"2B411BC",
    x"2B40EB8",
    x"2B40BB5",
    x"2B408B2",
    x"2B405B0",
    x"2B402AF",
    x"2B3FFAF",
    x"2B3FCAF",
    x"2B3F9B1",
    x"2B3F6B2",
    x"2B3F3B5",
    x"2B3F0B9",
    x"2B3EDBD",
    x"2B3EAC2",
    x"2B3E7C7",
    x"2B3E4CE",
    x"2B3E1D5",
    x"2B3DEDD",
    x"2B3DBE6",
    x"2B3D8EF",
    x"2B3D5F9",
    x"2B3D304",
    x"2B3D010",
    x"2B3CD1C",
    x"2B3CA29",
    x"2B3C737",
    x"2B3C445",
    x"2B3C155",
    x"2B3BE65",
    x"2B3BB76",
    x"2B3B887",
    x"2B3B599",
    x"2B3B2AC",
    x"2B3AFC0",
    x"2B3ACD4",
    x"2B3A9EA",
    x"2B3A6FF",
    x"2B3A416",
    x"2B3A12D",
    x"2B39E45",
    x"2B39B5E",
    x"2B39878",
    x"2B39592",
    x"2B392AD",
    x"2B38FC9",
    x"2B38CE5",
    x"2B38A02",
    x"2B38720",
    x"2B3843F",
    x"2B3815E",
    x"2B37E7E",
    x"2B37B9F",
    x"2B378C0",
    x"2B375E2",
    x"2B37305",
    x"2B37029",
    x"2B36D4D",
    x"2B36A72",
    x"2B36798",
    x"2B364BE",
    x"2B361E6",
    x"2B35F0D",
    x"2B35C36",
    x"2B3595F",
    x"2B35689",
    x"2B353B4",
    x"2B350DF",
    x"2B34E0C",
    x"2B34B38",
    x"2B34866",
    x"2B34594",
    x"2B342C3",
    x"2B33FF3",
    x"2B33D23",
    x"2B33A54",
    x"2B33786",
    x"2B334B9",
    x"2B331EC",
    x"2B32F20",
    x"2B32C54",
    x"2B32989",
    x"2B326BF",
    x"2B323F6",
    x"2B3212D",
    x"2B31E65",
    x"2B31B9E",
    x"2B318D8",
    x"2B31612",
    x"2B3134D",
    x"2B31088",
    x"2B30DC4",
    x"2B30B01",
    x"2B3083F",
    x"2B3057D",
    x"2B302BC",
    x"2B2FFFC",
    x"2B2FD3C",
    x"2B2FA7D",
    x"2B2F7BF",
    x"2B2F501",
    x"2B2F244",
    x"2B2EF88",
    x"2B2ECCD",
    x"2B2EA12",
    x"2B2E758",
    x"2B2E49E",
    x"2B2E1E5",
    x"2B2DF2D",
    x"2B2DC76",
    x"2B2D9BF",
    x"2B2D709",
    x"2B2D453",
    x"2B2D19F",
    x"2B2CEEB",
    x"2B2CC37",
    x"2B2C984",
    x"2B2C6D2",
    x"2B2C421",
    x"2B2C170",
    x"2B2BEC0",
    x"2B2BC11",
    x"2B2B962",
    x"2B2B6B4",
    x"2B2B407",
    x"2B2B15A",
    x"2B2AEAE",
    x"2B2AC03",
    x"2B2A958",
    x"2B2A6AE",
    x"2B2A405",
    x"2B2A15C",
    x"2B29EB4",
    x"2B29C0D",
    x"2B29966",
    x"2B296C0",
    x"2B2941B",
    x"2B29176",
    x"2B28ED2",
    x"2B28C2F",
    x"2B2898C",
    x"2B286EA",
    x"2B28449",
    x"2B281A8",
    x"2B27F08",
    x"2B27C68",
    x"2B279C9",
    x"2B2772B",
    x"2B2748E",
    x"2B271F1",
    x"2B26F55",
    x"2B26CB9",
    x"2B26A1F",
    x"2B26784",
    x"2B264EB",
    x"2B26252",
    x"2B25FBA",
    x"2B25D22",
    x"2B25A8B",
    x"2B257F5",
    x"2B2555F",
    x"2B252CA",
    x"2B25036",
    x"2B24DA2",
    x"2B24B0F",
    x"2B2487C",
    x"2B245EB",
    x"2B24359",
    x"2B240C9",
    x"2B23E39",
    x"2B23BAA",
    x"2B2391B",
    x"2B2368D",
    x"2B23400",
    x"2B23173",
    x"2B22EE7",
    x"2B22C5C",
    x"2B229D1",
    x"2B22747",
    x"2B224BD",
    x"2B22235",
    x"2B21FAC",
    x"2B21D25",
    x"2B21A9E",
    x"2B21817",
    x"2B21592",
    x"2B2130D",
    x"2B21088",
    x"2B20E04",
    x"2B20B81",
    x"2B208FF",
    x"2B2067D",
    x"2B203FB",
    x"2B2017B",
    x"2B1FEFB",
    x"2B1FC7B",
    x"2B1F9FC",
    x"2B1F77E",
    x"2B1F501",
    x"2B1F284",
    x"2B1F007",
    x"2B1ED8C",
    x"2B1EB11",
    x"2B1E896",
    x"2B1E61C",
    x"2B1E3A3",
    x"2B1E12A",
    x"2B1DEB2",
    x"2B1DC3B",
    x"2B1D9C4",
    x"2B1D74E",
    x"2B1D4D9",
    x"2B1D264",
    x"2B1CFF0",
    x"2B1CD7C",
    x"2B1CB09",
    x"2B1C896",
    x"2B1C624",
    x"2B1C3B3",
    x"2B1C143",
    x"2B1BED3",
    x"2B1BC63",
    x"2B1B9F4",
    x"2B1B786",
    x"2B1B519",
    x"2B1B2AC",
    x"2B1B03F",
    x"2B1ADD4",
    x"2B1AB68",
    x"2B1A8FE",
    x"2B1A694",
    x"2B1A42B",
    x"2B1A1C2",
    x"2B19F5A",
    x"2B19CF2",
    x"2B19A8B",
    x"2B19825",
    x"2B195BF",
    x"2B1935A",
    x"2B190F5",
    x"2B18E92",
    x"2B18C2E",
    x"2B189CB",
    x"2B18769",
    x"2B18508",
    x"2B182A7",
    x"2B18046",
    x"2B17DE7",
    x"2B17B87",
    x"2B17929",
    x"2B176CB",
    x"2B1746D",
    x"2B17211",
    x"2B16FB4",
    x"2B16D59",
    x"2B16AFE",
    x"2B168A3",
    x"2B16649",
    x"2B163F0",
    x"2B16197",
    x"2B15F3F",
    x"2B15CE8",
    x"2B15A91",
    x"2B1583B",
    x"2B155E5",
    x"2B15390",
    x"2B1513B",
    x"2B14EE7",
    x"2B14C94",
    x"2B14A41",
    x"2B147EE",
    x"2B1459D",
    x"2B1434C",
    x"2B140FB",
    x"2B13EAB",
    x"2B13C5C",
    x"2B13A0D",
    x"2B137BF",
    x"2B13571",
    x"2B13324",
    x"2B130D8",
    x"2B12E8C",
    x"2B12C40",
    x"2B129F5",
    x"2B127AB",
    x"2B12562",
    x"2B12319",
    x"2B120D0",
    x"2B11E88",
    x"2B11C41",
    x"2B119FA",
    x"2B117B4",
    x"2B1156E",
    x"2B11329",
    x"2B110E5",
    x"2B10EA1",
    x"2B10C5D",
    x"2B10A1A",
    x"2B107D8",
    x"2B10597",
    x"2B10355",
    x"2B10115",
    x"2B0FED5",
    x"2B0FC95",
    x"2B0FA57",
    x"2B0F818",
    x"2B0F5DB",
    x"2B0F39D",
    x"2B0F161",
    x"2B0EF25",
    x"2B0ECE9",
    x"2B0EAAE",
    x"2B0E874",
    x"2B0E63A",
    x"2B0E401",
    x"2B0E1C8",
    x"2B0DF90",
    x"2B0DD58",
    x"2B0DB21",
    x"2B0D8EB",
    x"2B0D6B5",
    x"2B0D47F",
    x"2B0D24A",
    x"2B0D016",
    x"2B0CDE2",
    x"2B0CBAF",
    x"2B0C97D",
    x"2B0C74A",
    x"2B0C519",
    x"2B0C2E8",
    x"2B0C0B7",
    x"2B0BE88",
    x"2B0BC58",
    x"2B0BA29",
    x"2B0B7FB",
    x"2B0B5CD",
    x"2B0B3A0",
    x"2B0B174",
    x"2B0AF47",
    x"2B0AD1C",
    x"2B0AAF1",
    x"2B0A8C6",
    x"2B0A69D",
    x"2B0A473",
    x"2B0A24A",
    x"2B0A022",
    x"2B09DFA",
    x"2B09BD3",
    x"2B099AC",
    x"2B09786",
    x"2B09561",
    x"2B0933B",
    x"2B09117",
    x"2B08EF3",
    x"2B08CCF",
    x"2B08AAD",
    x"2B0888A",
    x"2B08668",
    x"2B08447",
    x"2B08226",
    x"2B08006",
    x"2B07DE6",
    x"2B07BC7",
    x"2B079A8",
    x"2B0778A",
    x"2B0756C",
    x"2B0734F",
    x"2B07133",
    x"2B06F17",
    x"2B06CFB",
    x"2B06AE0",
    x"2B068C6",
    x"2B066AC",
    x"2B06492",
    x"2B0627A",
    x"2B06061",
    x"2B05E49",
    x"2B05C32",
    x"2B05A1B",
    x"2B05805",
    x"2B055EF",
    x"2B053DA",
    x"2B051C5",
    x"2B04FB1",
    x"2B04D9E",
    x"2B04B8A",
    x"2B04978",
    x"2B04766",
    x"2B04554",
    x"2B04343",
    x"2B04132",
    x"2B03F22",
    x"2B03D13",
    x"2B03B04",
    x"2B038F5",
    x"2B036E7",
    x"2B034DA",
    x"2B032CD",
    x"2B030C0",
    x"2B02EB5",
    x"2B02CA9",
    x"2B02A9E",
    x"2B02894",
    x"2B0268A",
    x"2B02481",
    x"2B02278",
    x"2B0206F",
    x"2B01E67",
    x"2B01C60",
    x"2B01A59",
    x"2B01853",
    x"2B0164D",
    x"2B01448",
    x"2B01243",
    x"2B0103F",
    x"2B00E3B",
    x"2B00C38",
    x"2B00A35",
    x"2B00832",
    x"2B00631",
    x"2B0042F",
    x"2B0022F",
    x"2B0002E",
    x"2AFFC5D",
    x"2AFF85F",
    x"2AFF461",
    x"2AFF065",
    x"2AFEC69",
    x"2AFE86E",
    x"2AFE475",
    x"2AFE07C",
    x"2AFDC85",
    x"2AFD88E",
    x"2AFD498",
    x"2AFD0A4",
    x"2AFCCB0",
    x"2AFC8BD",
    x"2AFC4CC",
    x"2AFC0DB",
    x"2AFBCEB",
    x"2AFB8FC",
    x"2AFB50F",
    x"2AFB122",
    x"2AFAD36",
    x"2AFA94B",
    x"2AFA561",
    x"2AFA179",
    x"2AF9D91",
    x"2AF99AA",
    x"2AF95C4",
    x"2AF91DF",
    x"2AF8DFB",
    x"2AF8A18",
    x"2AF8636",
    x"2AF8255",
    x"2AF7E75",
    x"2AF7A96",
    x"2AF76B7",
    x"2AF72DA",
    x"2AF6EFE",
    x"2AF6B23",
    x"2AF6748",
    x"2AF636F",
    x"2AF5F97",
    x"2AF5BBF",
    x"2AF57E9",
    x"2AF5413",
    x"2AF503F",
    x"2AF4C6B",
    x"2AF4899",
    x"2AF44C7",
    x"2AF40F6",
    x"2AF3D26",
    x"2AF3958",
    x"2AF358A",
    x"2AF31BD",
    x"2AF2DF1",
    x"2AF2A26",
    x"2AF265C",
    x"2AF2293",
    x"2AF1ECA",
    x"2AF1B03",
    x"2AF173D",
    x"2AF1378",
    x"2AF0FB3",
    x"2AF0BF0",
    x"2AF082D",
    x"2AF046C",
    x"2AF00AB",
    x"2AEFCEB",
    x"2AEF92D",
    x"2AEF56F",
    x"2AEF1B2",
    x"2AEEDF6",
    x"2AEEA3B",
    x"2AEE681",
    x"2AEE2C8",
    x"2AEDF0F",
    x"2AEDB58",
    x"2AED7A2",
    x"2AED3EC",
    x"2AED038",
    x"2AECC84",
    x"2AEC8D2",
    x"2AEC520",
    x"2AEC16F",
    x"2AEBDBF",
    x"2AEBA10",
    x"2AEB662",
    x"2AEB2B5",
    x"2AEAF09",
    x"2AEAB5D",
    x"2AEA7B3",
    x"2AEA40A",
    x"2AEA061",
    x"2AE9CB9",
    x"2AE9913",
    x"2AE956D",
    x"2AE91C8",
    x"2AE8E24",
    x"2AE8A81",
    x"2AE86DF",
    x"2AE833D",
    x"2AE7F9D",
    x"2AE7BFE",
    x"2AE785F",
    x"2AE74C1",
    x"2AE7125",
    x"2AE6D89",
    x"2AE69EE",
    x"2AE6654",
    x"2AE62BB",
    x"2AE5F22",
    x"2AE5B8B",
    x"2AE57F5",
    x"2AE545F",
    x"2AE50CB",
    x"2AE4D37",
    x"2AE49A4",
    x"2AE4612",
    x"2AE4281",
    x"2AE3EF1",
    x"2AE3B61",
    x"2AE37D3",
    x"2AE3446",
    x"2AE30B9",
    x"2AE2D2D",
    x"2AE29A2",
    x"2AE2618",
    x"2AE228F",
    x"2AE1F07",
    x"2AE1B80",
    x"2AE17F9",
    x"2AE1474",
    x"2AE10EF",
    x"2AE0D6B",
    x"2AE09E8",
    x"2AE0666",
    x"2AE02E5",
    x"2ADFF65",
    x"2ADFBE5",
    x"2ADF867",
    x"2ADF4E9",
    x"2ADF16C",
    x"2ADEDF1",
    x"2ADEA75",
    x"2ADE6FB",
    x"2ADE382",
    x"2ADE00A",
    x"2ADDC92",
    x"2ADD91B",
    x"2ADD5A5",
    x"2ADD230",
    x"2ADCEBC",
    x"2ADCB49",
    x"2ADC7D7",
    x"2ADC465",
    x"2ADC0F4",
    x"2ADBD85",
    x"2ADBA16",
    x"2ADB6A8",
    x"2ADB33A",
    x"2ADAFCE",
    x"2ADAC62",
    x"2ADA8F8",
    x"2ADA58E",
    x"2ADA225",
    x"2AD9EBD",
    x"2AD9B56",
    x"2AD97EF",
    x"2AD948A",
    x"2AD9125",
    x"2AD8DC1",
    x"2AD8A5E",
    x"2AD86FC",
    x"2AD839B",
    x"2AD803A",
    x"2AD7CDB",
    x"2AD797C",
    x"2AD761E",
    x"2AD72C1",
    x"2AD6F64",
    x"2AD6C09",
    x"2AD68AE",
    x"2AD6555",
    x"2AD61FC",
    x"2AD5EA4",
    x"2AD5B4C",
    x"2AD57F6",
    x"2AD54A0",
    x"2AD514C",
    x"2AD4DF8",
    x"2AD4AA5",
    x"2AD4752",
    x"2AD4401",
    x"2AD40B0",
    x"2AD3D61",
    x"2AD3A12",
    x"2AD36C4",
    x"2AD3376",
    x"2AD302A",
    x"2AD2CDE",
    x"2AD2993",
    x"2AD2649",
    x"2AD2300",
    x"2AD1FB8",
    x"2AD1C70",
    x"2AD192A",
    x"2AD15E4",
    x"2AD129F",
    x"2AD0F5B",
    x"2AD0C17",
    x"2AD08D5",
    x"2AD0593",
    x"2AD0252",
    x"2ACFF12",
    x"2ACFBD2",
    x"2ACF894",
    x"2ACF556",
    x"2ACF219",
    x"2ACEEDD",
    x"2ACEBA2",
    x"2ACE867",
    x"2ACE52D",
    x"2ACE1F4",
    x"2ACDEBC",
    x"2ACDB85",
    x"2ACD84F",
    x"2ACD519",
    x"2ACD1E4",
    x"2ACCEB0",
    x"2ACCB7D",
    x"2ACC84A",
    x"2ACC519",
    x"2ACC1E8",
    x"2ACBEB8",
    x"2ACBB88",
    x"2ACB85A",
    x"2ACB52C",
    x"2ACB1FF",
    x"2ACAED3",
    x"2ACABA8",
    x"2ACA87D",
    x"2ACA554",
    x"2ACA22B",
    x"2AC9F03",
    x"2AC9BDB",
    x"2AC98B5",
    x"2AC958F",
    x"2AC926A",
    x"2AC8F46",
    x"2AC8C22",
    x"2AC8900",
    x"2AC85DE",
    x"2AC82BD",
    x"2AC7F9C",
    x"2AC7C7D",
    x"2AC795E",
    x"2AC7640",
    x"2AC7323",
    x"2AC7007",
    x"2AC6CEB",
    x"2AC69D0",
    x"2AC66B6",
    x"2AC639D",
    x"2AC6084",
    x"2AC5D6C",
    x"2AC5A55",
    x"2AC573F",
    x"2AC542A",
    x"2AC5115",
    x"2AC4E01",
    x"2AC4AEE",
    x"2AC47DC",
    x"2AC44CA",
    x"2AC41B9",
    x"2AC3EA9",
    x"2AC3B9A",
    x"2AC388C",
    x"2AC357E",
    x"2AC3271",
    x"2AC2F65",
    x"2AC2C59",
    x"2AC294E",
    x"2AC2645",
    x"2AC233B",
    x"2AC2033",
    x"2AC1D2B",
    x"2AC1A24",
    x"2AC171E",
    x"2AC1419",
    x"2AC1114",
    x"2AC0E10",
    x"2AC0B0D",
    x"2AC080B",
    x"2AC0509",
    x"2AC0208",
    x"2ABFF08",
    x"2ABFC09",
    x"2ABF90A",
    x"2ABF60C",
    x"2ABF30F",
    x"2ABF013",
    x"2ABED17",
    x"2ABEA1C",
    x"2ABE722",
    x"2ABE428",
    x"2ABE130",
    x"2ABDE38",
    x"2ABDB41",
    x"2ABD84A",
    x"2ABD555",
    x"2ABD260",
    x"2ABCF6B",
    x"2ABCC78",
    x"2ABC985",
    x"2ABC693",
    x"2ABC3A2",
    x"2ABC0B1",
    x"2ABBDC1",
    x"2ABBAD2",
    x"2ABB7E4",
    x"2ABB4F6",
    x"2ABB20A",
    x"2ABAF1D",
    x"2ABAC32",
    x"2ABA947",
    x"2ABA65D",
    x"2ABA374",
    x"2ABA08C",
    x"2AB9DA4",
    x"2AB9ABD",
    x"2AB97D7",
    x"2AB94F1",
    x"2AB920C",
    x"2AB8F28",
    x"2AB8C44",
    x"2AB8962",
    x"2AB8680",
    x"2AB839F",
    x"2AB80BE",
    x"2AB7DDE",
    x"2AB7AFF",
    x"2AB7821",
    x"2AB7543",
    x"2AB7266",
    x"2AB6F8A",
    x"2AB6CAE",
    x"2AB69D3",
    x"2AB66F9",
    x"2AB6420",
    x"2AB6147",
    x"2AB5E6F",
    x"2AB5B98",
    x"2AB58C2",
    x"2AB55EC",
    x"2AB5317",
    x"2AB5042",
    x"2AB4D6E",
    x"2AB4A9B",
    x"2AB47C9",
    x"2AB44F8",
    x"2AB4227",
    x"2AB3F56",
    x"2AB3C87",
    x"2AB39B8",
    x"2AB36EA",
    x"2AB341D",
    x"2AB3150",
    x"2AB2E84",
    x"2AB2BB9",
    x"2AB28EE",
    x"2AB2624",
    x"2AB235B",
    x"2AB2093",
    x"2AB1DCB",
    x"2AB1B04",
    x"2AB183D",
    x"2AB1578",
    x"2AB12B3",
    x"2AB0FEE",
    x"2AB0D2B",
    x"2AB0A68",
    x"2AB07A5",
    x"2AB04E4",
    x"2AB0223",
    x"2AAFF63",
    x"2AAFCA3",
    x"2AAF9E4",
    x"2AAF726",
    x"2AAF469",
    x"2AAF1AC",
    x"2AAEEF0",
    x"2AAEC35",
    x"2AAE97A",
    x"2AAE6C0",
    x"2AAE407",
    x"2AAE14E",
    x"2AADE96",
    x"2AADBDF",
    x"2AAD928",
    x"2AAD672",
    x"2AAD3BD",
    x"2AAD108",
    x"2AACE54",
    x"2AACBA1",
    x"2AAC8EE",
    x"2AAC63D",
    x"2AAC38B",
    x"2AAC0DB",
    x"2AABE2B",
    x"2AABB7C",
    x"2AAB8CD",
    x"2AAB61F",
    x"2AAB372",
    x"2AAB0C6",
    x"2AAAE1A",
    x"2AAAB6E",
    x"2AAA8C4",
    x"2AAA61A",
    x"2AAA371",
    x"2AAA0C8",
    x"2AA9E21",
    x"2AA9B79",
    x"2AA98D3",
    x"2AA962D",
    x"2AA9388",
    x"2AA90E3",
    x"2AA8E3F",
    x"2AA8B9C",
    x"2AA88F9",
    x"2AA8658",
    x"2AA83B6",
    x"2AA8116",
    x"2AA7E76",
    x"2AA7BD6",
    x"2AA7938",
    x"2AA769A",
    x"2AA73FD",
    x"2AA7160",
    x"2AA6EC4",
    x"2AA6C28",
    x"2AA698E",
    x"2AA66F4",
    x"2AA645A",
    x"2AA61C1",
    x"2AA5F29",
    x"2AA5C92",
    x"2AA59FB",
    x"2AA5765",
    x"2AA54CF",
    x"2AA523B",
    x"2AA4FA6",
    x"2AA4D13",
    x"2AA4A80",
    x"2AA47ED",
    x"2AA455C",
    x"2AA42CB",
    x"2AA403A",
    x"2AA3DAB",
    x"2AA3B1C",
    x"2AA388D",
    x"2AA35FF",
    x"2AA3372",
    x"2AA30E6",
    x"2AA2E5A",
    x"2AA2BCE",
    x"2AA2944",
    x"2AA26BA",
    x"2AA2430",
    x"2AA21A8",
    x"2AA1F20",
    x"2AA1C98",
    x"2AA1A11",
    x"2AA178B",
    x"2AA1505",
    x"2AA1281",
    x"2AA0FFC",
    x"2AA0D79",
    x"2AA0AF5",
    x"2AA0873",
    x"2AA05F1",
    x"2AA0370",
    x"2AA00F0",
    x"2A9FE70",
    x"2A9FBF0",
    x"2A9F972",
    x"2A9F6F4",
    x"2A9F476",
    x"2A9F1F9",
    x"2A9EF7D",
    x"2A9ED02",
    x"2A9EA87",
    x"2A9E80C",
    x"2A9E593",
    x"2A9E31A",
    x"2A9E0A1",
    x"2A9DE29",
    x"2A9DBB2",
    x"2A9D93B",
    x"2A9D6C5",
    x"2A9D450",
    x"2A9D1DB",
    x"2A9CF67",
    x"2A9CCF4",
    x"2A9CA81",
    x"2A9C80E",
    x"2A9C59D",
    x"2A9C32B",
    x"2A9C0BB",
    x"2A9BE4B",
    x"2A9BBDC",
    x"2A9B96D",
    x"2A9B6FF",
    x"2A9B492",
    x"2A9B225",
    x"2A9AFB9",
    x"2A9AD4D",
    x"2A9AAE2",
    x"2A9A878",
    x"2A9A60E",
    x"2A9A3A5",
    x"2A9A13C",
    x"2A99ED4",
    x"2A99C6C",
    x"2A99A06",
    x"2A9979F",
    x"2A9953A",
    x"2A992D5",
    x"2A99070",
    x"2A98E0D",
    x"2A98BA9",
    x"2A98947",
    x"2A986E5",
    x"2A98483",
    x"2A98223",
    x"2A97FC2",
    x"2A97D63",
    x"2A97B04",
    x"2A978A5",
    x"2A97647",
    x"2A973EA",
    x"2A9718D",
    x"2A96F31",
    x"2A96CD6",
    x"2A96A7B",
    x"2A96820",
    x"2A965C7",
    x"2A9636E",
    x"2A96115",
    x"2A95EBD",
    x"2A95C66",
    x"2A95A0F",
    x"2A957B9",
    x"2A95563",
    x"2A9530E",
    x"2A950B9",
    x"2A94E66",
    x"2A94C12",
    x"2A949C0",
    x"2A9476D",
    x"2A9451C",
    x"2A942CB",
    x"2A9407A",
    x"2A93E2B",
    x"2A93BDB",
    x"2A9398D",
    x"2A9373F",
    x"2A934F1",
    x"2A932A4",
    x"2A93058",
    x"2A92E0C",
    x"2A92BC1",
    x"2A92976",
    x"2A9272C",
    x"2A924E2",
    x"2A9229A",
    x"2A92051",
    x"2A91E09",
    x"2A91BC2",
    x"2A9197B",
    x"2A91735",
    x"2A914F0",
    x"2A912AB",
    x"2A91067",
    x"2A90E23",
    x"2A90BDF",
    x"2A9099D",
    x"2A9075B",
    x"2A90519",
    x"2A902D8",
    x"2A90098",
    x"2A8FE58",
    x"2A8FC19",
    x"2A8F9DA",
    x"2A8F79C",
    x"2A8F55E",
    x"2A8F321",
    x"2A8F0E4",
    x"2A8EEA8",
    x"2A8EC6D",
    x"2A8EA32",
    x"2A8E7F8",
    x"2A8E5BE",
    x"2A8E385",
    x"2A8E14C",
    x"2A8DF14",
    x"2A8DCDD",
    x"2A8DAA6",
    x"2A8D870",
    x"2A8D63A",
    x"2A8D405",
    x"2A8D1D0",
    x"2A8CF9C",
    x"2A8CD68",
    x"2A8CB35",
    x"2A8C902",
    x"2A8C6D0",
    x"2A8C49F",
    x"2A8C26E",
    x"2A8C03E",
    x"2A8BE0E",
    x"2A8BBDF",
    x"2A8B9B0",
    x"2A8B782",
    x"2A8B554",
    x"2A8B327",
    x"2A8B0FB",
    x"2A8AECF",
    x"2A8ACA3",
    x"2A8AA78",
    x"2A8A84E",
    x"2A8A624",
    x"2A8A3FB",
    x"2A8A1D2",
    x"2A89FAA",
    x"2A89D82",
    x"2A89B5B",
    x"2A89935",
    x"2A8970F",
    x"2A894E9",
    x"2A892C4",
    x"2A890A0",
    x"2A88E7C",
    x"2A88C59",
    x"2A88A36",
    x"2A88813",
    x"2A885F2",
    x"2A883D1",
    x"2A881B0",
    x"2A87F90",
    x"2A87D70",
    x"2A87B51",
    x"2A87932",
    x"2A87714",
    x"2A874F7",
    x"2A872DA",
    x"2A870BD",
    x"2A86EA1",
    x"2A86C86",
    x"2A86A6B",
    x"2A86851",
    x"2A86637",
    x"2A8641E",
    x"2A86205",
    x"2A85FED",
    x"2A85DD5",
    x"2A85BBE",
    x"2A859A7",
    x"2A85791",
    x"2A8557B",
    x"2A85366",
    x"2A85152",
    x"2A84F3E",
    x"2A84D2A",
    x"2A84B17",
    x"2A84905",
    x"2A846F3",
    x"2A844E1",
    x"2A842D0",
    x"2A840C0",
    x"2A83EB0",
    x"2A83CA0",
    x"2A83A91",
    x"2A83883",
    x"2A83675",
    x"2A83468",
    x"2A8325B",
    x"2A8304F",
    x"2A82E43",
    x"2A82C37",
    x"2A82A2D",
    x"2A82822",
    x"2A82619",
    x"2A8240F",
    x"2A82207",
    x"2A81FFE",
    x"2A81DF7",
    x"2A81BEF",
    x"2A819E9",
    x"2A817E2",
    x"2A815DD",
    x"2A813D7",
    x"2A811D3",
    x"2A80FCF",
    x"2A80DCB",
    x"2A80BC8",
    x"2A809C5",
    x"2A807C3",
    x"2A805C1",
    x"2A803C0",
    x"2A801BF",
    x"2A7FF7E",
    x"2A7FB7F",
    x"2A7F781",
    x"2A7F383",
    x"2A7EF87",
    x"2A7EB8C",
    x"2A7E791",
    x"2A7E398",
    x"2A7DF9F",
    x"2A7DBA8",
    x"2A7D7B2",
    x"2A7D3BC",
    x"2A7CFC8",
    x"2A7CBD4",
    x"2A7C7E2",
    x"2A7C3F0",
    x"2A7C000",
    x"2A7BC10",
    x"2A7B822",
    x"2A7B434",
    x"2A7B048",
    x"2A7AC5C",
    x"2A7A871",
    x"2A7A488",
    x"2A7A09F",
    x"2A79CB8",
    x"2A798D1",
    x"2A794EB",
    x"2A79106",
    x"2A78D23",
    x"2A78940",
    x"2A7855E",
    x"2A7817D",
    x"2A77D9D",
    x"2A779BE",
    x"2A775E0",
    x"2A77203",
    x"2A76E27",
    x"2A76A4C",
    x"2A76672",
    x"2A76299",
    x"2A75EC1",
    x"2A75AEA",
    x"2A75713",
    x"2A7533E",
    x"2A74F6A",
    x"2A74B96",
    x"2A747C4",
    x"2A743F3",
    x"2A74022",
    x"2A73C53",
    x"2A73884",
    x"2A734B6",
    x"2A730EA",
    x"2A72D1E",
    x"2A72953",
    x"2A72589",
    x"2A721C0",
    x"2A71DF8",
    x"2A71A31",
    x"2A7166B",
    x"2A712A6",
    x"2A70EE2",
    x"2A70B1F",
    x"2A7075C",
    x"2A7039B",
    x"2A6FFDA",
    x"2A6FC1B",
    x"2A6F85C",
    x"2A6F49F",
    x"2A6F0E2",
    x"2A6ED26",
    x"2A6E96C",
    x"2A6E5B2",
    x"2A6E1F9",
    x"2A6DE41",
    x"2A6DA8A",
    x"2A6D6D3",
    x"2A6D31E",
    x"2A6CF6A",
    x"2A6CBB6",
    x"2A6C804",
    x"2A6C452",
    x"2A6C0A2",
    x"2A6BCF2",
    x"2A6B943",
    x"2A6B595",
    x"2A6B1E9",
    x"2A6AE3D",
    x"2A6AA91",
    x"2A6A6E7",
    x"2A6A33E",
    x"2A69F96",
    x"2A69BEE",
    x"2A69848",
    x"2A694A2",
    x"2A690FD",
    x"2A68D5A",
    x"2A689B7",
    x"2A68615",
    x"2A68274",
    x"2A67ED3",
    x"2A67B34",
    x"2A67796",
    x"2A673F8",
    x"2A6705C",
    x"2A66CC0",
    x"2A66925",
    x"2A6658C",
    x"2A661F3",
    x"2A65E5B",
    x"2A65AC4",
    x"2A6572D",
    x"2A65398",
    x"2A65003",
    x"2A64C70",
    x"2A648DD",
    x"2A6454B",
    x"2A641BB",
    x"2A63E2B",
    x"2A63A9C",
    x"2A6370D",
    x"2A63380",
    x"2A62FF4",
    x"2A62C68",
    x"2A628DD",
    x"2A62554",
    x"2A621CB",
    x"2A61E43",
    x"2A61ABC",
    x"2A61735",
    x"2A613B0",
    x"2A6102B",
    x"2A60CA8",
    x"2A60925",
    x"2A605A3",
    x"2A60222",
    x"2A5FEA2",
    x"2A5FB23",
    x"2A5F7A5",
    x"2A5F427",
    x"2A5F0AB",
    x"2A5ED2F",
    x"2A5E9B4",
    x"2A5E63A",
    x"2A5E2C1",
    x"2A5DF49",
    x"2A5DBD1",
    x"2A5D85B",
    x"2A5D4E5",
    x"2A5D170",
    x"2A5CDFC",
    x"2A5CA89",
    x"2A5C717",
    x"2A5C3A6",
    x"2A5C035",
    x"2A5BCC6",
    x"2A5B957",
    x"2A5B5E9",
    x"2A5B27C",
    x"2A5AF10",
    x"2A5ABA4",
    x"2A5A83A",
    x"2A5A4D0",
    x"2A5A167",
    x"2A59E00",
    x"2A59A98",
    x"2A59732",
    x"2A593CD",
    x"2A59068",
    x"2A58D05",
    x"2A589A2",
    x"2A58640",
    x"2A582DF",
    x"2A57F7E",
    x"2A57C1F",
    x"2A578C0",
    x"2A57563",
    x"2A57206",
    x"2A56EAA",
    x"2A56B4E",
    x"2A567F4",
    x"2A5649A",
    x"2A56142",
    x"2A55DEA",
    x"2A55A93",
    x"2A5573C",
    x"2A553E7",
    x"2A55092",
    x"2A54D3F",
    x"2A549EC",
    x"2A5469A",
    x"2A54349",
    x"2A53FF8",
    x"2A53CA9",
    x"2A5395A",
    x"2A5360C",
    x"2A532BF",
    x"2A52F73",
    x"2A52C27",
    x"2A528DC",
    x"2A52593",
    x"2A5224A",
    x"2A51F01",
    x"2A51BBA",
    x"2A51874",
    x"2A5152E",
    x"2A511E9",
    x"2A50EA5",
    x"2A50B62",
    x"2A5081F",
    x"2A504DE",
    x"2A5019D",
    x"2A4FE5D",
    x"2A4FB1E",
    x"2A4F7DF",
    x"2A4F4A2",
    x"2A4F165",
    x"2A4EE29",
    x"2A4EAEE",
    x"2A4E7B4",
    x"2A4E47A",
    x"2A4E141",
    x"2A4DE09",
    x"2A4DAD2",
    x"2A4D79C",
    x"2A4D466",
    x"2A4D132",
    x"2A4CDFE",
    x"2A4CACB",
    x"2A4C799",
    x"2A4C467",
    x"2A4C136",
    x"2A4BE06",
    x"2A4BAD7",
    x"2A4B7A9",
    x"2A4B47B",
    x"2A4B14F",
    x"2A4AE23",
    x"2A4AAF8",
    x"2A4A7CD",
    x"2A4A4A4",
    x"2A4A17B",
    x"2A49E53",
    x"2A49B2C",
    x"2A49805",
    x"2A494E0",
    x"2A491BB",
    x"2A48E97",
    x"2A48B74",
    x"2A48851",
    x"2A48530",
    x"2A4820F",
    x"2A47EEF",
    x"2A47BCF",
    x"2A478B1",
    x"2A47593",
    x"2A47276",
    x"2A46F5A",
    x"2A46C3E",
    x"2A46923",
    x"2A4660A",
    x"2A462F0",
    x"2A45FD8",
    x"2A45CC1",
    x"2A459AA",
    x"2A45694",
    x"2A4537E",
    x"2A4506A",
    x"2A44D56",
    x"2A44A43",
    x"2A44731",
    x"2A44420",
    x"2A4410F",
    x"2A43DFF",
    x"2A43AF0",
    x"2A437E2",
    x"2A434D4",
    x"2A431C7",
    x"2A42EBB",
    x"2A42BB0",
    x"2A428A5",
    x"2A4259C",
    x"2A42293",
    x"2A41F8A",
    x"2A41C83",
    x"2A4197C",
    x"2A41676",
    x"2A41371",
    x"2A4106C",
    x"2A40D69",
    x"2A40A66",
    x"2A40763",
    x"2A40462",
    x"2A40161",
    x"2A3FE61",
    x"2A3FB62",
    x"2A3F864",
    x"2A3F566",
    x"2A3F269",
    x"2A3EF6D",
    x"2A3EC71",
    x"2A3E976",
    x"2A3E67C",
    x"2A3E383",
    x"2A3E08B",
    x"2A3DD93",
    x"2A3DA9C",
    x"2A3D7A6",
    x"2A3D4B0",
    x"2A3D1BB",
    x"2A3CEC7",
    x"2A3CBD4",
    x"2A3C8E1",
    x"2A3C5EF",
    x"2A3C2FE",
    x"2A3C00E",
    x"2A3BD1E",
    x"2A3BA2F",
    x"2A3B741",
    x"2A3B454",
    x"2A3B167",
    x"2A3AE7B",
    x"2A3AB90",
    x"2A3A8A5",
    x"2A3A5BB",
    x"2A3A2D2",
    x"2A39FEA",
    x"2A39D02",
    x"2A39A1B",
    x"2A39735",
    x"2A39450",
    x"2A3916B",
    x"2A38E87",
    x"2A38BA4",
    x"2A388C1",
    x"2A385E0",
    x"2A382FE",
    x"2A3801E",
    x"2A37D3E",
    x"2A37A5F",
    x"2A37781",
    x"2A374A4",
    x"2A371C7",
    x"2A36EEB",
    x"2A36C0F",
    x"2A36935",
    x"2A3665B",
    x"2A36382",
    x"2A360A9",
    x"2A35DD1",
    x"2A35AFA",
    x"2A35824",
    x"2A3554E",
    x"2A35279",
    x"2A34FA5",
    x"2A34CD1",
    x"2A349FE",
    x"2A3472C",
    x"2A3445B",
    x"2A3418A",
    x"2A33EBA",
    x"2A33BEB",
    x"2A3391C",
    x"2A3364E",
    x"2A33381",
    x"2A330B4",
    x"2A32DE9",
    x"2A32B1D",
    x"2A32853",
    x"2A32589",
    x"2A322C0",
    x"2A31FF8",
    x"2A31D30",
    x"2A31A69",
    x"2A317A3",
    x"2A314DD",
    x"2A31219",
    x"2A30F54",
    x"2A30C91",
    x"2A309CE",
    x"2A3070C",
    x"2A3044B",
    x"2A3018A",
    x"2A2FECA",
    x"2A2FC0B",
    x"2A2F94C",
    x"2A2F68E",
    x"2A2F3D1",
    x"2A2F114",
    x"2A2EE58",
    x"2A2EB9D",
    x"2A2E8E2",
    x"2A2E628",
    x"2A2E36F",
    x"2A2E0B7",
    x"2A2DDFF",
    x"2A2DB48",
    x"2A2D891",
    x"2A2D5DB",
    x"2A2D326",
    x"2A2D072",
    x"2A2CDBE",
    x"2A2CB0B",
    x"2A2C858",
    x"2A2C5A7",
    x"2A2C2F6",
    x"2A2C045",
    x"2A2BD95",
    x"2A2BAE6",
    x"2A2B838",
    x"2A2B58A",
    x"2A2B2DD",
    x"2A2B031",
    x"2A2AD85",
    x"2A2AADA",
    x"2A2A830",
    x"2A2A586",
    x"2A2A2DD",
    x"2A2A035",
    x"2A29D8D",
    x"2A29AE6",
    x"2A2983F",
    x"2A2959A",
    x"2A292F5",
    x"2A29050",
    x"2A28DAC",
    x"2A28B09",
    x"2A28867",
    x"2A285C5",
    x"2A28324",
    x"2A28084",
    x"2A27DE4",
    x"2A27B45",
    x"2A278A6",
    x"2A27608",
    x"2A2736B",
    x"2A270CF",
    x"2A26E33",
    x"2A26B98",
    x"2A268FD",
    x"2A26663",
    x"2A263CA",
    x"2A26131",
    x"2A25E99",
    x"2A25C02",
    x"2A2596B",
    x"2A256D5",
    x"2A25440",
    x"2A251AB",
    x"2A24F17",
    x"2A24C83",
    x"2A249F1",
    x"2A2475E",
    x"2A244CD",
    x"2A2423C",
    x"2A23FAC",
    x"2A23D1C",
    x"2A23A8D",
    x"2A237FF",
    x"2A23571",
    x"2A232E4",
    x"2A23058",
    x"2A22DCC",
    x"2A22B41",
    x"2A228B6",
    x"2A2262D",
    x"2A223A3",
    x"2A2211B",
    x"2A21E93",
    x"2A21C0B",
    x"2A21985",
    x"2A216FF",
    x"2A21479",
    x"2A211F4",
    x"2A20F70",
    x"2A20CED",
    x"2A20A6A",
    x"2A207E8",
    x"2A20566",
    x"2A202E5",
    x"2A20064",
    x"2A1FDE5",
    x"2A1FB65",
    x"2A1F8E7",
    x"2A1F669",
    x"2A1F3EC",
    x"2A1F16F",
    x"2A1EEF3",
    x"2A1EC78",
    x"2A1E9FD",
    x"2A1E783",
    x"2A1E509",
    x"2A1E290",
    x"2A1E018",
    x"2A1DDA0",
    x"2A1DB29",
    x"2A1D8B2",
    x"2A1D63D",
    x"2A1D3C7",
    x"2A1D153",
    x"2A1CEDF",
    x"2A1CC6B",
    x"2A1C9F8",
    x"2A1C786",
    x"2A1C515",
    x"2A1C2A4",
    x"2A1C033",
    x"2A1BDC4",
    x"2A1BB55",
    x"2A1B8E6",
    x"2A1B678",
    x"2A1B40B",
    x"2A1B19E",
    x"2A1AF32",
    x"2A1ACC6",
    x"2A1AA5C",
    x"2A1A7F1",
    x"2A1A588",
    x"2A1A31E",
    x"2A1A0B6",
    x"2A19E4E",
    x"2A19BE7",
    x"2A19980",
    x"2A1971A",
    x"2A194B5",
    x"2A19250",
    x"2A18FEB",
    x"2A18D88",
    x"2A18B25",
    x"2A188C2",
    x"2A18660",
    x"2A183FF",
    x"2A1819E",
    x"2A17F3E",
    x"2A17CDF",
    x"2A17A80",
    x"2A17821",
    x"2A175C4",
    x"2A17367",
    x"2A1710A",
    x"2A16EAE",
    x"2A16C53",
    x"2A169F8",
    x"2A1679E",
    x"2A16544",
    x"2A162EB",
    x"2A16093",
    x"2A15E3B",
    x"2A15BE3",
    x"2A1598D",
    x"2A15737",
    x"2A154E1",
    x"2A1528C",
    x"2A15038",
    x"2A14DE4",
    x"2A14B91",
    x"2A1493E",
    x"2A146EC",
    x"2A1449B",
    x"2A1424A",
    x"2A13FFA",
    x"2A13DAA",
    x"2A13B5B",
    x"2A1390C",
    x"2A136BE",
    x"2A13471",
    x"2A13224",
    x"2A12FD8",
    x"2A12D8C",
    x"2A12B41",
    x"2A128F7",
    x"2A126AD",
    x"2A12463",
    x"2A1221A",
    x"2A11FD2",
    x"2A11D8B",
    x"2A11B43",
    x"2A118FD",
    x"2A116B7",
    x"2A11472",
    x"2A1122D",
    x"2A10FE9",
    x"2A10DA5",
    x"2A10B62",
    x"2A1091F",
    x"2A106DD",
    x"2A1049C",
    x"2A1025B",
    x"2A1001B",
    x"2A0FDDB",
    x"2A0FB9C",
    x"2A0F95D",
    x"2A0F71F",
    x"2A0F4E1",
    x"2A0F2A4",
    x"2A0F068",
    x"2A0EE2C",
    x"2A0EBF1",
    x"2A0E9B6",
    x"2A0E77C",
    x"2A0E543",
    x"2A0E309",
    x"2A0E0D1",
    x"2A0DE99",
    x"2A0DC62",
    x"2A0DA2B",
    x"2A0D7F5",
    x"2A0D5BF",
    x"2A0D38A",
    x"2A0D155",
    x"2A0CF21",
    x"2A0CCEE",
    x"2A0CABB",
    x"2A0C888",
    x"2A0C656",
    x"2A0C425",
    x"2A0C1F4",
    x"2A0BFC4",
    x"2A0BD94",
    x"2A0BB65",
    x"2A0B937",
    x"2A0B709",
    x"2A0B4DB",
    x"2A0B2AE",
    x"2A0B082",
    x"2A0AE56",
    x"2A0AC2B",
    x"2A0AA00",
    x"2A0A7D6",
    x"2A0A5AC",
    x"2A0A383",
    x"2A0A15A",
    x"2A09F32",
    x"2A09D0B",
    x"2A09AE4",
    x"2A098BD",
    x"2A09697",
    x"2A09472",
    x"2A0924D",
    x"2A09029",
    x"2A08E05",
    x"2A08BE2",
    x"2A089BF",
    x"2A0879D",
    x"2A0857B",
    x"2A0835A",
    x"2A0813A",
    x"2A07F19",
    x"2A07CFA",
    x"2A07ADB",
    x"2A078BD",
    x"2A0769F",
    x"2A07481",
    x"2A07264",
    x"2A07048",
    x"2A06E2C",
    x"2A06C11",
    x"2A069F6",
    x"2A067DC",
    x"2A065C2",
    x"2A063A9",
    x"2A06190",
    x"2A05F78",
    x"2A05D61",
    x"2A05B4A",
    x"2A05933",
    x"2A0571D",
    x"2A05508",
    x"2A052F3",
    x"2A050DE",
    x"2A04ECA",
    x"2A04CB7",
    x"2A04AA4",
    x"2A04891",
    x"2A0467F",
    x"2A0446E",
    x"2A0425D",
    x"2A0404D",
    x"2A03E3D",
    x"2A03C2E",
    x"2A03A1F",
    x"2A03811",
    x"2A03603",
    x"2A033F6",
    x"2A031E9",
    x"2A02FDD",
    x"2A02DD1",
    x"2A02BC6",
    x"2A029BB",
    x"2A027B1",
    x"2A025A7",
    x"2A0239E",
    x"2A02195",
    x"2A01F8D",
    x"2A01D86",
    x"2A01B7F",
    x"2A01978",
    x"2A01772",
    x"2A0156C",
    x"2A01367",
    x"2A01163",
    x"2A00F5E",
    x"2A00D5B",
    x"2A00B58",
    x"2A00955",
    x"2A00753",
    x"2A00552",
    x"2A00350",
    x"2A00150",
    x"29FFEA0",
    x"29FFAA1",
    x"29FF6A3",
    x"29FF2A6",
    x"29FEEA9",
    x"29FEAAE",
    x"29FE6B4",
    x"29FE2BB",
    x"29FDEC3",
    x"29FDACB",
    x"29FD6D5",
    x"29FD2E0",
    x"29FCEEC",
    x"29FCAF9",
    x"29FC706",
    x"29FC315",
    x"29FBF25",
    x"29FBB35",
    x"29FB747",
    x"29FB35A",
    x"29FAF6E",
    x"29FAB82",
    x"29FA798",
    x"29FA3AE",
    x"29F9FC6",
    x"29F9BDE",
    x"29F97F8",
    x"29F9412",
    x"29F902E",
    x"29F8C4A",
    x"29F8868",
    x"29F8486",
    x"29F80A6",
    x"29F7CC6",
    x"29F78E7",
    x"29F7509",
    x"29F712D",
    x"29F6D51",
    x"29F6976",
    x"29F659C",
    x"29F61C3",
    x"29F5DEB",
    x"29F5A14",
    x"29F563E",
    x"29F5269",
    x"29F4E95",
    x"29F4AC2",
    x"29F46F0",
    x"29F431E",
    x"29F3F4E",
    x"29F3B7F",
    x"29F37B0",
    x"29F33E3",
    x"29F3016",
    x"29F2C4B",
    x"29F2880",
    x"29F24B7",
    x"29F20EE",
    x"29F1D26",
    x"29F195F",
    x"29F1599",
    x"29F11D4",
    x"29F0E10",
    x"29F0A4D",
    x"29F068B",
    x"29F02CA",
    x"29EFF0A",
    x"29EFB4B",
    x"29EF78C",
    x"29EF3CF",
    x"29EF012",
    x"29EEC57",
    x"29EE89C",
    x"29EE4E2",
    x"29EE12A",
    x"29EDD72",
    x"29ED9BB",
    x"29ED605",
    x"29ED250",
    x"29ECE9C",
    x"29ECAE9",
    x"29EC736",
    x"29EC385",
    x"29EBFD5",
    x"29EBC25",
    x"29EB877",
    x"29EB4C9",
    x"29EB11C",
    x"29EAD70",
    x"29EA9C5",
    x"29EA61B",
    x"29EA272",
    x"29E9ECA",
    x"29E9B23",
    x"29E977D",
    x"29E93D7",
    x"29E9033",
    x"29E8C8F",
    x"29E88EC",
    x"29E854B",
    x"29E81AA",
    x"29E7E0A",
    x"29E7A6B",
    x"29E76CD",
    x"29E732F",
    x"29E6F93",
    x"29E6BF8",
    x"29E685D",
    x"29E64C3",
    x"29E612B",
    x"29E5D93",
    x"29E59FC",
    x"29E5666",
    x"29E52D1",
    x"29E4F3C",
    x"29E4BA9",
    x"29E4817",
    x"29E4485",
    x"29E40F4",
    x"29E3D65",
    x"29E39D6",
    x"29E3648",
    x"29E32BB",
    x"29E2F2E",
    x"29E2BA3",
    x"29E2818",
    x"29E248F",
    x"29E2106",
    x"29E1D7E",
    x"29E19F7",
    x"29E1671",
    x"29E12EC",
    x"29E0F68",
    x"29E0BE5",
    x"29E0862",
    x"29E04E0",
    x"29E0160",
    x"29DFDE0",
    x"29DFA61",
    x"29DF6E2",
    x"29DF365",
    x"29DEFE9",
    x"29DEC6D",
    x"29DE8F3",
    x"29DE579",
    x"29DE200",
    x"29DDE88",
    x"29DDB11",
    x"29DD79A",
    x"29DD425",
    x"29DD0B0",
    x"29DCD3C",
    x"29DC9CA",
    x"29DC657",
    x"29DC2E6",
    x"29DBF76",
    x"29DBC07",
    x"29DB898",
    x"29DB52A",
    x"29DB1BD",
    x"29DAE51",
    x"29DAAE6",
    x"29DA77C",
    x"29DA413",
    x"29DA0AA",
    x"29D9D42",
    x"29D99DB",
    x"29D9675",
    x"29D9310",
    x"29D8FAC",
    x"29D8C48",
    x"29D88E6",
    x"29D8584",
    x"29D8223",
    x"29D7EC3",
    x"29D7B63",
    x"29D7805",
    x"29D74A7",
    x"29D714B",
    x"29D6DEF",
    x"29D6A94",
    x"29D673A",
    x"29D63E0",
    x"29D6088",
    x"29D5D30",
    x"29D59D9",
    x"29D5683",
    x"29D532E",
    x"29D4FD9",
    x"29D4C86",
    x"29D4933",
    x"29D45E1",
    x"29D4290",
    x"29D3F40",
    x"29D3BF1",
    x"29D38A2",
    x"29D3554",
    x"29D3207",
    x"29D2EBB",
    x"29D2B70",
    x"29D2825",
    x"29D24DC",
    x"29D2193",
    x"29D1E4B",
    x"29D1B04",
    x"29D17BE",
    x"29D1478",
    x"29D1133",
    x"29D0DEF",
    x"29D0AAC",
    x"29D076A",
    x"29D0429",
    x"29D00E8",
    x"29CFDA8",
    x"29CFA69",
    x"29CF72B",
    x"29CF3EE",
    x"29CF0B1",
    x"29CED75",
    x"29CEA3A",
    x"29CE700",
    x"29CE3C7",
    x"29CE08E",
    x"29CDD56",
    x"29CDA20",
    x"29CD6E9",
    x"29CD3B4",
    x"29CD080",
    x"29CCD4C",
    x"29CCA19",
    x"29CC6E7",
    x"29CC3B5",
    x"29CC085",
    x"29CBD55",
    x"29CBA26",
    x"29CB6F8",
    x"29CB3CB",
    x"29CB09E",
    x"29CAD72",
    x"29CAA48",
    x"29CA71D",
    x"29CA3F4",
    x"29CA0CB",
    x"29C9DA4",
    x"29C9A7D",
    x"29C9756",
    x"29C9431",
    x"29C910C",
    x"29C8DE8",
    x"29C8AC5",
    x"29C87A3",
    x"29C8481",
    x"29C8161",
    x"29C7E41",
    x"29C7B22",
    x"29C7803",
    x"29C74E6",
    x"29C71C9",
    x"29C6EAD",
    x"29C6B91",
    x"29C6877",
    x"29C655D",
    x"29C6244",
    x"29C5F2C",
    x"29C5C15",
    x"29C58FE",
    x"29C55E8",
    x"29C52D3",
    x"29C4FBF",
    x"29C4CAB",
    x"29C4998",
    x"29C4686",
    x"29C4375",
    x"29C4065",
    x"29C3D55",
    x"29C3A46",
    x"29C3738",
    x"29C342A",
    x"29C311E",
    x"29C2E12",
    x"29C2B07",
    x"29C27FC",
    x"29C24F3",
    x"29C21EA",
    x"29C1EE2",
    x"29C1BDA",
    x"29C18D4",
    x"29C15CE",
    x"29C12C9",
    x"29C0FC5",
    x"29C0CC1",
    x"29C09BE",
    x"29C06BC",
    x"29C03BB",
    x"29C00BA",
    x"29BFDBA",
    x"29BFABB",
    x"29BF7BD",
    x"29BF4C0",
    x"29BF1C3",
    x"29BEEC7",
    x"29BEBCB",
    x"29BE8D1",
    x"29BE5D7",
    x"29BE2DE",
    x"29BDFE5",
    x"29BDCEE",
    x"29BD9F7",
    x"29BD701",
    x"29BD40C",
    x"29BD117",
    x"29BCE23",
    x"29BCB30",
    x"29BC83D",
    x"29BC54C",
    x"29BC25B",
    x"29BBF6A",
    x"29BBC7B",
    x"29BB98C",
    x"29BB69E",
    x"29BB3B1",
    x"29BB0C4",
    x"29BADD9",
    x"29BAAED",
    x"29BA803",
    x"29BA519",
    x"29BA231",
    x"29B9F48",
    x"29B9C61",
    x"29B997A",
    x"29B9694",
    x"29B93AF",
    x"29B90CA",
    x"29B8DE6",
    x"29B8B03",
    x"29B8821",
    x"29B853F",
    x"29B825E",
    x"29B7F7E",
    x"29B7C9F",
    x"29B79C0",
    x"29B76E2",
    x"29B7404",
    x"29B7128",
    x"29B6E4C",
    x"29B6B71",
    x"29B6896",
    x"29B65BC",
    x"29B62E3",
    x"29B600B",
    x"29B5D33",
    x"29B5A5C",
    x"29B5786",
    x"29B54B0",
    x"29B51DC",
    x"29B4F08",
    x"29B4C34",
    x"29B4961",
    x"29B468F",
    x"29B43BE",
    x"29B40EE",
    x"29B3E1E",
    x"29B3B4F",
    x"29B3880",
    x"29B35B2",
    x"29B32E5",
    x"29B3019",
    x"29B2D4D",
    x"29B2A82",
    x"29B27B8",
    x"29B24EE",
    x"29B2225",
    x"29B1F5D",
    x"29B1C96",
    x"29B19CF",
    x"29B1709",
    x"29B1443",
    x"29B117F",
    x"29B0EBB",
    x"29B0BF7",
    x"29B0935",
    x"29B0673",
    x"29B03B1",
    x"29B00F1",
    x"29AFE31",
    x"29AFB72",
    x"29AF8B3",
    x"29AF5F5",
    x"29AF338",
    x"29AF07C",
    x"29AEDC0",
    x"29AEB05",
    x"29AE84B",
    x"29AE591",
    x"29AE2D8",
    x"29AE01F",
    x"29ADD68",
    x"29ADAB1",
    x"29AD7FA",
    x"29AD545",
    x"29AD290",
    x"29ACFDB",
    x"29ACD28",
    x"29ACA75",
    x"29AC7C3",
    x"29AC511",
    x"29AC260",
    x"29ABFB0",
    x"29ABD00",
    x"29ABA51",
    x"29AB7A3",
    x"29AB4F5",
    x"29AB249",
    x"29AAF9C",
    x"29AACF1",
    x"29AAA46",
    x"29AA79C",
    x"29AA4F2",
    x"29AA249",
    x"29A9FA1",
    x"29A9CF9",
    x"29A9A52",
    x"29A97AC",
    x"29A9507",
    x"29A9262",
    x"29A8FBD",
    x"29A8D1A",
    x"29A8A77",
    x"29A87D4",
    x"29A8533",
    x"29A8292",
    x"29A7FF2",
    x"29A7D52",
    x"29A7AB3",
    x"29A7815",
    x"29A7577",
    x"29A72DA",
    x"29A703D",
    x"29A6DA2",
    x"29A6B07",
    x"29A686C",
    x"29A65D2",
    x"29A6339",
    x"29A60A1",
    x"29A5E09",
    x"29A5B72",
    x"29A58DB",
    x"29A5645",
    x"29A53B0",
    x"29A511C",
    x"29A4E88",
    x"29A4BF4",
    x"29A4962",
    x"29A46D0",
    x"29A443E",
    x"29A41AD",
    x"29A3F1D",
    x"29A3C8E",
    x"29A39FF",
    x"29A3771",
    x"29A34E3",
    x"29A3256",
    x"29A2FCA",
    x"29A2D3F",
    x"29A2AB4",
    x"29A2829",
    x"29A259F",
    x"29A2316",
    x"29A208E",
    x"29A1E06",
    x"29A1B7F",
    x"29A18F8",
    x"29A1672",
    x"29A13ED",
    x"29A1168",
    x"29A0EE4",
    x"29A0C61",
    x"29A09DE",
    x"29A075C",
    x"29A04DB",
    x"29A025A",
    x"299FFD9",
    x"299FD5A",
    x"299FADB",
    x"299F85C",
    x"299F5DF",
    x"299F361",
    x"299F0E5",
    x"299EE69",
    x"299EBEE",
    x"299E973",
    x"299E6F9",
    x"299E47F",
    x"299E207",
    x"299DF8E",
    x"299DD17",
    x"299DAA0",
    x"299D82A",
    x"299D5B4",
    x"299D33F",
    x"299D0CA",
    x"299CE56",
    x"299CBE3",
    x"299C970",
    x"299C6FE",
    x"299C48D",
    x"299C21C",
    x"299BFAC",
    x"299BD3C",
    x"299BACD",
    x"299B85F",
    x"299B5F1",
    x"299B384",
    x"299B117",
    x"299AEAB",
    x"299AC40",
    x"299A9D5",
    x"299A76B",
    x"299A501",
    x"299A298",
    x"299A030",
    x"2999DC8",
    x"2999B61",
    x"29998FB",
    x"2999695",
    x"299942F",
    x"29991CB",
    x"2998F67",
    x"2998D03",
    x"2998AA0",
    x"299883E",
    x"29985DC",
    x"299837B",
    x"299811A",
    x"2997EBA",
    x"2997C5B",
    x"29979FC",
    x"299779E",
    x"2997540",
    x"29972E3",
    x"2997087",
    x"2996E2B",
    x"2996BD0",
    x"2996975",
    x"299671B",
    x"29964C1",
    x"2996269",
    x"2996010",
    x"2995DB8",
    x"2995B61",
    x"299590B",
    x"29956B5",
    x"299545F",
    x"299520B",
    x"2994FB6",
    x"2994D63",
    x"2994B10",
    x"29948BD",
    x"299466B",
    x"299441A",
    x"29941C9",
    x"2993F79",
    x"2993D2A",
    x"2993ADB",
    x"299388C",
    x"299363E",
    x"29933F1",
    x"29931A4",
    x"2992F58",
    x"2992D0D",
    x"2992AC2",
    x"2992877",
    x"299262D",
    x"29923E4",
    x"299219B",
    x"2991F53",
    x"2991D0C",
    x"2991AC5",
    x"299187E",
    x"2991639",
    x"29913F3",
    x"29911AF",
    x"2990F6A",
    x"2990D27",
    x"2990AE4",
    x"29908A1",
    x"2990660",
    x"299041E",
    x"29901DE",
    x"298FF9D",
    x"298FD5E",
    x"298FB1F",
    x"298F8E0",
    x"298F6A2",
    x"298F465",
    x"298F228",
    x"298EFEC",
    x"298EDB0",
    x"298EB75",
    x"298E93A",
    x"298E700",
    x"298E4C7",
    x"298E28E",
    x"298E056",
    x"298DE1E",
    x"298DBE7",
    x"298D9B0",
    x"298D77A",
    x"298D544",
    x"298D30F",
    x"298D0DB",
    x"298CEA7",
    x"298CC73",
    x"298CA40",
    x"298C80E",
    x"298C5DC",
    x"298C3AB",
    x"298C17B",
    x"298BF4A",
    x"298BD1B",
    x"298BAEC",
    x"298B8BD",
    x"298B68F",
    x"298B462",
    x"298B235",
    x"298B009",
    x"298ADDD",
    x"298ABB2",
    x"298A987",
    x"298A75D",
    x"298A534",
    x"298A30B",
    x"298A0E2",
    x"2989EBA",
    x"2989C93",
    x"2989A6C",
    x"2989846",
    x"2989620",
    x"29893FB",
    x"29891D6",
    x"2988FB2",
    x"2988D8E",
    x"2988B6B",
    x"2988948",
    x"2988726",
    x"2988505",
    x"29882E4",
    x"29880C3",
    x"2987EA3",
    x"2987C84",
    x"2987A65",
    x"2987847",
    x"2987629",
    x"298740C",
    x"29871EF",
    x"2986FD3",
    x"2986DB7",
    x"2986B9C",
    x"2986981",
    x"2986767",
    x"298654E",
    x"2986334",
    x"298611C",
    x"2985F04",
    x"2985CEC",
    x"2985AD5",
    x"29858BF",
    x"29856A9",
    x"2985494",
    x"298527F",
    x"298506A",
    x"2984E57",
    x"2984C43",
    x"2984A30",
    x"298481E",
    x"298460C",
    x"29843FB",
    x"29841EA",
    x"2983FDA",
    x"2983DCA",
    x"2983BBB",
    x"29839AD",
    x"298379E",
    x"2983591",
    x"2983384",
    x"2983177",
    x"2982F6B",
    x"2982D5F",
    x"2982B54",
    x"298294A",
    x"2982740",
    x"2982536",
    x"298232D",
    x"2982124",
    x"2981F1C",
    x"2981D15",
    x"2981B0E",
    x"2981907",
    x"2981701",
    x"29814FC",
    x"29812F7",
    x"29810F2",
    x"2980EEE",
    x"2980CEB",
    x"2980AE8",
    x"29808E5",
    x"29806E3",
    x"29804E2",
    x"29802E1",
    x"29800E1",
    x"297FDC2",
    x"297F9C3",
    x"297F5C5",
    x"297F1C8",
    x"297EDCC",
    x"297E9D1",
    x"297E5D7",
    x"297E1DE",
    x"297DDE6",
    x"297D9EF",
    x"297D5F9",
    x"297D204",
    x"297CE10",
    x"297CA1D",
    x"297C62B",
    x"297C23A",
    x"297BE4A",
    x"297BA5B",
    x"297B66D",
    x"297B280",
    x"297AE93",
    x"297AAA8",
    x"297A6BE",
    x"297A2D5",
    x"2979EED",
    x"2979B05",
    x"297971F",
    x"297933A",
    x"2978F56",
    x"2978B72",
    x"2978790",
    x"29783AE",
    x"2977FCE",
    x"2977BEE",
    x"2977810",
    x"2977432",
    x"2977056",
    x"2976C7A",
    x"29768A0",
    x"29764C6",
    x"29760ED",
    x"2975D16",
    x"297593F",
    x"2975569",
    x"2975194",
    x"2974DC0",
    x"29749ED",
    x"297461B",
    x"297424A",
    x"2973E7A",
    x"2973AAB",
    x"29736DD",
    x"297330F",
    x"2972F43",
    x"2972B78",
    x"29727AD",
    x"29723E4",
    x"297201B",
    x"2971C54",
    x"297188D",
    x"29714C8",
    x"2971103",
    x"2970D3F",
    x"297097C",
    x"29705BA",
    x"29701F9",
    x"296FE39",
    x"296FA7A",
    x"296F6BC",
    x"296F2FF",
    x"296EF43",
    x"296EB87",
    x"296E7CD",
    x"296E413",
    x"296E05B",
    x"296DCA3",
    x"296D8ED",
    x"296D537",
    x"296D182",
    x"296CDCE",
    x"296CA1B",
    x"296C669",
    x"296C2B8",
    x"296BF08",
    x"296BB58",
    x"296B7AA",
    x"296B3FC",
    x"296B050",
    x"296ACA4",
    x"296A8FA",
    x"296A550",
    x"296A1A7",
    x"2969DFF",
    x"2969A58",
    x"29696B2",
    x"296930D",
    x"2968F68",
    x"2968BC5",
    x"2968822",
    x"2968481",
    x"29680E0",
    x"2967D40",
    x"29679A2",
    x"2967604",
    x"2967267",
    x"2966ECA",
    x"2966B2F",
    x"2966795",
    x"29663FB",
    x"2966063",
    x"2965CCB",
    x"2965934",
    x"296559F",
    x"296520A",
    x"2964E75",
    x"2964AE2",
    x"2964750",
    x"29643BF",
    x"296402E",
    x"2963C9F",
    x"2963910",
    x"2963582",
    x"29631F5",
    x"2962E69",
    x"2962ADE",
    x"2962754",
    x"29623CA",
    x"2962042",
    x"2961CBA",
    x"2961933",
    x"29615AE",
    x"2961229",
    x"2960EA4",
    x"2960B21",
    x"296079F",
    x"296041D",
    x"296009D",
    x"295FD1D",
    x"295F99E",
    x"295F620",
    x"295F2A3",
    x"295EF27",
    x"295EBAC",
    x"295E831",
    x"295E4B8",
    x"295E13F",
    x"295DDC7",
    x"295DA50",
    x"295D6DA",
    x"295D364",
    x"295CFF0",
    x"295CC7C",
    x"295C90A",
    x"295C598",
    x"295C227",
    x"295BEB7",
    x"295BB48",
    x"295B7D9",
    x"295B46C",
    x"295B0FF",
    x"295AD93",
    x"295AA28",
    x"295A6BE",
    x"295A355",
    x"2959FEC",
    x"2959C85",
    x"295991E",
    x"29595B8",
    x"2959253",
    x"2958EEF",
    x"2958B8C",
    x"2958829",
    x"29584C8",
    x"2958167",
    x"2957E07",
    x"2957AA8",
    x"295774A",
    x"29573EC",
    x"2957090",
    x"2956D34",
    x"29569D9",
    x"295667F",
    x"2956326",
    x"2955FCE",
    x"2955C76",
    x"295591F",
    x"29555C9",
    x"2955274",
    x"2954F20",
    x"2954BCD",
    x"295487A",
    x"2954529",
    x"29541D8",
    x"2953E88",
    x"2953B38",
    x"29537EA",
    x"295349D",
    x"2953150",
    x"2952E04",
    x"2952AB9",
    x"295276F",
    x"2952425",
    x"29520DC",
    x"2951D95",
    x"2951A4E",
    x"2951707",
    x"29513C2",
    x"295107E",
    x"2950D3A",
    x"29509F7",
    x"29506B5",
    x"2950374",
    x"2950033",
    x"294FCF4",
    x"294F9B5",
    x"294F677",
    x"294F339",
    x"294EFFD",
    x"294ECC1",
    x"294E987",
    x"294E64D",
    x"294E314",
    x"294DFDB",
    x"294DCA4",
    x"294D96D",
    x"294D637",
    x"294D302",
    x"294CFCD",
    x"294CC9A",
    x"294C967",
    x"294C635",
    x"294C304",
    x"294BFD4",
    x"294BCA4",
    x"294B975",
    x"294B647",
    x"294B31A",
    x"294AFEE",
    x"294ACC2",
    x"294A997",
    x"294A66D",
    x"294A344",
    x"294A01C",
    x"2949CF4",
    x"29499CD",
    x"29496A7",
    x"2949382",
    x"294905D",
    x"2948D3A",
    x"2948A17",
    x"29486F5",
    x"29483D3",
    x"29480B3",
    x"2947D93",
    x"2947A74",
    x"2947756",
    x"2947438",
    x"294711C",
    x"2946E00",
    x"2946AE5",
    x"29467CA",
    x"29464B1",
    x"2946198",
    x"2945E80",
    x"2945B69",
    x"2945852",
    x"294553D",
    x"2945228",
    x"2944F14",
    x"2944C00",
    x"29448EE",
    x"29445DC",
    x"29442CB",
    x"2943FBA",
    x"2943CAB",
    x"294399C",
    x"294368E",
    x"2943381",
    x"2943074",
    x"2942D68",
    x"2942A5D",
    x"2942753",
    x"294244A",
    x"2942141",
    x"2941E39",
    x"2941B32",
    x"294182C",
    x"2941526",
    x"2941221",
    x"2940F1D",
    x"2940C19",
    x"2940917",
    x"2940615",
    x"2940314",
    x"2940013",
    x"293FD14",
    x"293FA15",
    x"293F717",
    x"293F419",
    x"293F11D",
    x"293EE21",
    x"293EB26",
    x"293E82B",
    x"293E531",
    x"293E239",
    x"293DF40",
    x"293DC49",
    x"293D952",
    x"293D65C",
    x"293D367",
    x"293D073",
    x"293CD7F",
    x"293CA8C",
    x"293C79A",
    x"293C4A8",
    x"293C1B7",
    x"293BEC7",
    x"293BBD8",
    x"293B8E9",
    x"293B5FB",
    x"293B30E",
    x"293B022",
    x"293AD36",
    x"293AA4B",
    x"293A761",
    x"293A478",
    x"293A18F",
    x"2939EA7",
    x"2939BBF",
    x"29398D9",
    x"29395F3",
    x"293930E",
    x"2939029",
    x"2938D46",
    x"2938A63",
    x"2938781",
    x"293849F",
    x"29381BE",
    x"2937EDE",
    x"2937BFF",
    x"2937920",
    x"2937642",
    x"2937365",
    x"2937089",
    x"2936DAD",
    x"2936AD2",
    x"29367F7",
    x"293651E",
    x"2936245",
    x"2935F6D",
    x"2935C95",
    x"29359BE",
    x"29356E8",
    x"2935413",
    x"293513E",
    x"2934E6A",
    x"2934B97",
    x"29348C4",
    x"29345F3",
    x"2934322",
    x"2934051",
    x"2933D81",
    x"2933AB2",
    x"29337E4",
    x"2933516",
    x"2933249",
    x"2932F7D",
    x"2932CB2",
    x"29329E7",
    x"293271D",
    x"2932453",
    x"293218B",
    x"2931EC3",
    x"2931BFB",
    x"2931935",
    x"293166F",
    x"29313A9",
    x"29310E5",
    x"2930E21",
    x"2930B5E",
    x"293089B",
    x"29305D9",
    x"2930318",
    x"2930058",
    x"292FD98",
    x"292FAD9",
    x"292F81B",
    x"292F55D",
    x"292F2A0",
    x"292EFE4",
    x"292ED28",
    x"292EA6D",
    x"292E7B3",
    x"292E4F9",
    x"292E240",
    x"292DF88",
    x"292DCD1",
    x"292DA1A",
    x"292D764",
    x"292D4AE",
    x"292D1F9",
    x"292CF45",
    x"292CC92",
    x"292C9DF",
    x"292C72D",
    x"292C47B",
    x"292C1CA",
    x"292BF1A",
    x"292BC6B",
    x"292B9BC",
    x"292B70E",
    x"292B461",
    x"292B1B4",
    x"292AF08",
    x"292AC5C",
    x"292A9B2",
    x"292A707",
    x"292A45E",
    x"292A1B5",
    x"2929F0D",
    x"2929C66",
    x"29299BF",
    x"2929719",
    x"2929473",
    x"29291CF",
    x"2928F2A",
    x"2928C87",
    x"29289E4",
    x"2928742",
    x"29284A1",
    x"2928200",
    x"2927F60",
    x"2927CC0",
    x"2927A21",
    x"2927783",
    x"29274E5",
    x"2927249",
    x"2926FAC",
    x"2926D11",
    x"2926A76",
    x"29267DB",
    x"2926542",
    x"29262A9",
    x"2926011",
    x"2925D79",
    x"2925AE2",
    x"292584B",
    x"29255B6",
    x"2925321",
    x"292508C",
    x"2924DF8",
    x"2924B65",
    x"29248D3",
    x"2924641",
    x"29243AF",
    x"292411F",
    x"2923E8F",
    x"2923C00",
    x"2923971",
    x"29236E3",
    x"2923455",
    x"29231C9",
    x"2922F3D",
    x"2922CB1",
    x"2922A26",
    x"292279C",
    x"2922512",
    x"2922289",
    x"2922001",
    x"2921D79",
    x"2921AF2",
    x"292186C",
    x"29215E6",
    x"2921361",
    x"29210DC",
    x"2920E59",
    x"2920BD5",
    x"2920953",
    x"29206D1",
    x"292044F",
    x"29201CE",
    x"291FF4E",
    x"291FCCF",
    x"291FA50",
    x"291F7D2",
    x"291F554",
    x"291F2D7",
    x"291F05B",
    x"291EDDF",
    x"291EB64",
    x"291E8E9",
    x"291E66F",
    x"291E3F6",
    x"291E17D",
    x"291DF05",
    x"291DC8E",
    x"291DA17",
    x"291D7A1",
    x"291D52B",
    x"291D2B6",
    x"291D042",
    x"291CDCE",
    x"291CB5B",
    x"291C8E8",
    x"291C676",
    x"291C405",
    x"291C194",
    x"291BF24",
    x"291BCB5",
    x"291BA46",
    x"291B7D8",
    x"291B56A",
    x"291B2FD",
    x"291B090",
    x"291AE25",
    x"291ABB9",
    x"291A94F",
    x"291A6E5",
    x"291A47B",
    x"291A213",
    x"2919FAA",
    x"2919D43",
    x"2919ADC",
    x"2919875",
    x"291960F",
    x"29193AA",
    x"2919146",
    x"2918EE2",
    x"2918C7E",
    x"2918A1B",
    x"29187B9",
    x"2918557",
    x"29182F6",
    x"2918096",
    x"2917E36",
    x"2917BD7",
    x"2917978",
    x"291771A",
    x"29174BD",
    x"2917260",
    x"2917003",
    x"2916DA8",
    x"2916B4D",
    x"29168F2",
    x"2916698",
    x"291643F",
    x"29161E6",
    x"2915F8E",
    x"2915D36",
    x"2915ADF",
    x"2915889",
    x"2915633",
    x"29153DE",
    x"2915189",
    x"2914F35",
    x"2914CE1",
    x"2914A8F",
    x"291483C",
    x"29145EA",
    x"2914399",
    x"2914149",
    x"2913EF9",
    x"2913CA9",
    x"2913A5A",
    x"291380C",
    x"29135BE",
    x"2913371",
    x"2913124",
    x"2912ED8",
    x"2912C8D",
    x"2912A42",
    x"29127F8",
    x"29125AE",
    x"2912365",
    x"291211D",
    x"2911ED5",
    x"2911C8D",
    x"2911A46",
    x"2911800",
    x"29115BA",
    x"2911375",
    x"2911131",
    x"2910EED",
    x"2910CA9",
    x"2910A66",
    x"2910824",
    x"29105E2",
    x"29103A1",
    x"2910160",
    x"290FF20",
    x"290FCE1",
    x"290FAA2",
    x"290F863",
    x"290F626",
    x"290F3E8",
    x"290F1AC",
    x"290EF70",
    x"290ED34",
    x"290EAF9",
    x"290E8BE",
    x"290E685",
    x"290E44B",
    x"290E212",
    x"290DFDA",
    x"290DDA2",
    x"290DB6B",
    x"290D935",
    x"290D6FF",
    x"290D4C9",
    x"290D294",
    x"290D060",
    x"290CE2C",
    x"290CBF9",
    x"290C9C6",
    x"290C794",
    x"290C562",
    x"290C331",
    x"290C101",
    x"290BED1",
    x"290BCA1",
    x"290BA72",
    x"290B844",
    x"290B616",
    x"290B3E9",
    x"290B1BC",
    x"290AF90",
    x"290AD65",
    x"290AB3A",
    x"290A90F",
    x"290A6E5",
    x"290A4BC",
    x"290A293",
    x"290A06A",
    x"2909E42",
    x"2909C1B",
    x"29099F4",
    x"29097CE",
    x"29095A8",
    x"2909383",
    x"290915F",
    x"2908F3B",
    x"2908D17",
    x"2908AF4",
    x"29088D2",
    x"29086B0",
    x"290848E",
    x"290826D",
    x"290804D",
    x"2907E2D",
    x"2907C0E",
    x"29079EF",
    x"29077D1",
    x"29075B3",
    x"2907396",
    x"2907179",
    x"2906F5D",
    x"2906D42",
    x"2906B27",
    x"290690C",
    x"29066F2",
    x"29064D9",
    x"29062C0",
    x"29060A7",
    x"2905E8F",
    x"2905C78",
    x"2905A61",
    x"290584B",
    x"2905635",
    x"2905420",
    x"290520B",
    x"2904FF7",
    x"2904DE3",
    x"2904BD0",
    x"29049BD",
    x"29047AB",
    x"2904599",
    x"2904388",
    x"2904178",
    x"2903F67",
    x"2903D58",
    x"2903B49",
    x"290393A",
    x"290372C",
    x"290351F",
    x"2903312",
    x"2903105",
    x"2902EF9",
    x"2902CEE",
    x"2902AE3",
    x"29028D8",
    x"29026CE",
    x"29024C5",
    x"29022BC",
    x"29020B3",
    x"2901EAB",
    x"2901CA4",
    x"2901A9D",
    x"2901897",
    x"2901691",
    x"290148B",
    x"2901287",
    x"2901082",
    x"2900E7E",
    x"2900C7B",
    x"2900A78",
    x"2900876",
    x"2900674",
    x"2900472",
    x"2900272",
    x"2900071",
    x"28FFCE3",
    x"28FF8E5",
    x"28FF4E7",
    x"28FF0EA",
    x"28FECEE",
    x"28FE8F4",
    x"28FE4FA",
    x"28FE101",
    x"28FDD09",
    x"28FD913",
    x"28FD51D",
    x"28FD128",
    x"28FCD34",
    x"28FC941",
    x"28FC550",
    x"28FC15F",
    x"28FBD6F",
    x"28FB980",
    x"28FB592",
    x"28FB1A5",
    x"28FADB9",
    x"28FA9CE",
    x"28FA5E4",
    x"28FA1FB",
    x"28F9E13",
    x"28F9A2C",
    x"28F9646",
    x"28F9261",
    x"28F8E7D",
    x"28F8A9A",
    x"28F86B8",
    x"28F82D7",
    x"28F7EF6",
    x"28F7B17",
    x"28F7739",
    x"28F735C",
    x"28F6F7F",
    x"28F6BA4",
    x"28F67C9",
    x"28F63F0",
    x"28F6017",
    x"28F5C40",
    x"28F5869",
    x"28F5494",
    x"28F50BF",
    x"28F4CEB",
    x"28F4919",
    x"28F4547",
    x"28F4176",
    x"28F3DA6",
    x"28F39D7",
    x"28F3609",
    x"28F323C",
    x"28F2E70",
    x"28F2AA5",
    x"28F26DB",
    x"28F2311",
    x"28F1F49",
    x"28F1B82",
    x"28F17BB",
    x"28F13F6",
    x"28F1031",
    x"28F0C6E",
    x"28F08AB",
    x"28F04E9",
    x"28F0129",
    x"28EFD69",
    x"28EF9AA",
    x"28EF5EC",
    x"28EF22F",
    x"28EEE73",
    x"28EEAB8",
    x"28EE6FE",
    x"28EE344",
    x"28EDF8C",
    x"28EDBD5",
    x"28ED81E",
    x"28ED468",
    x"28ED0B4",
    x"28ECD00",
    x"28EC94D",
    x"28EC59B",
    x"28EC1EB",
    x"28EBE3B",
    x"28EBA8B",
    x"28EB6DD",
    x"28EB330",
    x"28EAF84",
    x"28EABD8",
    x"28EA82E",
    x"28EA484",
    x"28EA0DB",
    x"28E9D34",
    x"28E998D",
    x"28E95E7",
    x"28E9242",
    x"28E8E9E",
    x"28E8AFB",
    x"28E8758",
    x"28E83B7",
    x"28E8016",
    x"28E7C77",
    x"28E78D8",
    x"28E753A",
    x"28E719E",
    x"28E6E02",
    x"28E6A67",
    x"28E66CC",
    x"28E6333",
    x"28E5F9B",
    x"28E5C03",
    x"28E586D",
    x"28E54D7",
    x"28E5142",
    x"28E4DAF",
    x"28E4A1C",
    x"28E468A",
    x"28E42F8",
    x"28E3F68",
    x"28E3BD9",
    x"28E384A",
    x"28E34BC",
    x"28E3130",
    x"28E2DA4",
    x"28E2A19",
    x"28E268F",
    x"28E2306",
    x"28E1F7D",
    x"28E1BF6",
    x"28E186F",
    x"28E14EA",
    x"28E1165",
    x"28E0DE1",
    x"28E0A5E",
    x"28E06DC",
    x"28E035B",
    x"28DFFDA",
    x"28DFC5B",
    x"28DF8DC",
    x"28DF55E",
    x"28DF1E1",
    x"28DEE65",
    x"28DEAEA",
    x"28DE770",
    x"28DE3F6",
    x"28DE07E",
    x"28DDD06",
    x"28DD98F",
    x"28DD619",
    x"28DD2A4",
    x"28DCF30",
    x"28DCBBD",
    x"28DC84A",
    x"28DC4D8",
    x"28DC168",
    x"28DBDF8",
    x"28DBA89",
    x"28DB71A",
    x"28DB3AD",
    x"28DB041",
    x"28DACD5",
    x"28DA96A",
    x"28DA600",
    x"28DA297",
    x"28D9F2F",
    x"28D9BC8",
    x"28D9861",
    x"28D94FB",
    x"28D9197",
    x"28D8E33",
    x"28D8AD0",
    x"28D876D",
    x"28D840C",
    x"28D80AB",
    x"28D7D4B",
    x"28D79ED",
    x"28D768F",
    x"28D7331",
    x"28D6FD5",
    x"28D6C79",
    x"28D691F",
    x"28D65C5",
    x"28D626C",
    x"28D5F14",
    x"28D5BBC",
    x"28D5866",
    x"28D5510",
    x"28D51BB",
    x"28D4E67",
    x"28D4B14",
    x"28D47C2",
    x"28D4470",
    x"28D411F",
    x"28D3DD0",
    x"28D3A81",
    x"28D3732",
    x"28D33E5",
    x"28D3098",
    x"28D2D4D",
    x"28D2A02",
    x"28D26B8",
    x"28D236E",
    x"28D2026",
    x"28D1CDE",
    x"28D1997",
    x"28D1651",
    x"28D130C",
    x"28D0FC8",
    x"28D0C84",
    x"28D0942",
    x"28D0600",
    x"28D02BF",
    x"28CFF7E",
    x"28CFC3F",
    x"28CF900",
    x"28CF5C2",
    x"28CF285",
    x"28CEF49",
    x"28CEC0E",
    x"28CE8D3",
    x"28CE599",
    x"28CE260",
    x"28CDF28",
    x"28CDBF1",
    x"28CD8BA",
    x"28CD584",
    x"28CD24F",
    x"28CCF1B",
    x"28CCBE8",
    x"28CC8B5",
    x"28CC584",
    x"28CC253",
    x"28CBF22",
    x"28CBBF3",
    x"28CB8C4",
    x"28CB597",
    x"28CB26A",
    x"28CAF3D",
    x"28CAC12",
    x"28CA8E7",
    x"28CA5BE",
    x"28CA294",
    x"28C9F6C",
    x"28C9C45",
    x"28C991E",
    x"28C95F8",
    x"28C92D3",
    x"28C8FAF",
    x"28C8C8B",
    x"28C8969",
    x"28C8647",
    x"28C8325",
    x"28C8005",
    x"28C7CE5",
    x"28C79C7",
    x"28C76A8",
    x"28C738B",
    x"28C706F",
    x"28C6D53",
    x"28C6A38",
    x"28C671E",
    x"28C6404",
    x"28C60EC",
    x"28C5DD4",
    x"28C5ABD",
    x"28C57A7",
    x"28C5491",
    x"28C517C",
    x"28C4E68",
    x"28C4B55",
    x"28C4843",
    x"28C4531",
    x"28C4220",
    x"28C3F10",
    x"28C3C01",
    x"28C38F2",
    x"28C35E4",
    x"28C32D7",
    x"28C2FCB",
    x"28C2CBF",
    x"28C29B4",
    x"28C26AA",
    x"28C23A1",
    x"28C2098",
    x"28C1D91",
    x"28C1A8A",
    x"28C1783",
    x"28C147E",
    x"28C1179",
    x"28C0E75",
    x"28C0B72",
    x"28C086F",
    x"28C056E",
    x"28C026D",
    x"28BFF6C",
    x"28BFC6D",
    x"28BF96E",
    x"28BF670",
    x"28BF373",
    x"28BF077",
    x"28BED7B",
    x"28BEA80",
    x"28BE786",
    x"28BE48C",
    x"28BE193",
    x"28BDE9B",
    x"28BDBA4",
    x"28BD8AD",
    x"28BD5B8",
    x"28BD2C3",
    x"28BCFCE",
    x"28BCCDB",
    x"28BC9E8",
    x"28BC6F6",
    x"28BC404",
    x"28BC114",
    x"28BBE24",
    x"28BBB35",
    x"28BB846",
    x"28BB559",
    x"28BB26C",
    x"28BAF7F",
    x"28BAC94",
    x"28BA9A9",
    x"28BA6BF",
    x"28BA3D6",
    x"28BA0ED",
    x"28B9E05",
    x"28B9B1E",
    x"28B9838",
    x"28B9552",
    x"28B926D",
    x"28B8F89",
    x"28B8CA5",
    x"28B89C2",
    x"28B86E0",
    x"28B83FF",
    x"28B811E",
    x"28B7E3E",
    x"28B7B5F",
    x"28B7881",
    x"28B75A3",
    x"28B72C6",
    x"28B6FEA",
    x"28B6D0E",
    x"28B6A33",
    x"28B6759",
    x"28B647F",
    x"28B61A7",
    x"28B5ECF",
    x"28B5BF7",
    x"28B5921",
    x"28B564B",
    x"28B5375",
    x"28B50A1",
    x"28B4DCD",
    x"28B4AFA",
    x"28B4828",
    x"28B4556",
    x"28B4285",
    x"28B3FB5",
    x"28B3CE5",
    x"28B3A16",
    x"28B3748",
    x"28B347B",
    x"28B31AE",
    x"28B2EE2",
    x"28B2C16",
    x"28B294C",
    x"28B2682",
    x"28B23B8",
    x"28B20F0",
    x"28B1E28",
    x"28B1B61",
    x"28B189A",
    x"28B15D4",
    x"28B130F",
    x"28B104B",
    x"28B0D87",
    x"28B0AC4",
    x"28B0802",
    x"28B0540",
    x"28B027F",
    x"28AFFBF",
    x"28AFCFF",
    x"28AFA40",
    x"28AF782",
    x"28AF4C5",
    x"28AF208",
    x"28AEF4C",
    x"28AEC90",
    x"28AE9D5",
    x"28AE71B",
    x"28AE462",
    x"28AE1A9",
    x"28ADEF1",
    x"28ADC3A",
    x"28AD983",
    x"28AD6CD",
    x"28AD417",
    x"28AD163",
    x"28ACEAF",
    x"28ACBFB",
    x"28AC949",
    x"28AC697",
    x"28AC3E5",
    x"28AC135",
    x"28ABE85",
    x"28ABBD6",
    x"28AB927",
    x"28AB679",
    x"28AB3CC",
    x"28AB11F",
    x"28AAE73",
    x"28AABC8",
    x"28AA91D",
    x"28AA673",
    x"28AA3CA",
    x"28AA121",
    x"28A9E79",
    x"28A9BD2",
    x"28A992C",
    x"28A9686",
    x"28A93E0",
    x"28A913C",
    x"28A8E98",
    x"28A8BF4",
    x"28A8952",
    x"28A86B0",
    x"28A840E",
    x"28A816E",
    x"28A7ECE",
    x"28A7C2E",
    x"28A7990",
    x"28A76F1",
    x"28A7454",
    x"28A71B7",
    x"28A6F1B",
    x"28A6C80",
    x"28A69E5",
    x"28A674B",
    x"28A64B1",
    x"28A6218",
    x"28A5F80",
    x"28A5CE9",
    x"28A5A52",
    x"28A57BC",
    x"28A5526",
    x"28A5291",
    x"28A4FFD",
    x"28A4D69",
    x"28A4AD6",
    x"28A4844",
    x"28A45B2",
    x"28A4321",
    x"28A4090",
    x"28A3E00",
    x"28A3B71",
    x"28A38E3",
    x"28A3655",
    x"28A33C8",
    x"28A313B",
    x"28A2EAF",
    x"28A2C24",
    x"28A2999",
    x"28A270F",
    x"28A2485",
    x"28A21FC",
    x"28A1F74",
    x"28A1CED",
    x"28A1A66",
    x"28A17E0",
    x"28A155A",
    x"28A12D5",
    x"28A1050",
    x"28A0DCD",
    x"28A0B4A",
    x"28A08C7",
    x"28A0645",
    x"28A03C4",
    x"28A0143",
    x"289FEC3",
    x"289FC44",
    x"289F9C5",
    x"289F747",
    x"289F4CA",
    x"289F24D",
    x"289EFD0",
    x"289ED55",
    x"289EADA",
    x"289E85F",
    x"289E5E6",
    x"289E36C",
    x"289E0F4",
    x"289DE7C",
    x"289DC05",
    x"289D98E",
    x"289D718",
    x"289D4A2",
    x"289D22D",
    x"289CFB9",
    x"289CD46",
    x"289CAD3",
    x"289C860",
    x"289C5EE",
    x"289C37D",
    x"289C10D",
    x"289BE9D",
    x"289BC2D",
    x"289B9BF",
    x"289B750",
    x"289B4E3",
    x"289B276",
    x"289B00A",
    x"289AD9E",
    x"289AB33",
    x"289A8C8",
    x"289A65F",
    x"289A3F5",
    x"289A18D",
    x"2899F24",
    x"2899CBD",
    x"2899A56",
    x"28997F0",
    x"289958A",
    x"2899325",
    x"28990C1",
    x"2898E5D",
    x"2898BF9",
    x"2898997",
    x"2898735",
    x"28984D3",
    x"2898272",
    x"2898012",
    x"2897DB2",
    x"2897B53",
    x"28978F4",
    x"2897697",
    x"2897439",
    x"28971DC",
    x"2896F80",
    x"2896D25",
    x"2896ACA",
    x"289686F",
    x"2896615",
    x"28963BC",
    x"2896164",
    x"2895F0C",
    x"2895CB4",
    x"2895A5D",
    x"2895807",
    x"28955B1",
    x"289535C",
    x"2895107",
    x"2894EB4",
    x"2894C60",
    x"2894A0D",
    x"28947BB",
    x"2894569",
    x"2894318",
    x"28940C8",
    x"2893E78",
    x"2893C29",
    x"28939DA",
    x"289378C",
    x"289353E",
    x"28932F1",
    x"28930A5",
    x"2892E59",
    x"2892C0D",
    x"28929C3",
    x"2892779",
    x"289252F",
    x"28922E6",
    x"289209E",
    x"2891E56",
    x"2891C0E",
    x"28919C8",
    x"2891782",
    x"289153C",
    x"28912F7",
    x"28910B2",
    x"2890E6F",
    x"2890C2B",
    x"28909E8",
    x"28907A6",
    x"2890565",
    x"2890324",
    x"28900E3",
    x"288FEA3",
    x"288FC64",
    x"288FA25",
    x"288F7E7",
    x"288F5A9",
    x"288F36C",
    x"288F12F",
    x"288EEF3",
    x"288ECB8",
    x"288EA7D",
    x"288E843",
    x"288E609",
    x"288E3D0",
    x"288E197",
    x"288DF5F",
    x"288DD27",
    x"288DAF0",
    x"288D8BA",
    x"288D684",
    x"288D44E",
    x"288D21A",
    x"288CFE5",
    x"288CDB2",
    x"288CB7F",
    x"288C94C",
    x"288C71A",
    x"288C4E8",
    x"288C2B7",
    x"288C087",
    x"288BE57",
    x"288BC28",
    x"288B9F9",
    x"288B7CB",
    x"288B59D",
    x"288B370",
    x"288B143",
    x"288AF17",
    x"288ACEC",
    x"288AAC1",
    x"288A897",
    x"288A66D",
    x"288A443",
    x"288A21B",
    x"2889FF2",
    x"2889DCB",
    x"2889BA3",
    x"288997D",
    x"2889757",
    x"2889531",
    x"288930C",
    x"28890E8",
    x"2888EC4",
    x"2888CA0",
    x"2888A7D",
    x"288885B",
    x"2888639",
    x"2888418",
    x"28881F7",
    x"2887FD7",
    x"2887DB7",
    x"2887B98",
    x"2887979",
    x"288775B",
    x"288753E",
    x"2887321",
    x"2887104",
    x"2886EE8",
    x"2886CCD",
    x"2886AB2",
    x"2886897",
    x"288667D",
    x"2886464",
    x"288624B",
    x"2886033",
    x"2885E1B",
    x"2885C04",
    x"28859ED",
    x"28857D7",
    x"28855C1",
    x"28853AC",
    x"2885197",
    x"2884F83",
    x"2884D70",
    x"2884B5C",
    x"288494A",
    x"2884738",
    x"2884526",
    x"2884315",
    x"2884105",
    x"2883EF5",
    x"2883CE5",
    x"2883AD6",
    x"28838C8",
    x"28836BA",
    x"28834AC",
    x"28832A0",
    x"2883093",
    x"2882E87",
    x"2882C7C",
    x"2882A71",
    x"2882867",
    x"288265D",
    x"2882454",
    x"288224B",
    x"2882042",
    x"2881E3B",
    x"2881C33",
    x"2881A2C",
    x"2881826",
    x"2881620",
    x"288141B",
    x"2881216",
    x"2881012",
    x"2880E0E",
    x"2880C0B",
    x"2880A08",
    x"2880806",
    x"2880604",
    x"2880403",
    x"2880202",
    x"2880002",
    x"287FC05",
    x"287F806",
    x"287F409",
    x"287F00C",
    x"287EC11",
    x"287E816",
    x"287E41D",
    x"287E024",
    x"287DC2D",
    x"287D836",
    x"287D441",
    x"287D04C",
    x"287CC59",
    x"287C866",
    x"287C474",
    x"287C084",
    x"287BC94",
    x"287B8A5",
    x"287B4B8",
    x"287B0CB",
    x"287ACDF",
    x"287A8F5",
    x"287A50B",
    x"287A122",
    x"2879D3A",
    x"2879953",
    x"287956E",
    x"2879189",
    x"2878DA5",
    x"28789C2",
    x"28785E0",
    x"28781FF",
    x"2877E1F",
    x"2877A40",
    x"2877662",
    x"2877285",
    x"2876EA9",
    x"2876ACD",
    x"28766F3",
    x"287631A",
    x"2875F42",
    x"2875B6A",
    x"2875794",
    x"28753BF",
    x"2874FEA",
    x"2874C17",
    x"2874844",
    x"2874472",
    x"28740A2",
    x"2873CD2",
    x"2873903",
    x"2873536",
    x"2873169",
    x"2872D9D",
    x"28729D2",
    x"2872608",
    x"287223F",
    x"2871E77",
    x"2871AB0",
    x"28716EA",
    x"2871324",
    x"2870F60",
    x"2870B9D",
    x"28707DA",
    x"2870419",
    x"2870058",
    x"286FC98",
    x"286F8DA",
    x"286F51C",
    x"286F15F",
    x"286EDA3",
    x"286E9E8",
    x"286E62E",
    x"286E275",
    x"286DEBD",
    x"286DB06",
    x"286D750",
    x"286D39A",
    x"286CFE6",
    x"286CC32",
    x"286C880",
    x"286C4CE",
    x"286C11D",
    x"286BD6E",
    x"286B9BF",
    x"286B611",
    x"286B264",
    x"286AEB7",
    x"286AB0C",
    x"286A762",
    x"286A3B9",
    x"286A010",
    x"2869C69",
    x"28698C2",
    x"286951C",
    x"2869177",
    x"2868DD3",
    x"2868A30",
    x"286868E",
    x"28682ED",
    x"2867F4D",
    x"2867BAD",
    x"286780F",
    x"2867471",
    x"28670D5",
    x"2866D39",
    x"286699E",
    x"2866604",
    x"286626B",
    x"2865ED3",
    x"2865B3C",
    x"28657A5",
    x"2865410",
    x"286507B",
    x"2864CE8",
    x"2864955",
    x"28645C3",
    x"2864232",
    x"2863EA2",
    x"2863B13",
    x"2863784",
    x"28633F7",
    x"286306A",
    x"2862CDF",
    x"2862954",
    x"28625CA",
    x"2862241",
    x"2861EB9",
    x"2861B32",
    x"28617AB",
    x"2861426",
    x"28610A1",
    x"2860D1E",
    x"286099B",
    x"2860619",
    x"2860298",
    x"285FF17",
    x"285FB98",
    x"285F81A",
    x"285F49C",
    x"285F11F",
    x"285EDA3",
    x"285EA29",
    x"285E6AE",
    x"285E335",
    x"285DFBD",
    x"285DC45",
    x"285D8CF",
    x"285D559",
    x"285D1E4",
    x"285CE70",
    x"285CAFD",
    x"285C78A",
    x"285C419",
    x"285C0A8",
    x"285BD39",
    x"285B9CA",
    x"285B65C",
    x"285B2EF",
    x"285AF82",
    x"285AC17",
    x"285A8AC",
    x"285A543",
    x"285A1DA",
    x"2859E72",
    x"2859B0A",
    x"28597A4",
    x"285943F",
    x"28590DA",
    x"2858D76",
    x"2858A13",
    x"28586B1",
    x"2858350",
    x"2857FEF",
    x"2857C90",
    x"2857931",
    x"28575D3",
    x"2857276",
    x"2856F1A",
    x"2856BBF",
    x"2856864",
    x"285650B",
    x"28561B2",
    x"2855E5A",
    x"2855B03",
    x"28557AC",
    x"2855457",
    x"2855102",
    x"2854DAE",
    x"2854A5B",
    x"2854709",
    x"28543B8",
    x"2854067",
    x"2853D17",
    x"28539C9",
    x"285367B",
    x"285332D",
    x"2852FE1",
    x"2852C95",
    x"285294B",
    x"2852601",
    x"28522B8",
    x"2851F6F",
    x"2851C28",
    x"28518E1",
    x"285159B",
    x"2851257",
    x"2850F12",
    x"2850BCF",
    x"285088C",
    x"285054B",
    x"285020A",
    x"284FECA",
    x"284FB8A",
    x"284F84C",
    x"284F50E",
    x"284F1D1",
    x"284EE95",
    x"284EB5A",
    x"284E820",
    x"284E4E6",
    x"284E1AD",
    x"284DE75",
    x"284DB3E",
    x"284D808",
    x"284D4D2",
    x"284D19D",
    x"284CE69",
    x"284CB36",
    x"284C804",
    x"284C4D2",
    x"284C1A1",
    x"284BE71",
    x"284BB42",
    x"284B813",
    x"284B4E6",
    x"284B1B9",
    x"284AE8D",
    x"284AB62",
    x"284A837",
    x"284A50E",
    x"284A1E5",
    x"2849EBD",
    x"2849B95",
    x"284986F",
    x"2849549",
    x"2849224",
    x"2848F00",
    x"2848BDD",
    x"28488BA",
    x"2848598",
    x"2848277",
    x"2847F57",
    x"2847C38",
    x"2847919",
    x"28475FB",
    x"28472DE",
    x"2846FC2",
    x"2846CA6",
    x"284698B",
    x"2846671",
    x"2846358",
    x"2846040",
    x"2845D28",
    x"2845A11",
    x"28456FB",
    x"28453E6",
    x"28450D1",
    x"2844DBD",
    x"2844AAA",
    x"2844798",
    x"2844486",
    x"2844176",
    x"2843E66",
    x"2843B56",
    x"2843848",
    x"284353A",
    x"284322D",
    x"2842F21",
    x"2842C16",
    x"284290B",
    x"2842601",
    x"28422F8",
    x"2841FF0",
    x"2841CE8",
    x"28419E1",
    x"28416DB",
    x"28413D6",
    x"28410D1",
    x"2840DCE",
    x"2840ACA",
    x"28407C8",
    x"28404C7",
    x"28401C6",
    x"283FEC6",
    x"283FBC6",
    x"283F8C8",
    x"283F5CA",
    x"283F2CD",
    x"283EFD1",
    x"283ECD5",
    x"283E9DA",
    x"283E6E0",
    x"283E3E7",
    x"283E0EE",
    x"283DDF6",
    x"283DAFF",
    x"283D809",
    x"283D513",
    x"283D21E",
    x"283CF2A",
    x"283CC37",
    x"283C944",
    x"283C652",
    x"283C361",
    x"283C070",
    x"283BD81",
    x"283BA92",
    x"283B7A3",
    x"283B4B6",
    x"283B1C9",
    x"283AEDD",
    x"283ABF1",
    x"283A907",
    x"283A61D",
    x"283A334",
    x"283A04B",
    x"2839D64",
    x"2839A7D",
    x"2839796",
    x"28394B1",
    x"28391CC",
    x"2838EE8",
    x"2838C05",
    x"2838922",
    x"2838640",
    x"283835F",
    x"283807E",
    x"2837D9F",
    x"2837AC0",
    x"28377E1",
    x"2837504",
    x"2837227",
    x"2836F4B",
    x"2836C6F",
    x"2836994",
    x"28366BA",
    x"28363E1",
    x"2836108",
    x"2835E30",
    x"2835B59",
    x"2835883",
    x"28355AD",
    x"28352D8",
    x"2835004",
    x"2834D30",
    x"2834A5D",
    x"283478B",
    x"28344B9",
    x"28341E8",
    x"2833F18",
    x"2833C49",
    x"283397A",
    x"28336AC",
    x"28333DF",
    x"2833112",
    x"2832E46",
    x"2832B7B",
    x"28328B0",
    x"28325E7",
    x"283231E",
    x"2832055",
    x"2831D8D",
    x"2831AC6",
    x"2831800",
    x"283153A",
    x"2831275",
    x"2830FB1",
    x"2830CED",
    x"2830A2B",
    x"2830768",
    x"28304A7",
    x"28301E6",
    x"282FF26",
    x"282FC67",
    x"282F9A8",
    x"282F6EA",
    x"282F42C",
    x"282F170",
    x"282EEB4",
    x"282EBF8",
    x"282E93E",
    x"282E684",
    x"282E3CA",
    x"282E112",
    x"282DE5A",
    x"282DBA3",
    x"282D8EC",
    x"282D636",
    x"282D381",
    x"282D0CC",
    x"282CE18",
    x"282CB65",
    x"282C8B3",
    x"282C601",
    x"282C350",
    x"282C09F",
    x"282BDEF",
    x"282BB40",
    x"282B892",
    x"282B5E4",
    x"282B337",
    x"282B08A",
    x"282ADDF",
    x"282AB33",
    x"282A889",
    x"282A5DF",
    x"282A336",
    x"282A08E",
    x"2829DE6",
    x"2829B3F",
    x"2829898",
    x"28295F2",
    x"282934D",
    x"28290A9",
    x"2828E05",
    x"2828B62",
    x"28288BF",
    x"282861D",
    x"282837C",
    x"28280DC",
    x"2827E3C",
    x"2827B9C",
    x"28278FE",
    x"2827660",
    x"28273C3",
    x"2827126",
    x"2826E8A",
    x"2826BEF",
    x"2826954",
    x"28266BA",
    x"2826421",
    x"2826188",
    x"2825EF0",
    x"2825C59",
    x"28259C2",
    x"282572C",
    x"2825496",
    x"2825201",
    x"2824F6D",
    x"2824CDA",
    x"2824A47",
    x"28247B5",
    x"2824523",
    x"2824292",
    x"2824002",
    x"2823D72",
    x"2823AE3",
    x"2823855",
    x"28235C7",
    x"282333A",
    x"28230AD",
    x"2822E21",
    x"2822B96",
    x"282290C",
    x"2822682",
    x"28223F8",
    x"2822170",
    x"2821EE8",
    x"2821C60",
    x"28219D9",
    x"2821753",
    x"28214CE",
    x"2821249",
    x"2820FC5",
    x"2820D41",
    x"2820ABE",
    x"282083C",
    x"28205BA",
    x"2820339",
    x"28200B8",
    x"281FE38",
    x"281FBB9",
    x"281F93A",
    x"281F6BC",
    x"281F43F",
    x"281F1C2",
    x"281EF46",
    x"281ECCB",
    x"281EA50",
    x"281E7D6",
    x"281E55C",
    x"281E2E3",
    x"281E06A",
    x"281DDF3",
    x"281DB7B",
    x"281D905",
    x"281D68F",
    x"281D41A",
    x"281D1A5",
    x"281CF31",
    x"281CCBD",
    x"281CA4A",
    x"281C7D8",
    x"281C567",
    x"281C2F5",
    x"281C085",
    x"281BE15",
    x"281BBA6",
    x"281B937",
    x"281B6C9",
    x"281B45C",
    x"281B1EF",
    x"281AF83",
    x"281AD17",
    x"281AAAC",
    x"281A842",
    x"281A5D8",
    x"281A36F",
    x"281A107",
    x"2819E9F",
    x"2819C37",
    x"28199D1",
    x"281976A",
    x"2819505",
    x"28192A0",
    x"281903C",
    x"2818DD8",
    x"2818B75",
    x"2818912",
    x"28186B0",
    x"281844F",
    x"28181EE",
    x"2817F8E",
    x"2817D2E",
    x"2817ACF",
    x"2817871",
    x"2817613",
    x"28173B6",
    x"2817159",
    x"2816EFD",
    x"2816CA2",
    x"2816A47",
    x"28167EC",
    x"2816593",
    x"281633A",
    x"28160E1",
    x"2815E89",
    x"2815C32",
    x"28159DB",
    x"2815785",
    x"281552F",
    x"28152DA",
    x"2815086",
    x"2814E32",
    x"2814BDF",
    x"281498C",
    x"281473A",
    x"28144E9",
    x"2814298",
    x"2814047",
    x"2813DF7",
    x"2813BA8",
    x"281395A",
    x"281370C",
    x"28134BE",
    x"2813271",
    x"2813025",
    x"2812DD9",
    x"2812B8E",
    x"2812943",
    x"28126F9",
    x"28124B0",
    x"2812267",
    x"281201F",
    x"2811DD7",
    x"2811B90",
    x"2811949",
    x"2811703",
    x"28114BE",
    x"2811279",
    x"2811034",
    x"2810DF1",
    x"2810BAD",
    x"281096B",
    x"2810729",
    x"28104E7",
    x"28102A6",
    x"2810066",
    x"280FE26",
    x"280FBE7",
    x"280F9A8",
    x"280F76A",
    x"280F52C",
    x"280F2EF",
    x"280F0B3",
    x"280EE77",
    x"280EC3C",
    x"280EA01",
    x"280E7C7",
    x"280E58D",
    x"280E354",
    x"280E11B",
    x"280DEE3",
    x"280DCAC",
    x"280DA75",
    x"280D83F",
    x"280D609",
    x"280D3D4",
    x"280D19F",
    x"280CF6B",
    x"280CD37",
    x"280CB04",
    x"280C8D2",
    x"280C6A0",
    x"280C46E",
    x"280C23E",
    x"280C00D",
    x"280BDDE",
    x"280BBAE",
    x"280B980",
    x"280B752",
    x"280B524",
    x"280B2F7",
    x"280B0CB",
    x"280AE9F",
    x"280AC73",
    x"280AA48",
    x"280A81E",
    x"280A5F4",
    x"280A3CB",
    x"280A1A3",
    x"2809F7A",
    x"2809D53",
    x"2809B2C",
    x"2809905",
    x"28096DF",
    x"28094BA",
    x"2809295",
    x"2809070",
    x"2808E4D",
    x"2808C29",
    x"2808A07",
    x"28087E4",
    x"28085C3",
    x"28083A1",
    x"2808181",
    x"2807F61",
    x"2807D41",
    x"2807B22",
    x"2807904",
    x"28076E6",
    x"28074C8",
    x"28072AB",
    x"280708F",
    x"2806E73",
    x"2806C57",
    x"2806A3D",
    x"2806822",
    x"2806609",
    x"28063EF",
    x"28061D7",
    x"2805FBE",
    x"2805DA7",
    x"2805B90",
    x"2805979",
    x"2805763",
    x"280554D",
    x"2805338",
    x"2805124",
    x"2804F10",
    x"2804CFC",
    x"2804AE9",
    x"28048D7",
    x"28046C5",
    x"28044B3",
    x"28042A2",
    x"2804092",
    x"2803E82",
    x"2803C73",
    x"2803A64",
    x"2803856",
    x"2803648",
    x"280343A",
    x"280322E",
    x"2803021",
    x"2802E16",
    x"2802C0A",
    x"28029FF",
    x"28027F5",
    x"28025EC",
    x"28023E2",
    x"28021DA",
    x"2801FD1",
    x"2801DCA",
    x"2801BC2",
    x"28019BC",
    x"28017B6",
    x"28015B0",
    x"28013AB",
    x"28011A6",
    x"2800FA2",
    x"2800D9E",
    x"2800B9B",
    x"2800998",
    x"2800796",
    x"2800595",
    x"2800394",
    x"2800193",
    x"27FFF26",
    x"27FFB27",
    x"27FF728",
    x"27FF32B",
    x"27FEF2F",
    x"27FEB33",
    x"27FE739",
    x"27FE340",
    x"27FDF48",
    x"27FDB50",
    x"27FD75A",
    x"27FD365",
    x"27FCF70",
    x"27FCB7D",
    x"27FC78A",
    x"27FC399",
    x"27FBFA9",
    x"27FBBB9",
    x"27FB7CB",
    x"27FB3DD",
    x"27FAFF1",
    x"27FAC05",
    x"27FA81B",
    x"27FA431",
    x"27FA049",
    x"27F9C61",
    x"27F987B",
    x"27F9495",
    x"27F90B0",
    x"27F8CCD",
    x"27F88EA",
    x"27F8508",
    x"27F8127",
    x"27F7D48",
    x"27F7969",
    x"27F758B",
    x"27F71AE",
    x"27F6DD2",
    x"27F69F7",
    x"27F661D",
    x"27F6244",
    x"27F5E6C",
    x"27F5A95",
    x"27F56BF",
    x"27F52E9",
    x"27F4F15",
    x"27F4B42",
    x"27F4770",
    x"27F439E",
    x"27F3FCE",
    x"27F3BFE",
    x"27F3830",
    x"27F3462",
    x"27F3096",
    x"27F2CCA",
    x"27F28FF",
    x"27F2535",
    x"27F216D",
    x"27F1DA5",
    x"27F19DE",
    x"27F1618",
    x"27F1253",
    x"27F0E8F",
    x"27F0ACB",
    x"27F0709",
    x"27F0348",
    x"27EFF87",
    x"27EFBC8",
    x"27EF80A",
    x"27EF44C",
    x"27EF08F",
    x"27EECD4",
    x"27EE919",
    x"27EE55F",
    x"27EE1A6",
    x"27EDDEE",
    x"27EDA37",
    x"27ED681",
    x"27ED2CC",
    x"27ECF18",
    x"27ECB65",
    x"27EC7B2",
    x"27EC401",
    x"27EC050",
    x"27EBCA1",
    x"27EB8F2",
    x"27EB544",
    x"27EB197",
    x"27EADEB",
    x"27EAA40",
    x"27EA696",
    x"27EA2ED",
    x"27E9F45",
    x"27E9B9D",
    x"27E97F7",
    x"27E9451",
    x"27E90AD",
    x"27E8D09",
    x"27E8966",
    x"27E85C4",
    x"27E8223",
    x"27E7E83",
    x"27E7AE4",
    x"27E7746",
    x"27E73A8",
    x"27E700C",
    x"27E6C70",
    x"27E68D6",
    x"27E653C",
    x"27E61A3",
    x"27E5E0B",
    x"27E5A74",
    x"27E56DE",
    x"27E5349",
    x"27E4FB4",
    x"27E4C21",
    x"27E488E",
    x"27E44FD",
    x"27E416C",
    x"27E3DDC",
    x"27E3A4D",
    x"27E36BF",
    x"27E3331",
    x"27E2FA5",
    x"27E2C1A",
    x"27E288F",
    x"27E2505",
    x"27E217D",
    x"27E1DF5",
    x"27E1A6E",
    x"27E16E7",
    x"27E1362",
    x"27E0FDE",
    x"27E0C5A",
    x"27E08D8",
    x"27E0556",
    x"27E01D5",
    x"27DFE55",
    x"27DFAD6",
    x"27DF757",
    x"27DF3DA",
    x"27DF05D",
    x"27DECE2",
    x"27DE967",
    x"27DE5ED",
    x"27DE274",
    x"27DDEFC",
    x"27DDB85",
    x"27DD80E",
    x"27DD499",
    x"27DD124",
    x"27DCDB0",
    x"27DCA3D",
    x"27DC6CB",
    x"27DC35A",
    x"27DBFE9",
    x"27DBC7A",
    x"27DB90B",
    x"27DB59D",
    x"27DB230",
    x"27DAEC4",
    x"27DAB59",
    x"27DA7EE",
    x"27DA485",
    x"27DA11C",
    x"27D9DB4",
    x"27D9A4D",
    x"27D96E7",
    x"27D9382",
    x"27D901D",
    x"27D8CBA",
    x"27D8957",
    x"27D85F5",
    x"27D8294",
    x"27D7F34",
    x"27D7BD4",
    x"27D7876",
    x"27D7518",
    x"27D71BB",
    x"27D6E5F",
    x"27D6B04",
    x"27D67AA",
    x"27D6450",
    x"27D60F8",
    x"27D5DA0",
    x"27D5A49",
    x"27D56F3",
    x"27D539D",
    x"27D5049",
    x"27D4CF5",
    x"27D49A2",
    x"27D4650",
    x"27D42FF",
    x"27D3FAF",
    x"27D3C5F",
    x"27D3911",
    x"27D35C3",
    x"27D3276",
    x"27D2F2A",
    x"27D2BDE",
    x"27D2894",
    x"27D254A",
    x"27D2201",
    x"27D1EB9",
    x"27D1B72",
    x"27D182B",
    x"27D14E6",
    x"27D11A1",
    x"27D0E5D",
    x"27D0B1A",
    x"27D07D7",
    x"27D0496",
    x"27D0155",
    x"27CFE15",
    x"27CFAD6",
    x"27CF798",
    x"27CF45A",
    x"27CF11D",
    x"27CEDE2",
    x"27CEAA6",
    x"27CE76C",
    x"27CE433",
    x"27CE0FA",
    x"27CDDC2",
    x"27CDA8B",
    x"27CD755",
    x"27CD420",
    x"27CD0EB",
    x"27CCDB7",
    x"27CCA84",
    x"27CC752",
    x"27CC420",
    x"27CC0F0",
    x"27CBDC0",
    x"27CBA91",
    x"27CB763",
    x"27CB435",
    x"27CB109",
    x"27CADDD",
    x"27CAAB2",
    x"27CA787",
    x"27CA45E",
    x"27CA135",
    x"27C9E0D",
    x"27C9AE6",
    x"27C97C0",
    x"27C949A",
    x"27C9175",
    x"27C8E51",
    x"27C8B2E",
    x"27C880C",
    x"27C84EA",
    x"27C81C9",
    x"27C7EA9",
    x"27C7B8A",
    x"27C786C",
    x"27C754E",
    x"27C7231",
    x"27C6F15",
    x"27C6BF9",
    x"27C68DF",
    x"27C65C5",
    x"27C62AC",
    x"27C5F94",
    x"27C5C7C",
    x"27C5965",
    x"27C564F",
    x"27C533A",
    x"27C5026",
    x"27C4D12",
    x"27C49FF",
    x"27C46ED",
    x"27C43DC",
    x"27C40CB",
    x"27C3DBB",
    x"27C3AAC",
    x"27C379E",
    x"27C3491",
    x"27C3184",
    x"27C2E78",
    x"27C2B6D",
    x"27C2862",
    x"27C2558",
    x"27C224F",
    x"27C1F47",
    x"27C1C40",
    x"27C1939",
    x"27C1633",
    x"27C132E",
    x"27C102A",
    x"27C0D26",
    x"27C0A23",
    x"27C0721",
    x"27C041F",
    x"27C011F",
    x"27BFE1F",
    x"27BFB20",
    x"27BF821",
    x"27BF524",
    x"27BF227",
    x"27BEF2B",
    x"27BEC2F",
    x"27BE934",
    x"27BE63B",
    x"27BE341",
    x"27BE049",
    x"27BDD51",
    x"27BDA5A",
    x"27BD764",
    x"27BD46F",
    x"27BD17A",
    x"27BCE86",
    x"27BCB93",
    x"27BC8A0",
    x"27BC5AE",
    x"27BC2BD",
    x"27BBFCD",
    x"27BBCDD",
    x"27BB9EE",
    x"27BB700",
    x"27BB413",
    x"27BB126",
    x"27BAE3A",
    x"27BAB4F",
    x"27BA865",
    x"27BA57B",
    x"27BA292",
    x"27B9FAA",
    x"27B9CC2",
    x"27B99DB",
    x"27B96F5",
    x"27B9410",
    x"27B912B",
    x"27B8E47",
    x"27B8B64",
    x"27B8882",
    x"27B85A0",
    x"27B82BF",
    x"27B7FDE",
    x"27B7CFF",
    x"27B7A20",
    x"27B7742",
    x"27B7464",
    x"27B7188",
    x"27B6EAC",
    x"27B6BD0",
    x"27B68F6",
    x"27B661C",
    x"27B6343",
    x"27B606A",
    x"27B5D92",
    x"27B5ABB",
    x"27B57E5",
    x"27B550F",
    x"27B523A",
    x"27B4F66",
    x"27B4C93",
    x"27B49C0",
    x"27B46EE",
    x"27B441C",
    x"27B414C",
    x"27B3E7C",
    x"27B3BAD",
    x"27B38DE",
    x"27B3610",
    x"27B3343",
    x"27B3076",
    x"27B2DAB",
    x"27B2AE0",
    x"27B2815",
    x"27B254C",
    x"27B2283",
    x"27B1FBA",
    x"27B1CF3",
    x"27B1A2C",
    x"27B1766",
    x"27B14A0",
    x"27B11DB",
    x"27B0F17",
    x"27B0C54",
    x"27B0991",
    x"27B06CF",
    x"27B040E",
    x"27B014D",
    x"27AFE8D",
    x"27AFBCE",
    x"27AF90F",
    x"27AF651",
    x"27AF394",
    x"27AF0D7",
    x"27AEE1C",
    x"27AEB60",
    x"27AE8A6",
    x"27AE5EC",
    x"27AE333",
    x"27AE07A",
    x"27ADDC3",
    x"27ADB0C",
    x"27AD855",
    x"27AD59F",
    x"27AD2EA",
    x"27AD036",
    x"27ACD82",
    x"27ACACF",
    x"27AC81D",
    x"27AC56B",
    x"27AC2BA",
    x"27AC00A",
    x"27ABD5A",
    x"27ABAAB",
    x"27AB7FD",
    x"27AB54F",
    x"27AB2A2",
    x"27AAFF6",
    x"27AAD4A",
    x"27AAA9F",
    x"27AA7F5",
    x"27AA54B",
    x"27AA2A2",
    x"27A9FFA",
    x"27A9D52",
    x"27A9AAB",
    x"27A9805",
    x"27A955F",
    x"27A92BA",
    x"27A9016",
    x"27A8D72",
    x"27A8ACF",
    x"27A882D",
    x"27A858B",
    x"27A82EA",
    x"27A804A",
    x"27A7DAA",
    x"27A7B0B",
    x"27A786C",
    x"27A75CE",
    x"27A7331",
    x"27A7095",
    x"27A6DF9",
    x"27A6B5E",
    x"27A68C3",
    x"27A662A",
    x"27A6390",
    x"27A60F8",
    x"27A5E60",
    x"27A5BC9",
    x"27A5932",
    x"27A569C",
    x"27A5407",
    x"27A5172",
    x"27A4EDE",
    x"27A4C4A",
    x"27A49B8",
    x"27A4726",
    x"27A4494",
    x"27A4203",
    x"27A3F73",
    x"27A3CE4",
    x"27A3A55",
    x"27A37C6",
    x"27A3539",
    x"27A32AC",
    x"27A301F",
    x"27A2D94",
    x"27A2B09",
    x"27A287E",
    x"27A25F4",
    x"27A236B",
    x"27A20E3",
    x"27A1E5B",
    x"27A1BD4",
    x"27A194D",
    x"27A16C7",
    x"27A1442",
    x"27A11BD",
    x"27A0F39",
    x"27A0CB5",
    x"27A0A32",
    x"27A07B0",
    x"27A052E",
    x"27A02AD",
    x"27A002D",
    x"279FDAD",
    x"279FB2E",
    x"279F8B0",
    x"279F632",
    x"279F3B5",
    x"279F138",
    x"279EEBC",
    x"279EC41",
    x"279E9C6",
    x"279E74C",
    x"279E4D2",
    x"279E259",
    x"279DFE1",
    x"279DD69",
    x"279DAF2",
    x"279D87C",
    x"279D606",
    x"279D391",
    x"279D11C",
    x"279CEA8",
    x"279CC35",
    x"279C9C2",
    x"279C750",
    x"279C4DF",
    x"279C26E",
    x"279BFFD",
    x"279BD8E",
    x"279BB1F",
    x"279B8B0",
    x"279B642",
    x"279B3D5",
    x"279B168",
    x"279AEFC",
    x"279AC91",
    x"279AA26",
    x"279A7BC",
    x"279A552",
    x"279A2E9",
    x"279A081",
    x"2799E19",
    x"2799BB2",
    x"279994B",
    x"27996E5",
    x"2799480",
    x"279921B",
    x"2798FB7",
    x"2798D53",
    x"2798AF0",
    x"279888D",
    x"279862C",
    x"27983CA",
    x"279816A",
    x"2797F0A",
    x"2797CAA",
    x"2797A4B",
    x"27977ED",
    x"279758F",
    x"2797332",
    x"27970D6",
    x"2796E7A",
    x"2796C1F",
    x"27969C4",
    x"279676A",
    x"2796510",
    x"27962B7",
    x"279605F",
    x"2795E07",
    x"2795BB0",
    x"2795959",
    x"2795703",
    x"27954AE",
    x"2795259",
    x"2795004",
    x"2794DB1",
    x"2794B5E",
    x"279490B",
    x"27946B9",
    x"2794468",
    x"2794217",
    x"2793FC7",
    x"2793D77",
    x"2793B28",
    x"27938D9",
    x"279368B",
    x"279343E",
    x"27931F1",
    x"2792FA5",
    x"2792D5A",
    x"2792B0E",
    x"27928C4",
    x"279267A",
    x"2792431",
    x"27921E8",
    x"2791FA0",
    x"2791D58",
    x"2791B11",
    x"27918CB",
    x"2791685",
    x"279143F",
    x"27911FB",
    x"2790FB6",
    x"2790D73",
    x"2790B30",
    x"27908ED",
    x"27906AB",
    x"279046A",
    x"2790229",
    x"278FFE9",
    x"278FDA9",
    x"278FB6A",
    x"278F92B",
    x"278F6ED",
    x"278F4B0",
    x"278F273",
    x"278F037",
    x"278EDFB",
    x"278EBC0",
    x"278E985",
    x"278E74B",
    x"278E511",
    x"278E2D8",
    x"278E0A0",
    x"278DE68",
    x"278DC31",
    x"278D9FA",
    x"278D7C4",
    x"278D58E",
    x"278D359",
    x"278D124",
    x"278CEF0",
    x"278CCBD",
    x"278CA8A",
    x"278C858",
    x"278C626",
    x"278C3F5",
    x"278C1C4",
    x"278BF94",
    x"278BD64",
    x"278BB35",
    x"278B906",
    x"278B6D8",
    x"278B4AB",
    x"278B27E",
    x"278B052",
    x"278AE26",
    x"278ABFB",
    x"278A9D0",
    x"278A7A6",
    x"278A57C",
    x"278A353",
    x"278A12A",
    x"2789F02",
    x"2789CDB",
    x"2789AB4",
    x"278988E",
    x"2789668",
    x"2789442",
    x"278921E",
    x"2788FF9",
    x"2788DD6",
    x"2788BB2",
    x"2788990",
    x"278876E",
    x"278854C",
    x"278832B",
    x"278810A",
    x"2787EEA",
    x"2787CCB",
    x"2787AAC",
    x"278788E",
    x"2787670",
    x"2787452",
    x"2787236",
    x"2787019",
    x"2786DFE",
    x"2786BE2",
    x"27869C8",
    x"27867AD",
    x"2786594",
    x"278637B",
    x"2786162",
    x"2785F4A",
    x"2785D32",
    x"2785B1B",
    x"2785905",
    x"27856EF",
    x"27854D9",
    x"27852C4",
    x"27850B0",
    x"2784E9C",
    x"2784C89",
    x"2784A76",
    x"2784863",
    x"2784652",
    x"2784440",
    x"2784230",
    x"278401F",
    x"2783E0F",
    x"2783C00",
    x"27839F1",
    x"27837E3",
    x"27835D6",
    x"27833C8",
    x"27831BC",
    x"2782FAF",
    x"2782DA4",
    x"2782B99",
    x"278298E",
    x"2782784",
    x"278257A",
    x"2782371",
    x"2782168",
    x"2781F60",
    x"2781D59",
    x"2781B52",
    x"278194B",
    x"2781745",
    x"2781540",
    x"278133A",
    x"2781136",
    x"2780F32",
    x"2780D2E",
    x"2780B2B",
    x"2780929",
    x"2780727",
    x"2780525",
    x"2780324",
    x"2780124",
    x"277FE48",
    x"277FA48",
    x"277F64A",
    x"277F24D",
    x"277EE51",
    x"277EA56",
    x"277E65C",
    x"277E263",
    x"277DE6B",
    x"277DA74",
    x"277D67E",
    x"277D289",
    x"277CE94",
    x"277CAA1",
    x"277C6AF",
    x"277C2BE",
    x"277BECE",
    x"277BADE",
    x"277B6F0",
    x"277B303",
    x"277AF17",
    x"277AB2B",
    x"277A741",
    x"277A358",
    x"2779F6F",
    x"2779B88",
    x"27797A2",
    x"27793BC",
    x"2778FD8",
    x"2778BF4",
    x"2778812",
    x"2778430",
    x"2778050",
    x"2777C70",
    x"2777892",
    x"27774B4",
    x"27770D7",
    x"2776CFB",
    x"2776921",
    x"2776547",
    x"277616E",
    x"2775D96",
    x"27759BF",
    x"27755E9",
    x"2775214",
    x"2774E40",
    x"2774A6D",
    x"277469B",
    x"27742CA",
    x"2773EFA",
    x"2773B2A",
    x"277375C",
    x"277338F",
    x"2772FC2",
    x"2772BF7",
    x"277282C",
    x"2772463",
    x"277209A",
    x"2771CD2",
    x"277190C",
    x"2771546",
    x"2771181",
    x"2770DBD",
    x"27709FA",
    x"2770638",
    x"2770277",
    x"276FEB7",
    x"276FAF8",
    x"276F739",
    x"276F37C",
    x"276EFC0",
    x"276EC04",
    x"276E84A",
    x"276E490",
    x"276E0D7",
    x"276DD20",
    x"276D969",
    x"276D5B3",
    x"276D1FE",
    x"276CE4A",
    x"276CA97",
    x"276C6E5",
    x"276C333",
    x"276BF83",
    x"276BBD4",
    x"276B825",
    x"276B478",
    x"276B0CB",
    x"276AD1F",
    x"276A974",
    x"276A5CA",
    x"276A221",
    x"2769E79",
    x"2769AD2",
    x"276972C",
    x"2769387",
    x"2768FE2",
    x"2768C3F",
    x"276889C",
    x"27684FA",
    x"276815A",
    x"2767DBA",
    x"2767A1B",
    x"276767D",
    x"27672DF",
    x"2766F43",
    x"2766BA8",
    x"276680D",
    x"2766474",
    x"27660DB",
    x"2765D43",
    x"27659AD",
    x"2765617",
    x"2765281",
    x"2764EED",
    x"2764B5A",
    x"27647C8",
    x"2764436",
    x"27640A6",
    x"2763D16",
    x"2763987",
    x"27635F9",
    x"276326C",
    x"2762EE0",
    x"2762B55",
    x"27627CA",
    x"2762441",
    x"27620B8",
    x"2761D30",
    x"27619A9",
    x"2761623",
    x"276129E",
    x"2760F1A",
    x"2760B97",
    x"2760814",
    x"2760493",
    x"2760112",
    x"275FD92",
    x"275FA13",
    x"275F695",
    x"275F318",
    x"275EF9C",
    x"275EC20",
    x"275E8A6",
    x"275E52C",
    x"275E1B3",
    x"275DE3B",
    x"275DAC4",
    x"275D74E",
    x"275D3D8",
    x"275D064",
    x"275CCF0",
    x"275C97D",
    x"275C60B",
    x"275C29A",
    x"275BF2A",
    x"275BBBB",
    x"275B84C",
    x"275B4DE",
    x"275B172",
    x"275AE06",
    x"275AA9B",
    x"275A730",
    x"275A3C7",
    x"275A05F",
    x"2759CF7",
    x"2759990",
    x"275962A",
    x"27592C5",
    x"2758F61",
    x"2758BFD",
    x"275889B",
    x"2758539",
    x"27581D8",
    x"2757E78",
    x"2757B19",
    x"27577BB",
    x"275745D",
    x"2757100",
    x"2756DA5",
    x"2756A4A",
    x"27566EF",
    x"2756396",
    x"275603E",
    x"2755CE6",
    x"275598F",
    x"2755639",
    x"27552E4",
    x"2754F90",
    x"2754C3C",
    x"27548EA",
    x"2754598",
    x"2754247",
    x"2753EF7",
    x"2753BA7",
    x"2753859",
    x"275350B",
    x"27531BE",
    x"2752E72",
    x"2752B27",
    x"27527DD",
    x"2752493",
    x"275214A",
    x"2751E02",
    x"2751ABB",
    x"2751775",
    x"2751430",
    x"27510EB",
    x"2750DA7",
    x"2750A64",
    x"2750722",
    x"27503E1",
    x"27500A0",
    x"274FD60",
    x"274FA21",
    x"274F6E3",
    x"274F3A6",
    x"274F069",
    x"274ED2E",
    x"274E9F3",
    x"274E6B9",
    x"274E37F",
    x"274E047",
    x"274DD0F",
    x"274D9D8",
    x"274D6A2",
    x"274D36D",
    x"274D039",
    x"274CD05",
    x"274C9D2",
    x"274C6A0",
    x"274C36F",
    x"274C03E",
    x"274BD0F",
    x"274B9E0",
    x"274B6B2",
    x"274B385",
    x"274B058",
    x"274AD2C",
    x"274AA01",
    x"274A6D7",
    x"274A3AE",
    x"274A086",
    x"2749D5E",
    x"2749A37",
    x"2749711",
    x"27493EB",
    x"27490C7",
    x"2748DA3",
    x"2748A80",
    x"274875E",
    x"274843C",
    x"274811C",
    x"2747DFC",
    x"2747ADD",
    x"27477BE",
    x"27474A1",
    x"2747184",
    x"2746E68",
    x"2746B4D",
    x"2746832",
    x"2746519",
    x"2746200",
    x"2745EE8",
    x"2745BD0",
    x"27458BA",
    x"27455A4",
    x"274528F",
    x"2744F7B",
    x"2744C67",
    x"2744954",
    x"2744642",
    x"2744331",
    x"2744021",
    x"2743D11",
    x"2743A02",
    x"27436F4",
    x"27433E7",
    x"27430DA",
    x"2742DCE",
    x"2742AC3",
    x"27427B9",
    x"27424AF",
    x"27421A7",
    x"2741E9F",
    x"2741B97",
    x"2741891",
    x"274158B",
    x"2741286",
    x"2740F82",
    x"2740C7E",
    x"274097C",
    x"274067A",
    x"2740378",
    x"2740078",
    x"273FD78",
    x"273FA79",
    x"273F77B",
    x"273F47D",
    x"273F181",
    x"273EE85",
    x"273EB89",
    x"273E88F",
    x"273E595",
    x"273E29C",
    x"273DFA4",
    x"273DCAC",
    x"273D9B5",
    x"273D6BF",
    x"273D3CA",
    x"273D0D5",
    x"273CDE2",
    x"273CAEF",
    x"273C7FC",
    x"273C50B",
    x"273C21A",
    x"273BF2A",
    x"273BC3A",
    x"273B94B",
    x"273B65D",
    x"273B370",
    x"273B084",
    x"273AD98",
    x"273AAAD",
    x"273A7C3",
    x"273A4D9",
    x"273A1F0",
    x"2739F08",
    x"2739C21",
    x"273993A",
    x"2739654",
    x"273936F",
    x"273908A",
    x"2738DA7",
    x"2738AC4",
    x"27387E1",
    x"2738500",
    x"273821F",
    x"2737F3F",
    x"2737C5F",
    x"2737980",
    x"27376A2",
    x"27373C5",
    x"27370E8",
    x"2736E0D",
    x"2736B31",
    x"2736857",
    x"273657D",
    x"27362A4",
    x"2735FCC",
    x"2735CF4",
    x"2735A1D",
    x"2735747",
    x"2735472",
    x"273519D",
    x"2734EC9",
    x"2734BF6",
    x"2734923",
    x"2734651",
    x"2734380",
    x"27340AF",
    x"2733DDF",
    x"2733B10",
    x"2733842",
    x"2733574",
    x"27332A7",
    x"2732FDB",
    x"2732D0F",
    x"2732A44",
    x"273277A",
    x"27324B1",
    x"27321E8",
    x"2731F20",
    x"2731C58",
    x"2731992",
    x"27316CB",
    x"2731406",
    x"2731141",
    x"2730E7D",
    x"2730BBA",
    x"27308F8",
    x"2730636",
    x"2730375",
    x"27300B4",
    x"272FDF4",
    x"272FB35",
    x"272F877",
    x"272F5B9",
    x"272F2FC",
    x"272F03F",
    x"272ED84",
    x"272EAC9",
    x"272E80E",
    x"272E555",
    x"272E29C",
    x"272DFE3",
    x"272DD2C",
    x"272DA75",
    x"272D7BE",
    x"272D509",
    x"272D254",
    x"272CFA0",
    x"272CCEC",
    x"272CA39",
    x"272C787",
    x"272C4D5",
    x"272C224",
    x"272BF74",
    x"272BCC5",
    x"272BA16",
    x"272B768",
    x"272B4BA",
    x"272B20D",
    x"272AF61",
    x"272ACB6",
    x"272AA0B",
    x"272A761",
    x"272A4B7",
    x"272A20E",
    x"2729F66",
    x"2729CBF",
    x"2729A18",
    x"2729772",
    x"27294CC",
    x"2729227",
    x"2728F83",
    x"2728CDF",
    x"2728A3C",
    x"272879A",
    x"27284F9",
    x"2728258",
    x"2727FB8",
    x"2727D18",
    x"2727A79",
    x"27277DB",
    x"272753D",
    x"27272A0",
    x"2727004",
    x"2726D68",
    x"2726ACD",
    x"2726833",
    x"2726599",
    x"2726300",
    x"2726067",
    x"2725DD0",
    x"2725B38",
    x"27258A2",
    x"272560C",
    x"2725377",
    x"27250E2",
    x"2724E4F",
    x"2724BBB",
    x"2724929",
    x"2724697",
    x"2724405",
    x"2724175",
    x"2723EE5",
    x"2723C55",
    x"27239C6",
    x"2723738",
    x"27234AB",
    x"272321E",
    x"2722F92",
    x"2722D06",
    x"2722A7B",
    x"27227F1",
    x"2722567",
    x"27222DE",
    x"2722056",
    x"2721DCE",
    x"2721B47",
    x"27218C0",
    x"272163B",
    x"27213B5",
    x"2721131",
    x"2720EAD",
    x"2720C29",
    x"27209A7",
    x"2720725",
    x"27204A3",
    x"2720222",
    x"271FFA2",
    x"271FD22",
    x"271FAA3",
    x"271F825",
    x"271F5A7",
    x"271F32A",
    x"271F0AE",
    x"271EE32",
    x"271EBB7",
    x"271E93C",
    x"271E6C2",
    x"271E449",
    x"271E1D0",
    x"271DF58",
    x"271DCE0",
    x"271DA69",
    x"271D7F3",
    x"271D57D",
    x"271D308",
    x"271D094",
    x"271CE20",
    x"271CBAD",
    x"271C93A",
    x"271C6C8",
    x"271C457",
    x"271C1E6",
    x"271BF76",
    x"271BD06",
    x"271BA97",
    x"271B829",
    x"271B5BB",
    x"271B34E",
    x"271B0E2",
    x"271AE76",
    x"271AC0A",
    x"271A9A0",
    x"271A736",
    x"271A4CC",
    x"271A263",
    x"2719FFB",
    x"2719D93",
    x"2719B2C",
    x"27198C6",
    x"2719660",
    x"27193FA",
    x"2719196",
    x"2718F32",
    x"2718CCE",
    x"2718A6B",
    x"2718809",
    x"27185A7",
    x"2718346",
    x"27180E6",
    x"2717E86",
    x"2717C26",
    x"27179C8",
    x"2717769",
    x"271750C",
    x"27172AF",
    x"2717053",
    x"2716DF7",
    x"2716B9C",
    x"2716941",
    x"27166E7",
    x"271648D",
    x"2716235",
    x"2715FDC",
    x"2715D85",
    x"2715B2E",
    x"27158D7",
    x"2715681",
    x"271542C",
    x"27151D7",
    x"2714F83",
    x"2714D2F",
    x"2714ADC",
    x"271488A",
    x"2714638",
    x"27143E7",
    x"2714196",
    x"2713F46",
    x"2713CF6",
    x"2713AA8",
    x"2713859",
    x"271360B",
    x"27133BE",
    x"2713171",
    x"2712F25",
    x"2712CDA",
    x"2712A8F",
    x"2712845",
    x"27125FB",
    x"27123B2",
    x"2712169",
    x"2711F21",
    x"2711CD9",
    x"2711A92",
    x"271184C",
    x"2711606",
    x"27113C1",
    x"271117C",
    x"2710F38",
    x"2710CF5",
    x"2710AB2",
    x"2710870",
    x"271062E",
    x"27103EC",
    x"27101AC",
    x"270FF6C",
    x"270FD2C",
    x"270FAED",
    x"270F8AF",
    x"270F671",
    x"270F433",
    x"270F1F7",
    x"270EFBA",
    x"270ED7F",
    x"270EB44",
    x"270E909",
    x"270E6CF",
    x"270E496",
    x"270E25D",
    x"270E024",
    x"270DDED",
    x"270DBB5",
    x"270D97F",
    x"270D749",
    x"270D513",
    x"270D2DE",
    x"270D0AA",
    x"270CE76",
    x"270CC43",
    x"270CA10",
    x"270C7DE",
    x"270C5AC",
    x"270C37B",
    x"270C14A",
    x"270BF1A",
    x"270BCEB",
    x"270BABC",
    x"270B88D",
    x"270B65F",
    x"270B432",
    x"270B205",
    x"270AFD9",
    x"270ADAD",
    x"270AB82",
    x"270A958",
    x"270A72D",
    x"270A504",
    x"270A2DB",
    x"270A0B2",
    x"2709E8B",
    x"2709C63",
    x"2709A3C",
    x"2709816",
    x"27095F0",
    x"27093CB",
    x"27091A6",
    x"2708F82",
    x"2708D5F",
    x"2708B3C",
    x"2708919",
    x"27086F7",
    x"27084D6",
    x"27082B5",
    x"2708094",
    x"2707E74",
    x"2707C55",
    x"2707A36",
    x"2707818",
    x"27075FA",
    x"27073DD",
    x"27071C0",
    x"2706FA4",
    x"2706D88",
    x"2706B6D",
    x"2706953",
    x"2706739",
    x"270651F",
    x"2706306",
    x"27060EE",
    x"2705ED6",
    x"2705CBE",
    x"2705AA7",
    x"2705891",
    x"270567B",
    x"2705466",
    x"2705251",
    x"270503C",
    x"2704E29",
    x"2704C15",
    x"2704A03",
    x"27047F0",
    x"27045DF",
    x"27043CD",
    x"27041BD",
    x"2703FAD",
    x"2703D9D",
    x"2703B8E",
    x"270397F",
    x"2703771",
    x"2703563",
    x"2703356",
    x"270314A",
    x"2702F3E",
    x"2702D32",
    x"2702B27",
    x"270291C",
    x"2702712",
    x"2702509",
    x"2702300",
    x"27020F7",
    x"2701EEF",
    x"2701CE8",
    x"2701AE1",
    x"27018DB",
    x"27016D5",
    x"27014CF",
    x"27012CA",
    x"27010C6",
    x"2700EC2",
    x"2700CBE",
    x"2700ABB",
    x"27008B9",
    x"27006B7",
    x"27004B6",
    x"27002B5",
    x"27000B4",
    x"26FFD69",
    x"26FF96A",
    x"26FF56C",
    x"26FF170",
    x"26FED74",
    x"26FE979",
    x"26FE57F",
    x"26FE186",
    x"26FDD8E",
    x"26FD997",
    x"26FD5A1",
    x"26FD1AD",
    x"26FCDB9",
    x"26FC9C6",
    x"26FC5D4",
    x"26FC1E3",
    x"26FBDF3",
    x"26FBA04",
    x"26FB616",
    x"26FB229",
    x"26FAE3D",
    x"26FAA52",
    x"26FA667",
    x"26FA27E",
    x"26F9E96",
    x"26F9AAF",
    x"26F96C9",
    x"26F92E4",
    x"26F8EFF",
    x"26F8B1C",
    x"26F873A",
    x"26F8359",
    x"26F7F78",
    x"26F7B99",
    x"26F77BA",
    x"26F73DD",
    x"26F7000",
    x"26F6C25",
    x"26F684A",
    x"26F6471",
    x"26F6098",
    x"26F5CC1",
    x"26F58EA",
    x"26F5514",
    x"26F513F",
    x"26F4D6B",
    x"26F4999",
    x"26F45C7",
    x"26F41F6",
    x"26F3E26",
    x"26F3A57",
    x"26F3689",
    x"26F32BB",
    x"26F2EEF",
    x"26F2B24",
    x"26F275A",
    x"26F2390",
    x"26F1FC8",
    x"26F1C00",
    x"26F183A",
    x"26F1474",
    x"26F10B0",
    x"26F0CEC",
    x"26F0929",
    x"26F0567",
    x"26F01A6",
    x"26EFDE6",
    x"26EFA27",
    x"26EF669",
    x"26EF2AC",
    x"26EEEF0",
    x"26EEB35",
    x"26EE77A",
    x"26EE3C1",
    x"26EE009",
    x"26EDC51",
    x"26ED89A",
    x"26ED4E5",
    x"26ED130",
    x"26ECD7C",
    x"26EC9C9",
    x"26EC617",
    x"26EC266",
    x"26EBEB6",
    x"26EBB07",
    x"26EB758",
    x"26EB3AB",
    x"26EAFFF",
    x"26EAC53",
    x"26EA8A8",
    x"26EA4FF",
    x"26EA156",
    x"26E9DAE",
    x"26E9A07",
    x"26E9661",
    x"26E92BC",
    x"26E8F18",
    x"26E8B74",
    x"26E87D2",
    x"26E8431",
    x"26E8090",
    x"26E7CF0",
    x"26E7951",
    x"26E75B4",
    x"26E7217",
    x"26E6E7B",
    x"26E6ADF",
    x"26E6745",
    x"26E63AC",
    x"26E6013",
    x"26E5C7C",
    x"26E58E5",
    x"26E554F",
    x"26E51BA",
    x"26E4E26",
    x"26E4A93",
    x"26E4701",
    x"26E4370",
    x"26E3FDF",
    x"26E3C50",
    x"26E38C1",
    x"26E3533",
    x"26E31A7",
    x"26E2E1B",
    x"26E2A90",
    x"26E2705",
    x"26E237C",
    x"26E1FF4",
    x"26E1C6C",
    x"26E18E5",
    x"26E1560",
    x"26E11DB",
    x"26E0E57",
    x"26E0AD4",
    x"26E0751",
    x"26E03D0",
    x"26E004F",
    x"26DFCD0",
    x"26DF951",
    x"26DF5D3",
    x"26DF256",
    x"26DEEDA",
    x"26DEB5F",
    x"26DE7E4",
    x"26DE46B",
    x"26DE0F2",
    x"26DDD7A",
    x"26DDA03",
    x"26DD68D",
    x"26DD318",
    x"26DCFA4",
    x"26DCC30",
    x"26DC8BE",
    x"26DC54C",
    x"26DC1DB",
    x"26DBE6B",
    x"26DBAFC",
    x"26DB78D",
    x"26DB420",
    x"26DB0B3",
    x"26DAD48",
    x"26DA9DD",
    x"26DA673",
    x"26DA309",
    x"26D9FA1",
    x"26D9C3A",
    x"26D98D3",
    x"26D956D",
    x"26D9208",
    x"26D8EA4",
    x"26D8B41",
    x"26D87DF",
    x"26D847D",
    x"26D811C",
    x"26D7DBC",
    x"26D7A5D",
    x"26D76FF",
    x"26D73A2",
    x"26D7045",
    x"26D6CEA",
    x"26D698F",
    x"26D6635",
    x"26D62DC",
    x"26D5F84",
    x"26D5C2C",
    x"26D58D6",
    x"26D5580",
    x"26D522B",
    x"26D4ED7",
    x"26D4B83",
    x"26D4831",
    x"26D44DF",
    x"26D418E",
    x"26D3E3E",
    x"26D3AEF",
    x"26D37A1",
    x"26D3453",
    x"26D3107",
    x"26D2DBB",
    x"26D2A70",
    x"26D2726",
    x"26D23DC",
    x"26D2094",
    x"26D1D4C",
    x"26D1A05",
    x"26D16BF",
    x"26D137A",
    x"26D1035",
    x"26D0CF2",
    x"26D09AF",
    x"26D066D",
    x"26D032C",
    x"26CFFEB",
    x"26CFCAC",
    x"26CF96D",
    x"26CF62F",
    x"26CF2F2",
    x"26CEFB6",
    x"26CEC7A",
    x"26CE93F",
    x"26CE605",
    x"26CE2CC",
    x"26CDF94",
    x"26CDC5C",
    x"26CD926",
    x"26CD5F0",
    x"26CD2BB",
    x"26CCF87",
    x"26CCC53",
    x"26CC920",
    x"26CC5EE",
    x"26CC2BD",
    x"26CBF8D",
    x"26CBC5E",
    x"26CB92F",
    x"26CB601",
    x"26CB2D4",
    x"26CAFA8",
    x"26CAC7C",
    x"26CA951",
    x"26CA627",
    x"26CA2FE",
    x"26C9FD6",
    x"26C9CAE",
    x"26C9988",
    x"26C9662",
    x"26C933C",
    x"26C9018",
    x"26C8CF4",
    x"26C89D2",
    x"26C86AF",
    x"26C838E",
    x"26C806E",
    x"26C7D4E",
    x"26C7A2F",
    x"26C7711",
    x"26C73F3",
    x"26C70D7",
    x"26C6DBB",
    x"26C6AA0",
    x"26C6786",
    x"26C646C",
    x"26C6154",
    x"26C5E3C",
    x"26C5B24",
    x"26C580E",
    x"26C54F8",
    x"26C51E4",
    x"26C4ECF",
    x"26C4BBC",
    x"26C48AA",
    x"26C4598",
    x"26C4287",
    x"26C3F77",
    x"26C3C67",
    x"26C3958",
    x"26C364A",
    x"26C333D",
    x"26C3031",
    x"26C2D25",
    x"26C2A1A",
    x"26C2710",
    x"26C2407",
    x"26C20FE",
    x"26C1DF6",
    x"26C1AEF",
    x"26C17E9",
    x"26C14E3",
    x"26C11DE",
    x"26C0EDA",
    x"26C0BD7",
    x"26C08D4",
    x"26C05D2",
    x"26C02D1",
    x"26BFFD1",
    x"26BFCD1",
    x"26BF9D3",
    x"26BF6D4",
    x"26BF3D7",
    x"26BF0DB",
    x"26BEDDF",
    x"26BEAE4",
    x"26BE7E9",
    x"26BE4F0",
    x"26BE1F7",
    x"26BDEFF",
    x"26BDC07",
    x"26BD911",
    x"26BD61B",
    x"26BD326",
    x"26BD031",
    x"26BCD3E",
    x"26BCA4B",
    x"26BC758",
    x"26BC467",
    x"26BC176",
    x"26BBE86",
    x"26BBB97",
    x"26BB8A8",
    x"26BB5BB",
    x"26BB2CE",
    x"26BAFE1",
    x"26BACF6",
    x"26BAA0B",
    x"26BA721",
    x"26BA437",
    x"26BA14E",
    x"26B9E66",
    x"26B9B7F",
    x"26B9899",
    x"26B95B3",
    x"26B92CE",
    x"26B8FEA",
    x"26B8D06",
    x"26B8A23",
    x"26B8741",
    x"26B845F",
    x"26B817F",
    x"26B7E9F",
    x"26B7BBF",
    x"26B78E1",
    x"26B7603",
    x"26B7326",
    x"26B7049",
    x"26B6D6E",
    x"26B6A93",
    x"26B67B8",
    x"26B64DF",
    x"26B6206",
    x"26B5F2E",
    x"26B5C56",
    x"26B5980",
    x"26B56AA",
    x"26B53D4",
    x"26B5100",
    x"26B4E2C",
    x"26B4B59",
    x"26B4886",
    x"26B45B4",
    x"26B42E3",
    x"26B4013",
    x"26B3D43",
    x"26B3A74",
    x"26B37A6",
    x"26B34D8",
    x"26B320C",
    x"26B2F3F",
    x"26B2C74",
    x"26B29A9",
    x"26B26DF",
    x"26B2416",
    x"26B214D",
    x"26B1E85",
    x"26B1BBE",
    x"26B18F7",
    x"26B1631",
    x"26B136C",
    x"26B10A8",
    x"26B0DE4",
    x"26B0B21",
    x"26B085E",
    x"26B059C",
    x"26B02DB",
    x"26B001B",
    x"26AFD5B",
    x"26AFA9C",
    x"26AF7DE",
    x"26AF520",
    x"26AF263",
    x"26AEFA7",
    x"26AECEC",
    x"26AEA31",
    x"26AE777",
    x"26AE4BD",
    x"26AE204",
    x"26ADF4C",
    x"26ADC95",
    x"26AD9DE",
    x"26AD728",
    x"26AD472",
    x"26AD1BD",
    x"26ACF09",
    x"26ACC56",
    x"26AC9A3",
    x"26AC6F1",
    x"26AC440",
    x"26AC18F",
    x"26ABEDF",
    x"26ABC2F",
    x"26AB981",
    x"26AB6D3",
    x"26AB425",
    x"26AB179",
    x"26AAECD",
    x"26AAC21",
    x"26AA977",
    x"26AA6CC",
    x"26AA423",
    x"26AA17A",
    x"26A9ED2",
    x"26A9C2B",
    x"26A9984",
    x"26A96DE",
    x"26A9439",
    x"26A9194",
    x"26A8EF0",
    x"26A8C4D",
    x"26A89AA",
    x"26A8708",
    x"26A8466",
    x"26A81C6",
    x"26A7F26",
    x"26A7C86",
    x"26A79E7",
    x"26A7749",
    x"26A74AC",
    x"26A720F",
    x"26A6F73",
    x"26A6CD7",
    x"26A6A3C",
    x"26A67A2",
    x"26A6508",
    x"26A626F",
    x"26A5FD7",
    x"26A5D3F",
    x"26A5AA8",
    x"26A5812",
    x"26A557C",
    x"26A52E7",
    x"26A5053",
    x"26A4DBF",
    x"26A4B2C",
    x"26A489A",
    x"26A4608",
    x"26A4377",
    x"26A40E6",
    x"26A3E56",
    x"26A3BC7",
    x"26A3938",
    x"26A36AA",
    x"26A341D",
    x"26A3190",
    x"26A2F04",
    x"26A2C79",
    x"26A29EE",
    x"26A2764",
    x"26A24DA",
    x"26A2251",
    x"26A1FC9",
    x"26A1D41",
    x"26A1ABA",
    x"26A1834",
    x"26A15AE",
    x"26A1329",
    x"26A10A5",
    x"26A0E21",
    x"26A0B9E",
    x"26A091B",
    x"26A0699",
    x"26A0418",
    x"26A0197",
    x"269FF17",
    x"269FC98",
    x"269FA19",
    x"269F79B",
    x"269F51D",
    x"269F2A0",
    x"269F024",
    x"269EDA8",
    x"269EB2D",
    x"269E8B2",
    x"269E638",
    x"269E3BF",
    x"269E147",
    x"269DECF",
    x"269DC57",
    x"269D9E0",
    x"269D76A",
    x"269D4F5",
    x"269D280",
    x"269D00B",
    x"269CD98",
    x"269CB25",
    x"269C8B2",
    x"269C640",
    x"269C3CF",
    x"269C15E",
    x"269BEEE",
    x"269BC7F",
    x"269BA10",
    x"269B7A2",
    x"269B534",
    x"269B2C7",
    x"269B05B",
    x"269ADEF",
    x"269AB84",
    x"269A919",
    x"269A6AF",
    x"269A446",
    x"269A1DD",
    x"2699F75",
    x"2699D0D",
    x"2699AA7",
    x"2699840",
    x"26995DA",
    x"2699375",
    x"2699111",
    x"2698EAD",
    x"2698C49",
    x"26989E7",
    x"2698784",
    x"2698523",
    x"26982C2",
    x"2698061",
    x"2697E02",
    x"2697BA2",
    x"2697944",
    x"26976E6",
    x"2697488",
    x"269722C",
    x"2696FCF",
    x"2696D74",
    x"2696B19",
    x"26968BE",
    x"2696664",
    x"269640B",
    x"26961B2",
    x"2695F5A",
    x"2695D02",
    x"2695AAC",
    x"2695855",
    x"26955FF",
    x"26953AA",
    x"2695156",
    x"2694F01",
    x"2694CAE",
    x"2694A5B",
    x"2694809",
    x"26945B7",
    x"2694366",
    x"2694115",
    x"2693EC5",
    x"2693C76",
    x"2693A27",
    x"26937D9",
    x"269358B",
    x"269333E",
    x"26930F2",
    x"2692EA6",
    x"2692C5A",
    x"2692A10",
    x"26927C5",
    x"269257C",
    x"2692333",
    x"26920EA",
    x"2691EA2",
    x"2691C5B",
    x"2691A14",
    x"26917CE",
    x"2691588",
    x"2691343",
    x"26910FE",
    x"2690EBA",
    x"2690C77",
    x"2690A34",
    x"26907F2",
    x"26905B0",
    x"269036F",
    x"269012E",
    x"268FEEE",
    x"268FCAF",
    x"268FA70",
    x"268F832",
    x"268F5F4",
    x"268F3B7",
    x"268F17A",
    x"268EF3E",
    x"268ED03",
    x"268EAC8",
    x"268E88D",
    x"268E653",
    x"268E41A",
    x"268E1E1",
    x"268DFA9",
    x"268DD71",
    x"268DB3A",
    x"268D904",
    x"268D6CE",
    x"268D498",
    x"268D264",
    x"268D02F",
    x"268CDFB",
    x"268CBC8",
    x"268C996",
    x"268C763",
    x"268C532",
    x"268C301",
    x"268C0D0",
    x"268BEA0",
    x"268BC71",
    x"268BA42",
    x"268B814",
    x"268B5E6",
    x"268B3B9",
    x"268B18C",
    x"268AF60",
    x"268AD35",
    x"268AB0A",
    x"268A8DF",
    x"268A6B5",
    x"268A48C",
    x"268A263",
    x"268A03B",
    x"2689E13",
    x"2689BEB",
    x"26899C5",
    x"268979F",
    x"2689579",
    x"2689354",
    x"268912F",
    x"2688F0B",
    x"2688CE8",
    x"2688AC5",
    x"26888A2",
    x"2688680",
    x"268845F",
    x"268823E",
    x"268801E",
    x"2687DFE",
    x"2687BDF",
    x"26879C0",
    x"26877A2",
    x"2687584",
    x"2687367",
    x"268714B",
    x"2686F2F",
    x"2686D13",
    x"2686AF8",
    x"26868DE",
    x"26866C4",
    x"26864AA",
    x"2686291",
    x"2686079",
    x"2685E61",
    x"2685C4A",
    x"2685A33",
    x"268581D",
    x"2685607",
    x"26853F2",
    x"26851DD",
    x"2684FC9",
    x"2684DB5",
    x"2684BA2",
    x"268498F",
    x"268477D",
    x"268456C",
    x"268435A",
    x"268414A",
    x"2683F3A",
    x"2683D2A",
    x"2683B1B",
    x"268390D",
    x"26836FF",
    x"26834F1",
    x"26832E4",
    x"26830D8",
    x"2682ECC",
    x"2682CC0",
    x"2682AB5",
    x"26828AB",
    x"26826A1",
    x"2682498",
    x"268228F",
    x"2682086",
    x"2681E7F",
    x"2681C77",
    x"2681A70",
    x"268186A",
    x"2681664",
    x"268145F",
    x"268125A",
    x"2681056",
    x"2680E52",
    x"2680C4E",
    x"2680A4C",
    x"2680849",
    x"2680647",
    x"2680446",
    x"2680245",
    x"2680045",
    x"267FC8B",
    x"267F88C",
    x"267F48F",
    x"267F092",
    x"267EC96",
    x"267E89C",
    x"267E4A2",
    x"267E0A9",
    x"267DCB2",
    x"267D8BB",
    x"267D4C5",
    x"267D0D1",
    x"267CCDD",
    x"267C8EA",
    x"267C4F8",
    x"267C108",
    x"267BD18",
    x"267B929",
    x"267B53B",
    x"267B14E",
    x"267AD63",
    x"267A978",
    x"267A58E",
    x"267A1A5",
    x"2679DBD",
    x"26799D6",
    x"26795F0",
    x"267920B",
    x"2678E27",
    x"2678A44",
    x"2678662",
    x"2678281",
    x"2677EA1",
    x"2677AC2",
    x"26776E3",
    x"2677306",
    x"2676F2A",
    x"2676B4F",
    x"2676774",
    x"267639B",
    x"2675FC2",
    x"2675BEB",
    x"2675814",
    x"267543F",
    x"267506A",
    x"2674C97",
    x"26748C4",
    x"26744F2",
    x"2674122",
    x"2673D52",
    x"2673983",
    x"26735B5",
    x"26731E8",
    x"2672E1C",
    x"2672A51",
    x"2672687",
    x"26722BE",
    x"2671EF5",
    x"2671B2E",
    x"2671768",
    x"26713A3",
    x"2670FDE",
    x"2670C1B",
    x"2670858",
    x"2670496",
    x"26700D6",
    x"266FD16",
    x"266F957",
    x"266F599",
    x"266F1DC",
    x"266EE20",
    x"266EA65",
    x"266E6AB",
    x"266E2F2",
    x"266DF3A",
    x"266DB82",
    x"266D7CC",
    x"266D416",
    x"266D062",
    x"266CCAE",
    x"266C8FC",
    x"266C54A",
    x"266C199",
    x"266BDE9",
    x"266BA3A",
    x"266B68C",
    x"266B2DF",
    x"266AF32",
    x"266AB87",
    x"266A7DD",
    x"266A433",
    x"266A08B",
    x"2669CE3",
    x"266993C",
    x"2669596",
    x"26691F1",
    x"2668E4D",
    x"2668AAA",
    x"2668708",
    x"2668367",
    x"2667FC6",
    x"2667C27",
    x"2667888",
    x"26674EA",
    x"266714E",
    x"2666DB2",
    x"2666A17",
    x"266667D",
    x"26662E4",
    x"2665F4B",
    x"2665BB4",
    x"266581E",
    x"2665488",
    x"26650F3",
    x"2664D5F",
    x"26649CD",
    x"266463B",
    x"26642A9",
    x"2663F19",
    x"2663B8A",
    x"26637FB",
    x"266346E",
    x"26630E1",
    x"2662D55",
    x"26629CB",
    x"2662641",
    x"26622B7",
    x"2661F2F",
    x"2661BA8",
    x"2661821",
    x"266149C",
    x"2661117",
    x"2660D93",
    x"2660A10",
    x"266068E",
    x"266030D",
    x"265FF8D",
    x"265FC0D",
    x"265F88F",
    x"265F511",
    x"265F194",
    x"265EE18",
    x"265EA9D",
    x"265E723",
    x"265E3A9",
    x"265E031",
    x"265DCB9",
    x"265D943",
    x"265D5CD",
    x"265D258",
    x"265CEE4",
    x"265CB70",
    x"265C7FE",
    x"265C48C",
    x"265C11C",
    x"265BDAC",
    x"265BA3D",
    x"265B6CF",
    x"265B361",
    x"265AFF5",
    x"265AC89",
    x"265A91F",
    x"265A5B5",
    x"265A24C",
    x"2659EE4",
    x"2659B7C",
    x"2659816",
    x"26594B0",
    x"265914C",
    x"2658DE8",
    x"2658A85",
    x"2658722",
    x"26583C1",
    x"2658061",
    x"2657D01",
    x"26579A2",
    x"2657644",
    x"26572E7",
    x"2656F8B",
    x"2656C2F",
    x"26568D4",
    x"265657B",
    x"2656222",
    x"2655ECA",
    x"2655B72",
    x"265581C",
    x"26554C6",
    x"2655172",
    x"2654E1E",
    x"2654ACA",
    x"2654778",
    x"2654427",
    x"26540D6",
    x"2653D86",
    x"2653A37",
    x"26536E9",
    x"265339C",
    x"265304F",
    x"2652D04",
    x"26529B9",
    x"265266F",
    x"2652326",
    x"2651FDD",
    x"2651C96",
    x"265194F",
    x"2651609",
    x"26512C4",
    x"2650F80",
    x"2650C3C",
    x"26508FA",
    x"26505B8",
    x"2650277",
    x"264FF37",
    x"264FBF7",
    x"264F8B9",
    x"264F57B",
    x"264F23E",
    x"264EF02",
    x"264EBC6",
    x"264E88C",
    x"264E552",
    x"264E219",
    x"264DEE1",
    x"264DBAA",
    x"264D873",
    x"264D53D",
    x"264D208",
    x"264CED4",
    x"264CBA1",
    x"264C86F",
    x"264C53D",
    x"264C20C",
    x"264BEDC",
    x"264BBAD",
    x"264B87E",
    x"264B550",
    x"264B223",
    x"264AEF7",
    x"264ABCC",
    x"264A8A1",
    x"264A578",
    x"264A24F",
    x"2649F26",
    x"2649BFF",
    x"26498D8",
    x"26495B3",
    x"264928E",
    x"2648F69",
    x"2648C46",
    x"2648923",
    x"2648601",
    x"26482E0",
    x"2647FC0",
    x"2647CA0",
    x"2647982",
    x"2647664",
    x"2647346",
    x"264702A",
    x"2646D0E",
    x"26469F3",
    x"26466D9",
    x"26463C0",
    x"26460A7",
    x"2645D90",
    x"2645A79",
    x"2645762",
    x"264544D",
    x"2645138",
    x"2644E24",
    x"2644B11",
    x"26447FF",
    x"26444ED",
    x"26441DC",
    x"2643ECC",
    x"2643BBD",
    x"26438AE",
    x"26435A1",
    x"2643294",
    x"2642F87",
    x"2642C7C",
    x"2642971",
    x"2642667",
    x"264235E",
    x"2642055",
    x"2641D4E",
    x"2641A47",
    x"2641741",
    x"264143B",
    x"2641136",
    x"2640E32",
    x"2640B2F",
    x"264082D",
    x"264052B",
    x"264022A",
    x"263FF2A",
    x"263FC2B",
    x"263F92C",
    x"263F62E",
    x"263F331",
    x"263F035",
    x"263ED39",
    x"263EA3E",
    x"263E744",
    x"263E44A",
    x"263E152",
    x"263DE5A",
    x"263DB62",
    x"263D86C",
    x"263D576",
    x"263D281",
    x"263CF8D",
    x"263CC99",
    x"263C9A7",
    x"263C6B5",
    x"263C3C3",
    x"263C0D3",
    x"263BDE3",
    x"263BAF4",
    x"263B805",
    x"263B518",
    x"263B22B",
    x"263AF3F",
    x"263AC53",
    x"263A969",
    x"263A67F",
    x"263A395",
    x"263A0AD",
    x"2639DC5",
    x"2639ADE",
    x"26397F7",
    x"2639512",
    x"263922D",
    x"2638F49",
    x"2638C65",
    x"2638983",
    x"26386A1",
    x"26383BF",
    x"26380DF",
    x"2637DFF",
    x"2637B20",
    x"2637841",
    x"2637564",
    x"2637287",
    x"2636FAA",
    x"2636CCF",
    x"26369F4",
    x"263671A",
    x"2636440",
    x"2636168",
    x"2635E90",
    x"2635BB8",
    x"26358E2",
    x"263560C",
    x"2635337",
    x"2635062",
    x"2634D8F",
    x"2634ABC",
    x"26347E9",
    x"2634518",
    x"2634247",
    x"2633F76",
    x"2633CA7",
    x"26339D8",
    x"263370A",
    x"263343D",
    x"2633170",
    x"2632EA4",
    x"2632BD9",
    x"263290E",
    x"2632644",
    x"263237B",
    x"26320B2",
    x"2631DEA",
    x"2631B23",
    x"263185D",
    x"2631597",
    x"26312D2",
    x"263100E",
    x"2630D4A",
    x"2630A87",
    x"26307C5",
    x"2630503",
    x"2630242",
    x"262FF82",
    x"262FCC3",
    x"262FA04",
    x"262F746",
    x"262F488",
    x"262F1CB",
    x"262EF0F",
    x"262EC54",
    x"262E999",
    x"262E6DF",
    x"262E426",
    x"262E16D",
    x"262DEB5",
    x"262DBFD",
    x"262D947",
    x"262D691",
    x"262D3DC",
    x"262D127",
    x"262CE73",
    x"262CBC0",
    x"262C90D",
    x"262C65B",
    x"262C3AA",
    x"262C0F9",
    x"262BE49",
    x"262BB9A",
    x"262B8EC",
    x"262B63E",
    x"262B390",
    x"262B0E4",
    x"262AE38",
    x"262AB8D",
    x"262A8E2",
    x"262A638",
    x"262A38F",
    x"262A0E7",
    x"2629E3F",
    x"2629B97",
    x"26298F1",
    x"262964B",
    x"26293A6",
    x"2629101",
    x"2628E5D",
    x"2628BBA",
    x"2628917",
    x"2628675",
    x"26283D4",
    x"2628134",
    x"2627E94",
    x"2627BF4",
    x"2627956",
    x"26276B8",
    x"262741A",
    x"262717E",
    x"2626EE1",
    x"2626C46",
    x"26269AB",
    x"2626711",
    x"2626478",
    x"26261DF",
    x"2625F47",
    x"2625CAF",
    x"2625A19",
    x"2625782",
    x"26254ED",
    x"2625258",
    x"2624FC4",
    x"2624D30",
    x"2624A9D",
    x"262480B",
    x"2624579",
    x"26242E8",
    x"2624058",
    x"2623DC8",
    x"2623B39",
    x"26238AA",
    x"262361C",
    x"262338F",
    x"2623103",
    x"2622E77",
    x"2622BEB",
    x"2622961",
    x"26226D7",
    x"262244D",
    x"26221C4",
    x"2621F3C",
    x"2621CB5",
    x"2621A2E",
    x"26217A8",
    x"2621522",
    x"262129D",
    x"2621019",
    x"2620D95",
    x"2620B12",
    x"2620890",
    x"262060E",
    x"262038D",
    x"262010C",
    x"261FE8C",
    x"261FC0D",
    x"261F98E",
    x"261F710",
    x"261F492",
    x"261F216",
    x"261EF99",
    x"261ED1E",
    x"261EAA3",
    x"261E829",
    x"261E5AF",
    x"261E336",
    x"261E0BD",
    x"261DE45",
    x"261DBCE",
    x"261D957",
    x"261D6E1",
    x"261D46C",
    x"261D1F7",
    x"261CF83",
    x"261CD0F",
    x"261CA9C",
    x"261C82A",
    x"261C5B8",
    x"261C347",
    x"261C0D7",
    x"261BE67",
    x"261BBF8",
    x"261B989",
    x"261B71B",
    x"261B4AD",
    x"261B240",
    x"261AFD4",
    x"261AD68",
    x"261AAFD",
    x"261A893",
    x"261A629",
    x"261A3C0",
    x"261A157",
    x"2619EEF",
    x"2619C88",
    x"2619A21",
    x"26197BB",
    x"2619555",
    x"26192F0",
    x"261908C",
    x"2618E28",
    x"2618BC5",
    x"2618962",
    x"2618700",
    x"261849E",
    x"261823E",
    x"2617FDD",
    x"2617D7E",
    x"2617B1F",
    x"26178C0",
    x"2617662",
    x"2617405",
    x"26171A8",
    x"2616F4C",
    x"2616CF1",
    x"2616A96",
    x"261683B",
    x"26165E1",
    x"2616388",
    x"2616130",
    x"2615ED8",
    x"2615C80",
    x"2615A29",
    x"26157D3",
    x"261557E",
    x"2615328",
    x"26150D4",
    x"2614E80",
    x"2614C2D",
    x"26149DA",
    x"2614788",
    x"2614536",
    x"26142E5",
    x"2614095",
    x"2613E45",
    x"2613BF6",
    x"26139A7",
    x"2613759",
    x"261350B",
    x"26132BE",
    x"2613072",
    x"2612E26",
    x"2612BDB",
    x"2612990",
    x"2612746",
    x"26124FC",
    x"26122B3",
    x"261206B",
    x"2611E23",
    x"2611BDC",
    x"2611995",
    x"261174F",
    x"261150A",
    x"26112C5",
    x"2611080",
    x"2610E3C",
    x"2610BF9",
    x"26109B6",
    x"2610774",
    x"2610533",
    x"26102F2",
    x"26100B1",
    x"260FE71",
    x"260FC32",
    x"260F9F3",
    x"260F7B5",
    x"260F577",
    x"260F33A",
    x"260F0FE",
    x"260EEC2",
    x"260EC86",
    x"260EA4C",
    x"260E811",
    x"260E5D8",
    x"260E39E",
    x"260E166",
    x"260DF2E",
    x"260DCF6",
    x"260DABF",
    x"260D889",
    x"260D653",
    x"260D41E",
    x"260D1E9",
    x"260CFB5",
    x"260CD81",
    x"260CB4E",
    x"260C91B",
    x"260C6E9",
    x"260C4B8",
    x"260C287",
    x"260C057",
    x"260BE27",
    x"260BBF8",
    x"260B9C9",
    x"260B79B",
    x"260B56D",
    x"260B340",
    x"260B113",
    x"260AEE7",
    x"260ACBC",
    x"260AA91",
    x"260A867",
    x"260A63D",
    x"260A414",
    x"260A1EB",
    x"2609FC3",
    x"2609D9B",
    x"2609B74",
    x"260994D",
    x"2609727",
    x"2609502",
    x"26092DD",
    x"26090B8",
    x"2608E94",
    x"2608C71",
    x"2608A4E",
    x"260882C",
    x"260860A",
    x"26083E9",
    x"26081C8",
    x"2607FA8",
    x"2607D88",
    x"2607B69",
    x"260794A",
    x"260772C",
    x"260750F",
    x"26072F2",
    x"26070D5",
    x"2606EB9",
    x"2606C9E",
    x"2606A83",
    x"2606869",
    x"260664F",
    x"2606436",
    x"260621D",
    x"2606005",
    x"2605DED",
    x"2605BD6",
    x"26059BF",
    x"26057A9",
    x"2605593",
    x"260537E",
    x"2605169",
    x"2604F55",
    x"2604D42",
    x"2604B2F",
    x"260491C",
    x"260470A",
    x"26044F9",
    x"26042E8",
    x"26040D7",
    x"2603EC7",
    x"2603CB8",
    x"2603AA9",
    x"260389A",
    x"260368C",
    x"260347F",
    x"2603272",
    x"2603066",
    x"2602E5A",
    x"2602C4F",
    x"2602A44",
    x"260283A",
    x"2602630",
    x"2602426",
    x"260221E",
    x"2602015",
    x"2601E0E",
    x"2601C06",
    x"2601A00",
    x"26017F9",
    x"26015F4",
    x"26013EE",
    x"26011EA",
    x"2600FE5",
    x"2600DE2",
    x"2600BDF",
    x"26009DC",
    x"26007DA",
    x"26005D8",
    x"26003D7",
    x"26001D6",
    x"25FFFAC",
    x"25FFBAD",
    x"25FF7AE",
    x"25FF3B1",
    x"25FEFB4",
    x"25FEBB9",
    x"25FE7BE",
    x"25FE3C5",
    x"25FDFCD",
    x"25FDBD5",
    x"25FD7DF",
    x"25FD3E9",
    x"25FCFF5",
    x"25FCC01",
    x"25FC80F",
    x"25FC41D",
    x"25FC02D",
    x"25FBC3D",
    x"25FB84E",
    x"25FB461",
    x"25FB074",
    x"25FAC89",
    x"25FA89E",
    x"25FA4B4",
    x"25FA0CC",
    x"25F9CE4",
    x"25F98FD",
    x"25F9517",
    x"25F9133",
    x"25F8D4F",
    x"25F896C",
    x"25F858A",
    x"25F81A9",
    x"25F7DC9",
    x"25F79EA",
    x"25F760C",
    x"25F722F",
    x"25F6E53",
    x"25F6A78",
    x"25F669E",
    x"25F62C5",
    x"25F5EED",
    x"25F5B15",
    x"25F573F",
    x"25F536A",
    x"25F4F95",
    x"25F4BC2",
    x"25F47EF",
    x"25F441E",
    x"25F404D",
    x"25F3C7E",
    x"25F38AF",
    x"25F34E1",
    x"25F3115",
    x"25F2D49",
    x"25F297E",
    x"25F25B4",
    x"25F21EB",
    x"25F1E23",
    x"25F1A5C",
    x"25F1696",
    x"25F12D1",
    x"25F0F0D",
    x"25F0B49",
    x"25F0787",
    x"25F03C6",
    x"25F0005",
    x"25EFC46",
    x"25EF887",
    x"25EF4C9",
    x"25EF10D",
    x"25EED51",
    x"25EE996",
    x"25EE5DC",
    x"25EE223",
    x"25EDE6B",
    x"25EDAB4",
    x"25ED6FE",
    x"25ED348",
    x"25ECF94",
    x"25ECBE0",
    x"25EC82E",
    x"25EC47C",
    x"25EC0CC",
    x"25EBD1C",
    x"25EB96D",
    x"25EB5BF",
    x"25EB212",
    x"25EAE66",
    x"25EAABB",
    x"25EA711",
    x"25EA368",
    x"25E9FBF",
    x"25E9C18",
    x"25E9871",
    x"25E94CB",
    x"25E9127",
    x"25E8D83",
    x"25E89E0",
    x"25E863E",
    x"25E829D",
    x"25E7EFD",
    x"25E7B5D",
    x"25E77BF",
    x"25E7421",
    x"25E7085",
    x"25E6CE9",
    x"25E694E",
    x"25E65B5",
    x"25E621C",
    x"25E5E84",
    x"25E5AEC",
    x"25E5756",
    x"25E53C1",
    x"25E502C",
    x"25E4C99",
    x"25E4906",
    x"25E4574",
    x"25E41E3",
    x"25E3E53",
    x"25E3AC4",
    x"25E3736",
    x"25E33A8",
    x"25E301C",
    x"25E2C90",
    x"25E2906",
    x"25E257C",
    x"25E21F3",
    x"25E1E6B",
    x"25E1AE4",
    x"25E175D",
    x"25E13D8",
    x"25E1053",
    x"25E0CD0",
    x"25E094D",
    x"25E05CB",
    x"25E024A",
    x"25DFECA",
    x"25DFB4B",
    x"25DF7CC",
    x"25DF44F",
    x"25DF0D2",
    x"25DED56",
    x"25DE9DC",
    x"25DE662",
    x"25DE2E8",
    x"25DDF70",
    x"25DDBF9",
    x"25DD882",
    x"25DD50C",
    x"25DD198",
    x"25DCE24",
    x"25DCAB0",
    x"25DC73E",
    x"25DC3CD",
    x"25DC05C",
    x"25DBCED",
    x"25DB97E",
    x"25DB610",
    x"25DB2A3",
    x"25DAF37",
    x"25DABCB",
    x"25DA861",
    x"25DA4F7",
    x"25DA18E",
    x"25D9E26",
    x"25D9ABF",
    x"25D9759",
    x"25D93F3",
    x"25D908F",
    x"25D8D2B",
    x"25D89C8",
    x"25D8666",
    x"25D8305",
    x"25D7FA5",
    x"25D7C45",
    x"25D78E7",
    x"25D7589",
    x"25D722C",
    x"25D6ED0",
    x"25D6B74",
    x"25D681A",
    x"25D64C0",
    x"25D6168",
    x"25D5E10",
    x"25D5AB9",
    x"25D5762",
    x"25D540D",
    x"25D50B8",
    x"25D4D65",
    x"25D4A12",
    x"25D46C0",
    x"25D436E",
    x"25D401E",
    x"25D3CCE",
    x"25D397F",
    x"25D3631",
    x"25D32E4",
    x"25D2F98",
    x"25D2C4D",
    x"25D2902",
    x"25D25B8",
    x"25D226F",
    x"25D1F27",
    x"25D1BDF",
    x"25D1899",
    x"25D1553",
    x"25D120E",
    x"25D0ECA",
    x"25D0B87",
    x"25D0844",
    x"25D0503",
    x"25D01C2",
    x"25CFE82",
    x"25CFB43",
    x"25CF804",
    x"25CF4C7",
    x"25CF18A",
    x"25CEE4E",
    x"25CEB13",
    x"25CE7D8",
    x"25CE49F",
    x"25CE166",
    x"25CDE2E",
    x"25CDAF7",
    x"25CD7C1",
    x"25CD48B",
    x"25CD156",
    x"25CCE22",
    x"25CCAEF",
    x"25CC7BD",
    x"25CC48B",
    x"25CC15B",
    x"25CBE2B",
    x"25CBAFB",
    x"25CB7CD",
    x"25CB4A0",
    x"25CB173",
    x"25CAE47",
    x"25CAB1C",
    x"25CA7F1",
    x"25CA4C8",
    x"25CA19F",
    x"25C9E77",
    x"25C9B50",
    x"25C9829",
    x"25C9504",
    x"25C91DF",
    x"25C8EBB",
    x"25C8B97",
    x"25C8875",
    x"25C8553",
    x"25C8232",
    x"25C7F12",
    x"25C7BF3",
    x"25C78D4",
    x"25C75B6",
    x"25C7299",
    x"25C6F7D",
    x"25C6C61",
    x"25C6947",
    x"25C662D",
    x"25C6314",
    x"25C5FFB",
    x"25C5CE4",
    x"25C59CD",
    x"25C56B7",
    x"25C53A1",
    x"25C508D",
    x"25C4D79",
    x"25C4A66",
    x"25C4754",
    x"25C4443",
    x"25C4132",
    x"25C3E22",
    x"25C3B13",
    x"25C3804",
    x"25C34F7",
    x"25C31EA",
    x"25C2EDE",
    x"25C2BD2",
    x"25C28C8",
    x"25C25BE",
    x"25C22B5",
    x"25C1FAD",
    x"25C1CA5",
    x"25C199E",
    x"25C1698",
    x"25C1393",
    x"25C108F",
    x"25C0D8B",
    x"25C0A88",
    x"25C0786",
    x"25C0484",
    x"25C0183",
    x"25BFE83",
    x"25BFB84",
    x"25BF886",
    x"25BF588",
    x"25BF28B",
    x"25BEF8F",
    x"25BEC93",
    x"25BE998",
    x"25BE69E",
    x"25BE3A5",
    x"25BE0AC",
    x"25BDDB5",
    x"25BDABE",
    x"25BD7C7",
    x"25BD4D2",
    x"25BD1DD",
    x"25BCEE9",
    x"25BCBF5",
    x"25BC903",
    x"25BC611",
    x"25BC320",
    x"25BC02F",
    x"25BBD40",
    x"25BBA51",
    x"25BB762",
    x"25BB475",
    x"25BB188",
    x"25BAE9C",
    x"25BABB1",
    x"25BA8C6",
    x"25BA5DD",
    x"25BA2F3",
    x"25BA00B",
    x"25B9D23",
    x"25B9A3C",
    x"25B9756",
    x"25B9471",
    x"25B918C",
    x"25B8EA8",
    x"25B8BC5",
    x"25B88E2",
    x"25B8600",
    x"25B831F",
    x"25B803F",
    x"25B7D5F",
    x"25B7A80",
    x"25B77A2",
    x"25B74C4",
    x"25B71E7",
    x"25B6F0B",
    x"25B6C30",
    x"25B6955",
    x"25B667B",
    x"25B63A2",
    x"25B60C9",
    x"25B5DF2",
    x"25B5B1A",
    x"25B5844",
    x"25B556E",
    x"25B5299",
    x"25B4FC5",
    x"25B4CF1",
    x"25B4A1E",
    x"25B474C",
    x"25B447B",
    x"25B41AA",
    x"25B3EDA",
    x"25B3C0B",
    x"25B393C",
    x"25B366E",
    x"25B33A1",
    x"25B30D4",
    x"25B2E08",
    x"25B2B3D",
    x"25B2873",
    x"25B25A9",
    x"25B22E0",
    x"25B2018",
    x"25B1D50",
    x"25B1A89",
    x"25B17C3",
    x"25B14FD",
    x"25B1238",
    x"25B0F74",
    x"25B0CB0",
    x"25B09EE",
    x"25B072B",
    x"25B046A",
    x"25B01A9",
    x"25AFEE9",
    x"25AFC2A",
    x"25AF96B",
    x"25AF6AD",
    x"25AF3F0",
    x"25AF133",
    x"25AEE77",
    x"25AEBBC",
    x"25AE901",
    x"25AE647",
    x"25AE38E",
    x"25AE0D6",
    x"25ADE1E",
    x"25ADB66",
    x"25AD8B0",
    x"25AD5FA",
    x"25AD345",
    x"25AD090",
    x"25ACDDD",
    x"25ACB2A",
    x"25AC877",
    x"25AC5C5",
    x"25AC314",
    x"25AC064",
    x"25ABDB4",
    x"25ABB05",
    x"25AB857",
    x"25AB5A9",
    x"25AB2FC",
    x"25AB04F",
    x"25AADA4",
    x"25AAAF8",
    x"25AA84E",
    x"25AA5A4",
    x"25AA2FB",
    x"25AA053",
    x"25A9DAB",
    x"25A9B04",
    x"25A985E",
    x"25A95B8",
    x"25A9313",
    x"25A906E",
    x"25A8DCA",
    x"25A8B27",
    x"25A8885",
    x"25A85E3",
    x"25A8342",
    x"25A80A1",
    x"25A7E02",
    x"25A7B62",
    x"25A78C4",
    x"25A7626",
    x"25A7389",
    x"25A70EC",
    x"25A6E50",
    x"25A6BB5",
    x"25A691B",
    x"25A6681",
    x"25A63E7",
    x"25A614F",
    x"25A5EB7",
    x"25A5C1F",
    x"25A5989",
    x"25A56F3",
    x"25A545D",
    x"25A51C8",
    x"25A4F34",
    x"25A4CA1",
    x"25A4A0E",
    x"25A477C",
    x"25A44EA",
    x"25A4259",
    x"25A3FC9",
    x"25A3D39",
    x"25A3AAA",
    x"25A381C",
    x"25A358E",
    x"25A3301",
    x"25A3075",
    x"25A2DE9",
    x"25A2B5E",
    x"25A28D3",
    x"25A2649",
    x"25A23C0",
    x"25A2138",
    x"25A1EB0",
    x"25A1C28",
    x"25A19A1",
    x"25A171B",
    x"25A1496",
    x"25A1211",
    x"25A0F8D",
    x"25A0D09",
    x"25A0A86",
    x"25A0804",
    x"25A0582",
    x"25A0301",
    x"25A0081",
    x"259FE01",
    x"259FB82",
    x"259F903",
    x"259F685",
    x"259F408",
    x"259F18B",
    x"259EF0F",
    x"259EC94",
    x"259EA19",
    x"259E79F",
    x"259E525",
    x"259E2AC",
    x"259E034",
    x"259DDBC",
    x"259DB45",
    x"259D8CE",
    x"259D659",
    x"259D3E3",
    x"259D16F",
    x"259CEFB",
    x"259CC87",
    x"259CA14",
    x"259C7A2",
    x"259C530",
    x"259C2BF",
    x"259C04F",
    x"259BDDF",
    x"259BB70",
    x"259B902",
    x"259B694",
    x"259B426",
    x"259B1BA",
    x"259AF4D",
    x"259ACE2",
    x"259AA77",
    x"259A80D",
    x"259A5A3",
    x"259A33A",
    x"259A0D1",
    x"2599E69",
    x"2599C02",
    x"259999B",
    x"2599735",
    x"25994D0",
    x"259926B",
    x"2599007",
    x"2598DA3",
    x"2598B40",
    x"25988DD",
    x"259867B",
    x"259841A",
    x"25981B9",
    x"2597F59",
    x"2597CFA",
    x"2597A9B",
    x"259783C",
    x"25975DF",
    x"2597381",
    x"2597125",
    x"2596EC9",
    x"2596C6D",
    x"2596A13",
    x"25967B8",
    x"259655F",
    x"2596306",
    x"25960AD",
    x"2595E55",
    x"2595BFE",
    x"25959A7",
    x"2595751",
    x"25954FC",
    x"25952A7",
    x"2595052",
    x"2594DFF",
    x"2594BAB",
    x"2594959",
    x"2594707",
    x"25944B5",
    x"2594264",
    x"2594014",
    x"2593DC4",
    x"2593B75",
    x"2593927",
    x"25936D9",
    x"259348B",
    x"259323E",
    x"2592FF2",
    x"2592DA6",
    x"2592B5B",
    x"2592911",
    x"25926C7",
    x"259247D",
    x"2592234",
    x"2591FEC",
    x"2591DA4",
    x"2591B5D",
    x"2591917",
    x"25916D1",
    x"259148B",
    x"2591247",
    x"2591002",
    x"2590DBF",
    x"2590B7B",
    x"2590939",
    x"25906F7",
    x"25904B5",
    x"2590274",
    x"2590034",
    x"258FDF4",
    x"258FBB5",
    x"258F976",
    x"258F738",
    x"258F4FB",
    x"258F2BE",
    x"258F081",
    x"258EE46",
    x"258EC0A",
    x"258E9D0",
    x"258E795",
    x"258E55C",
    x"258E323",
    x"258E0EA",
    x"258DEB2",
    x"258DC7B",
    x"258DA44",
    x"258D80E",
    x"258D5D8",
    x"258D3A3",
    x"258D16E",
    x"258CF3A",
    x"258CD07",
    x"258CAD4",
    x"258C8A1",
    x"258C66F",
    x"258C43E",
    x"258C20D",
    x"258BFDD",
    x"258BDAD",
    x"258BB7E",
    x"258B94F",
    x"258B721",
    x"258B4F4",
    x"258B2C7",
    x"258B09B",
    x"258AE6F",
    x"258AC43",
    x"258AA19",
    x"258A7EE",
    x"258A5C5",
    x"258A39B",
    x"258A173",
    x"2589F4B",
    x"2589D23",
    x"2589AFC",
    x"25898D6",
    x"25896B0",
    x"258948A",
    x"2589265",
    x"2589041",
    x"2588E1D",
    x"2588BFA",
    x"25889D7",
    x"25887B5",
    x"2588593",
    x"2588372",
    x"2588152",
    x"2587F32",
    x"2587D12",
    x"2587AF3",
    x"25878D5",
    x"25876B7",
    x"2587499",
    x"258727C",
    x"2587060",
    x"2586E44",
    x"2586C29",
    x"2586A0E",
    x"25867F4",
    x"25865DA",
    x"25863C1",
    x"25861A8",
    x"2585F90",
    x"2585D78",
    x"2585B61",
    x"258594B",
    x"2585735",
    x"258551F",
    x"258530A",
    x"25850F6",
    x"2584EE2",
    x"2584CCE",
    x"2584ABB",
    x"25848A9",
    x"2584697",
    x"2584486",
    x"2584275",
    x"2584064",
    x"2583E54",
    x"2583C45",
    x"2583A36",
    x"2583828",
    x"258361A",
    x"258340D",
    x"2583200",
    x"2582FF4",
    x"2582DE8",
    x"2582BDD",
    x"25829D2",
    x"25827C8",
    x"25825BE",
    x"25823B5",
    x"25821AD",
    x"2581FA4",
    x"2581D9D",
    x"2581B96",
    x"258198F",
    x"2581789",
    x"2581583",
    x"258137E",
    x"2581179",
    x"2580F75",
    x"2580D72",
    x"2580B6F",
    x"258096C",
    x"258076A",
    x"2580568",
    x"2580367",
    x"2580167",
    x"257FECD",
    x"257FACE",
    x"257F6D0",
    x"257F2D3",
    x"257EED7",
    x"257EADB",
    x"257E6E1",
    x"257E2E8",
    x"257DEF0",
    x"257DAF9",
    x"257D702",
    x"257D30D",
    x"257CF19",
    x"257CB25",
    x"257C733",
    x"257C342",
    x"257BF52",
    x"257BB62",
    x"257B774",
    x"257B386",
    x"257AF9A",
    x"257ABAF",
    x"257A7C4",
    x"257A3DB",
    x"2579FF2",
    x"2579C0B",
    x"2579824",
    x"257943F",
    x"257905A",
    x"2578C77",
    x"2578894",
    x"25784B2",
    x"25780D2",
    x"2577CF2",
    x"2577913",
    x"2577535",
    x"2577159",
    x"2576D7D",
    x"25769A2",
    x"25765C8",
    x"25761EF",
    x"2575E17",
    x"2575A40",
    x"257566A",
    x"2575295",
    x"2574EC0",
    x"2574AED",
    x"257471B",
    x"257434A",
    x"2573F79",
    x"2573BAA",
    x"25737DC",
    x"257340E",
    x"2573041",
    x"2572C76",
    x"25728AB",
    x"25724E2",
    x"2572119",
    x"2571D51",
    x"257198A",
    x"25715C4",
    x"25711FF",
    x"2570E3B",
    x"2570A78",
    x"25706B6",
    x"25702F5",
    x"256FF35",
    x"256FB75",
    x"256F7B7",
    x"256F3F9",
    x"256F03D",
    x"256EC81",
    x"256E8C7",
    x"256E50D",
    x"256E154",
    x"256DD9C",
    x"256D9E5",
    x"256D62F",
    x"256D27A",
    x"256CEC6",
    x"256CB13",
    x"256C760",
    x"256C3AF",
    x"256BFFF",
    x"256BC4F",
    x"256B8A0",
    x"256B4F3",
    x"256B146",
    x"256AD9A",
    x"256A9EF",
    x"256A645",
    x"256A29C",
    x"2569EF4",
    x"2569B4D",
    x"25697A6",
    x"2569401",
    x"256905C",
    x"2568CB9",
    x"2568916",
    x"2568574",
    x"25681D3",
    x"2567E33",
    x"2567A94",
    x"25676F6",
    x"2567359",
    x"2566FBC",
    x"2566C21",
    x"2566886",
    x"25664EC",
    x"2566154",
    x"2565DBC",
    x"2565A25",
    x"256568F",
    x"25652F9",
    x"2564F65",
    x"2564BD2",
    x"256483F",
    x"25644AE",
    x"256411D",
    x"2563D8D",
    x"25639FE",
    x"2563670",
    x"25632E3",
    x"2562F57",
    x"2562BCB",
    x"2562841",
    x"25624B7",
    x"256212E",
    x"2561DA7",
    x"2561A20",
    x"2561699",
    x"2561314",
    x"2560F90",
    x"2560C0C",
    x"256088A",
    x"2560508",
    x"2560187",
    x"255FE07",
    x"255FA88",
    x"255F70A",
    x"255F38D",
    x"255F010",
    x"255EC95",
    x"255E91A",
    x"255E5A0",
    x"255E227",
    x"255DEAF",
    x"255DB38",
    x"255D7C2",
    x"255D44C",
    x"255D0D7",
    x"255CD64",
    x"255C9F1",
    x"255C67F",
    x"255C30D",
    x"255BF9D",
    x"255BC2E",
    x"255B8BF",
    x"255B551",
    x"255B1E4",
    x"255AE78",
    x"255AB0D",
    x"255A7A3",
    x"255A439",
    x"255A0D1",
    x"2559D69",
    x"2559A02",
    x"255969C",
    x"2559337",
    x"2558FD2",
    x"2558C6F",
    x"255890C",
    x"25585AA",
    x"2558249",
    x"2557EE9",
    x"2557B8A",
    x"255782B",
    x"25574CE",
    x"2557171",
    x"2556E15",
    x"2556ABA",
    x"2556760",
    x"2556406",
    x"25560AE",
    x"2555D56",
    x"25559FF",
    x"25556A9",
    x"2555354",
    x"2554FFF",
    x"2554CAC",
    x"2554959",
    x"2554607",
    x"25542B6",
    x"2553F66",
    x"2553C16",
    x"25538C8",
    x"255357A",
    x"255322D",
    x"2552EE1",
    x"2552B95",
    x"255284B",
    x"2552501",
    x"25521B8",
    x"2551E70",
    x"2551B29",
    x"25517E3",
    x"255149D",
    x"2551158",
    x"2550E15",
    x"2550AD1",
    x"255078F",
    x"255044E",
    x"255010D",
    x"254FDCD",
    x"254FA8E",
    x"254F750",
    x"254F412",
    x"254F0D6",
    x"254ED9A",
    x"254EA5F",
    x"254E725",
    x"254E3EB",
    x"254E0B3",
    x"254DD7B",
    x"254DA44",
    x"254D70E",
    x"254D3D9",
    x"254D0A4",
    x"254CD70",
    x"254CA3D",
    x"254C70B",
    x"254C3DA",
    x"254C0A9",
    x"254BD79",
    x"254BA4A",
    x"254B71C",
    x"254B3EF",
    x"254B0C2",
    x"254AD97",
    x"254AA6C",
    x"254A741",
    x"254A418",
    x"254A0EF",
    x"2549DC7",
    x"2549AA0",
    x"254977A",
    x"2549455",
    x"2549130",
    x"2548E0C",
    x"2548AE9",
    x"25487C7",
    x"25484A5",
    x"2548184",
    x"2547E64",
    x"2547B45",
    x"2547827",
    x"2547509",
    x"25471EC",
    x"2546ED0",
    x"2546BB5",
    x"254689A",
    x"2546580",
    x"2546267",
    x"2545F4F",
    x"2545C38",
    x"2545921",
    x"254560B",
    x"25452F6",
    x"2544FE2",
    x"2544CCE",
    x"25449BB",
    x"25446A9",
    x"2544398",
    x"2544087",
    x"2543D78",
    x"2543A69",
    x"254375B",
    x"254344D",
    x"2543140",
    x"2542E34",
    x"2542B29",
    x"254281F",
    x"2542515",
    x"254220C",
    x"2541F04",
    x"2541BFD",
    x"25418F6",
    x"25415F0",
    x"25412EB",
    x"2540FE7",
    x"2540CE3",
    x"25409E0",
    x"25406DE",
    x"25403DD",
    x"25400DC",
    x"253FDDD",
    x"253FADD",
    x"253F7DF",
    x"253F4E2",
    x"253F1E5",
    x"253EEE9",
    x"253EBED",
    x"253E8F3",
    x"253E5F9",
    x"253E300",
    x"253E007",
    x"253DD10",
    x"253DA19",
    x"253D723",
    x"253D42D",
    x"253D138",
    x"253CE45",
    x"253CB51",
    x"253C85F",
    x"253C56D",
    x"253C27C",
    x"253BF8C",
    x"253BC9C",
    x"253B9AE",
    x"253B6C0",
    x"253B3D2",
    x"253B0E6",
    x"253ADFA",
    x"253AB0F",
    x"253A824",
    x"253A53B",
    x"253A252",
    x"2539F69",
    x"2539C82",
    x"253999B",
    x"25396B5",
    x"25393D0",
    x"25390EB",
    x"2538E07",
    x"2538B24",
    x"2538842",
    x"2538560",
    x"253827F",
    x"2537F9F",
    x"2537CBF",
    x"25379E0",
    x"2537702",
    x"2537425",
    x"2537148",
    x"2536E6C",
    x"2536B91",
    x"25368B6",
    x"25365DD",
    x"2536304",
    x"253602B",
    x"2535D53",
    x"2535A7C",
    x"25357A6",
    x"25354D1",
    x"25351FC",
    x"2534F28",
    x"2534C54",
    x"2534982",
    x"25346AF",
    x"25343DE",
    x"253410E",
    x"2533E3E",
    x"2533B6E",
    x"25338A0",
    x"25335D2",
    x"2533305",
    x"2533039",
    x"2532D6D",
    x"2532AA2",
    x"25327D8",
    x"253250E",
    x"2532245",
    x"2531F7D",
    x"2531CB5",
    x"25319EE",
    x"2531728",
    x"2531463",
    x"253119E",
    x"2530EDA",
    x"2530C17",
    x"2530954",
    x"2530692",
    x"25303D1",
    x"2530110",
    x"252FE50",
    x"252FB91",
    x"252F8D2",
    x"252F615",
    x"252F357",
    x"252F09B",
    x"252EDDF",
    x"252EB24",
    x"252E86A",
    x"252E5B0",
    x"252E2F7",
    x"252E03E",
    x"252DD87",
    x"252DAD0",
    x"252D819",
    x"252D563",
    x"252D2AE",
    x"252CFFA",
    x"252CD46",
    x"252CA93",
    x"252C7E1",
    x"252C530",
    x"252C27F",
    x"252BFCE",
    x"252BD1F",
    x"252BA70",
    x"252B7C1",
    x"252B514",
    x"252B267",
    x"252AFBB",
    x"252AD0F",
    x"252AA64",
    x"252A7BA",
    x"252A510",
    x"252A267",
    x"2529FBF",
    x"2529D17",
    x"2529A71",
    x"25297CA",
    x"2529525",
    x"2529280",
    x"2528FDB",
    x"2528D38",
    x"2528A95",
    x"25287F2",
    x"2528551",
    x"25282B0",
    x"252800F",
    x"2527D70",
    x"2527AD1",
    x"2527832",
    x"2527595",
    x"25272F8",
    x"252705B",
    x"2526DBF",
    x"2526B24",
    x"252688A",
    x"25265F0",
    x"2526357",
    x"25260BE",
    x"2525E26",
    x"2525B8F",
    x"25258F9",
    x"2525663",
    x"25253CD",
    x"2525139",
    x"2524EA5",
    x"2524C12",
    x"252497F",
    x"25246ED",
    x"252445B",
    x"25241CB",
    x"2523F3A",
    x"2523CAB",
    x"2523A1C",
    x"252378E",
    x"2523500",
    x"2523273",
    x"2522FE7",
    x"2522D5B",
    x"2522AD0",
    x"2522846",
    x"25225BC",
    x"2522333",
    x"25220AB",
    x"2521E23",
    x"2521B9C",
    x"2521915",
    x"252168F",
    x"252140A",
    x"2521185",
    x"2520F01",
    x"2520C7E",
    x"25209FB",
    x"2520779",
    x"25204F7",
    x"2520276",
    x"251FFF6",
    x"251FD76",
    x"251FAF7",
    x"251F879",
    x"251F5FB",
    x"251F37E",
    x"251F101",
    x"251EE85",
    x"251EC0A",
    x"251E98F",
    x"251E715",
    x"251E49C",
    x"251E223",
    x"251DFAB",
    x"251DD33",
    x"251DABC",
    x"251D846",
    x"251D5D0",
    x"251D35B",
    x"251D0E6",
    x"251CE72",
    x"251CBFF",
    x"251C98C",
    x"251C71A",
    x"251C4A9",
    x"251C238",
    x"251BFC8",
    x"251BD58",
    x"251BAE9",
    x"251B87A",
    x"251B60D",
    x"251B39F",
    x"251B133",
    x"251AEC7",
    x"251AC5B",
    x"251A9F1",
    x"251A786",
    x"251A51D",
    x"251A2B4",
    x"251A04B",
    x"2519DE4",
    x"2519B7D",
    x"2519916",
    x"25196B0",
    x"251944B",
    x"25191E6",
    x"2518F82",
    x"2518D1E",
    x"2518ABB",
    x"2518859",
    x"25185F7",
    x"2518396",
    x"2518135",
    x"2517ED5",
    x"2517C76",
    x"2517A17",
    x"25177B9",
    x"251755B",
    x"25172FE",
    x"25170A2",
    x"2516E46",
    x"2516BEA",
    x"2516990",
    x"2516736",
    x"25164DC",
    x"2516283",
    x"251602B",
    x"2515DD3",
    x"2515B7C",
    x"2515925",
    x"25156CF",
    x"251547A",
    x"2515225",
    x"2514FD1",
    x"2514D7D",
    x"2514B2A",
    x"25148D8",
    x"2514686",
    x"2514434",
    x"25141E4",
    x"2513F93",
    x"2513D44",
    x"2513AF5",
    x"25138A6",
    x"2513658",
    x"251340B",
    x"25131BE",
    x"2512F72",
    x"2512D27",
    x"2512ADC",
    x"2512891",
    x"2512647",
    x"25123FE",
    x"25121B5",
    x"2511F6D",
    x"2511D26",
    x"2511ADF",
    x"2511898",
    x"2511652",
    x"251140D",
    x"25111C8",
    x"2510F84",
    x"2510D41",
    x"2510AFE",
    x"25108BB",
    x"2510679",
    x"2510438",
    x"25101F7",
    x"250FFB7",
    x"250FD77",
    x"250FB38",
    x"250F8FA",
    x"250F6BC",
    x"250F47E",
    x"250F241",
    x"250F005",
    x"250EDC9",
    x"250EB8E",
    x"250E954",
    x"250E71A",
    x"250E4E0",
    x"250E2A7",
    x"250E06F",
    x"250DE37",
    x"250DC00",
    x"250D9C9",
    x"250D793",
    x"250D55D",
    x"250D328",
    x"250D0F4",
    x"250CEC0",
    x"250CC8C",
    x"250CA59",
    x"250C827",
    x"250C5F5",
    x"250C3C4",
    x"250C193",
    x"250BF63",
    x"250BD34",
    x"250BB05",
    x"250B8D6",
    x"250B6A8",
    x"250B47B",
    x"250B24E",
    x"250B022",
    x"250ADF6",
    x"250ABCB",
    x"250A9A0",
    x"250A776",
    x"250A54C",
    x"250A323",
    x"250A0FB",
    x"2509ED3",
    x"2509CAB",
    x"2509A84",
    x"250985E",
    x"2509638",
    x"2509413",
    x"25091EE",
    x"2508FCA",
    x"2508DA6",
    x"2508B83",
    x"2508961",
    x"250873E",
    x"250851D",
    x"25082FC",
    x"25080DB",
    x"2507EBB",
    x"2507C9C",
    x"2507A7D",
    x"250785F",
    x"2507641",
    x"2507424",
    x"2507207",
    x"2506FEB",
    x"2506DCF",
    x"2506BB4",
    x"2506999",
    x"250677F",
    x"2506565",
    x"250634C",
    x"2506134",
    x"2505F1C",
    x"2505D04",
    x"2505AED",
    x"25058D7",
    x"25056C1",
    x"25054AB",
    x"2505296",
    x"2505082",
    x"2504E6E",
    x"2504C5B",
    x"2504A48",
    x"2504836",
    x"2504624",
    x"2504413",
    x"2504202",
    x"2503FF2",
    x"2503DE2",
    x"2503BD3",
    x"25039C4",
    x"25037B6",
    x"25035A8",
    x"250339B",
    x"250318E",
    x"2502F82",
    x"2502D77",
    x"2502B6B",
    x"2502961",
    x"2502757",
    x"250254D",
    x"2502344",
    x"250213C",
    x"2501F33",
    x"2501D2C",
    x"2501B25",
    x"250191E",
    x"2501718",
    x"2501513",
    x"250130E",
    x"2501109",
    x"2500F05",
    x"2500D02",
    x"2500AFF",
    x"25008FC",
    x"25006FA",
    x"25004F9",
    x"25002F8",
    x"25000F7",
    x"24FFDEF",
    x"24FF9F0",
    x"24FF5F2",
    x"24FF1F5",
    x"24FEDF9",
    x"24FE9FE",
    x"24FE604",
    x"24FE20B",
    x"24FDE13",
    x"24FDA1C",
    x"24FD626",
    x"24FD231",
    x"24FCE3D",
    x"24FCA4A",
    x"24FC658",
    x"24FC267",
    x"24FBE77",
    x"24FBA87",
    x"24FB699",
    x"24FB2AC",
    x"24FAEC0",
    x"24FAAD5",
    x"24FA6EB",
    x"24FA301",
    x"24F9F19",
    x"24F9B32",
    x"24F974B",
    x"24F9366",
    x"24F8F82",
    x"24F8B9E",
    x"24F87BC",
    x"24F83DB",
    x"24F7FFA",
    x"24F7C1B",
    x"24F783C",
    x"24F745E",
    x"24F7082",
    x"24F6CA6",
    x"24F68CB",
    x"24F64F2",
    x"24F6119",
    x"24F5D41",
    x"24F596A",
    x"24F5594",
    x"24F51C0",
    x"24F4DEC",
    x"24F4A19",
    x"24F4647",
    x"24F4275",
    x"24F3EA5",
    x"24F3AD6",
    x"24F3708",
    x"24F333B",
    x"24F2F6E",
    x"24F2BA3",
    x"24F27D8",
    x"24F240F",
    x"24F2046",
    x"24F1C7F",
    x"24F18B8",
    x"24F14F2",
    x"24F112E",
    x"24F0D6A",
    x"24F09A7",
    x"24F05E5",
    x"24F0224",
    x"24EFE64",
    x"24EFAA5",
    x"24EF6E7",
    x"24EF329",
    x"24EEF6D",
    x"24EEBB2",
    x"24EE7F7",
    x"24EE43E",
    x"24EE085",
    x"24EDCCD",
    x"24ED917",
    x"24ED561",
    x"24ED1AC",
    x"24ECDF8",
    x"24ECA45",
    x"24EC693",
    x"24EC2E2",
    x"24EBF31",
    x"24EBB82",
    x"24EB7D4",
    x"24EB426",
    x"24EB07A",
    x"24EACCE",
    x"24EA923",
    x"24EA579",
    x"24EA1D1",
    x"24E9E29",
    x"24E9A81",
    x"24E96DB",
    x"24E9336",
    x"24E8F92",
    x"24E8BEE",
    x"24E884C",
    x"24E84AA",
    x"24E8109",
    x"24E7D6A",
    x"24E79CB",
    x"24E762D",
    x"24E7290",
    x"24E6EF3",
    x"24E6B58",
    x"24E67BE",
    x"24E6424",
    x"24E608C",
    x"24E5CF4",
    x"24E595D",
    x"24E55C7",
    x"24E5232",
    x"24E4E9E",
    x"24E4B0B",
    x"24E4779",
    x"24E43E7",
    x"24E4057",
    x"24E3CC7",
    x"24E3938",
    x"24E35AA",
    x"24E321D",
    x"24E2E91",
    x"24E2B06",
    x"24E277C",
    x"24E23F2",
    x"24E206A",
    x"24E1CE2",
    x"24E195B",
    x"24E15D6",
    x"24E1251",
    x"24E0ECC",
    x"24E0B49",
    x"24E07C7",
    x"24E0445",
    x"24E00C5",
    x"24DFD45",
    x"24DF9C6",
    x"24DF648",
    x"24DF2CB",
    x"24DEF4F",
    x"24DEBD3",
    x"24DE859",
    x"24DE4DF",
    x"24DE166",
    x"24DDDEE",
    x"24DDA77",
    x"24DD701",
    x"24DD38C",
    x"24DD017",
    x"24DCCA4",
    x"24DC931",
    x"24DC5BF",
    x"24DC24E",
    x"24DBEDE",
    x"24DBB6F",
    x"24DB800",
    x"24DB493",
    x"24DB126",
    x"24DADBA",
    x"24DAA4F",
    x"24DA6E5",
    x"24DA37C",
    x"24DA013",
    x"24D9CAC",
    x"24D9945",
    x"24D95DF",
    x"24D927A",
    x"24D8F16",
    x"24D8BB2",
    x"24D8850",
    x"24D84EE",
    x"24D818D",
    x"24D7E2D",
    x"24D7ACE",
    x"24D7770",
    x"24D7413",
    x"24D70B6",
    x"24D6D5A",
    x"24D69FF",
    x"24D66A5",
    x"24D634C",
    x"24D5FF4",
    x"24D5C9C",
    x"24D5945",
    x"24D55EF",
    x"24D529A",
    x"24D4F46",
    x"24D4BF3",
    x"24D48A0",
    x"24D454E",
    x"24D41FD",
    x"24D3EAD",
    x"24D3B5E",
    x"24D3810",
    x"24D34C2",
    x"24D3175",
    x"24D2E29",
    x"24D2ADE",
    x"24D2794",
    x"24D244A",
    x"24D2102",
    x"24D1DBA",
    x"24D1A73",
    x"24D172D",
    x"24D13E7",
    x"24D10A3",
    x"24D0D5F",
    x"24D0A1C",
    x"24D06DA",
    x"24D0399",
    x"24D0058",
    x"24CFD18",
    x"24CF9DA",
    x"24CF69C",
    x"24CF35E",
    x"24CF022",
    x"24CECE6",
    x"24CE9AB",
    x"24CE671",
    x"24CE338",
    x"24CE000",
    x"24CDCC8",
    x"24CD991",
    x"24CD65B",
    x"24CD326",
    x"24CCFF2",
    x"24CCCBE",
    x"24CC98B",
    x"24CC659",
    x"24CC328",
    x"24CBFF8",
    x"24CBCC8",
    x"24CB999",
    x"24CB66B",
    x"24CB33E",
    x"24CB012",
    x"24CACE6",
    x"24CA9BB",
    x"24CA691",
    x"24CA368",
    x"24CA040",
    x"24C9D18",
    x"24C99F1",
    x"24C96CB",
    x"24C93A6",
    x"24C9081",
    x"24C8D5D",
    x"24C8A3B",
    x"24C8718",
    x"24C83F7",
    x"24C80D6",
    x"24C7DB7",
    x"24C7A98",
    x"24C7779",
    x"24C745C",
    x"24C713F",
    x"24C6E23",
    x"24C6B08",
    x"24C67EE",
    x"24C64D4",
    x"24C61BB",
    x"24C5EA3",
    x"24C5B8C",
    x"24C5875",
    x"24C5560",
    x"24C524B",
    x"24C4F37",
    x"24C4C23",
    x"24C4910",
    x"24C45FF",
    x"24C42ED",
    x"24C3FDD",
    x"24C3CCE",
    x"24C39BF",
    x"24C36B1",
    x"24C33A3",
    x"24C3097",
    x"24C2D8B",
    x"24C2A80",
    x"24C2776",
    x"24C246C",
    x"24C2164",
    x"24C1E5C",
    x"24C1B54",
    x"24C184E",
    x"24C1548",
    x"24C1243",
    x"24C0F3F",
    x"24C0C3C",
    x"24C0939",
    x"24C0637",
    x"24C0336",
    x"24C0035",
    x"24BFD36",
    x"24BFA37",
    x"24BF739",
    x"24BF43B",
    x"24BF13F",
    x"24BEE43",
    x"24BEB47",
    x"24BE84D",
    x"24BE553",
    x"24BE25A",
    x"24BDF62",
    x"24BDC6B",
    x"24BD974",
    x"24BD67E",
    x"24BD389",
    x"24BD094",
    x"24BCDA0",
    x"24BCAAD",
    x"24BC7BB",
    x"24BC4C9",
    x"24BC1D9",
    x"24BBEE9",
    x"24BBBF9",
    x"24BB90B",
    x"24BB61D",
    x"24BB32F",
    x"24BB043",
    x"24BAD57",
    x"24BAA6C",
    x"24BA782",
    x"24BA499",
    x"24BA1B0",
    x"24B9EC8",
    x"24B9BE0",
    x"24B98FA",
    x"24B9614",
    x"24B932F",
    x"24B904A",
    x"24B8D67",
    x"24B8A84",
    x"24B87A1",
    x"24B84C0",
    x"24B81DF",
    x"24B7EFF",
    x"24B7C20",
    x"24B7941",
    x"24B7663",
    x"24B7386",
    x"24B70A9",
    x"24B6DCD",
    x"24B6AF2",
    x"24B6818",
    x"24B653E",
    x"24B6265",
    x"24B5F8D",
    x"24B5CB5",
    x"24B59DF",
    x"24B5709",
    x"24B5433",
    x"24B515E",
    x"24B4E8A",
    x"24B4BB7",
    x"24B48E5",
    x"24B4613",
    x"24B4342",
    x"24B4071",
    x"24B3DA1",
    x"24B3AD2",
    x"24B3804",
    x"24B3536",
    x"24B3269",
    x"24B2F9D",
    x"24B2CD1",
    x"24B2A07",
    x"24B273C",
    x"24B2473",
    x"24B21AA",
    x"24B1EE2",
    x"24B1C1B",
    x"24B1954",
    x"24B168E",
    x"24B13C9",
    x"24B1104",
    x"24B0E40",
    x"24B0B7D",
    x"24B08BB",
    x"24B05F9",
    x"24B0338",
    x"24B0077",
    x"24AFDB7",
    x"24AFAF8",
    x"24AF83A",
    x"24AF57C",
    x"24AF2BF",
    x"24AF003",
    x"24AED47",
    x"24AEA8C",
    x"24AE7D2",
    x"24AE518",
    x"24AE25F",
    x"24ADFA7",
    x"24ADCEF",
    x"24ADA39",
    x"24AD782",
    x"24AD4CD",
    x"24AD218",
    x"24ACF64",
    x"24ACCB0",
    x"24AC9FD",
    x"24AC74B",
    x"24AC49A",
    x"24AC1E9",
    x"24ABF39",
    x"24ABC89",
    x"24AB9DB",
    x"24AB72C",
    x"24AB47F",
    x"24AB1D2",
    x"24AAF26",
    x"24AAC7B",
    x"24AA9D0",
    x"24AA726",
    x"24AA47C",
    x"24AA1D3",
    x"24A9F2B",
    x"24A9C84",
    x"24A99DD",
    x"24A9737",
    x"24A9491",
    x"24A91ED",
    x"24A8F48",
    x"24A8CA5",
    x"24A8A02",
    x"24A8760",
    x"24A84BE",
    x"24A821E",
    x"24A7F7D",
    x"24A7CDE",
    x"24A7A3F",
    x"24A77A1",
    x"24A7503",
    x"24A7266",
    x"24A6FCA",
    x"24A6D2E",
    x"24A6A93",
    x"24A67F9",
    x"24A655F",
    x"24A62C6",
    x"24A602E",
    x"24A5D96",
    x"24A5AFF",
    x"24A5869",
    x"24A55D3",
    x"24A533E",
    x"24A50A9",
    x"24A4E16",
    x"24A4B82",
    x"24A48F0",
    x"24A465E",
    x"24A43CD",
    x"24A413C",
    x"24A3EAC",
    x"24A3C1D",
    x"24A398E",
    x"24A3700",
    x"24A3472",
    x"24A31E6",
    x"24A2F59",
    x"24A2CCE",
    x"24A2A43",
    x"24A27B9",
    x"24A252F",
    x"24A22A6",
    x"24A201E",
    x"24A1D96",
    x"24A1B0F",
    x"24A1889",
    x"24A1603",
    x"24A137E",
    x"24A10F9",
    x"24A0E75",
    x"24A0BF2",
    x"24A096F",
    x"24A06ED",
    x"24A046C",
    x"24A01EB",
    x"249FF6B",
    x"249FCEB",
    x"249FA6C",
    x"249F7EE",
    x"249F570",
    x"249F2F3",
    x"249F077",
    x"249EDFB",
    x"249EB80",
    x"249E905",
    x"249E68B",
    x"249E412",
    x"249E199",
    x"249DF21",
    x"249DCAA",
    x"249DA33",
    x"249D7BD",
    x"249D547",
    x"249D2D2",
    x"249D05E",
    x"249CDEA",
    x"249CB77",
    x"249C904",
    x"249C692",
    x"249C421",
    x"249C1B0",
    x"249BF40",
    x"249BCD0",
    x"249BA62",
    x"249B7F3",
    x"249B586",
    x"249B318",
    x"249B0AC",
    x"249AE40",
    x"249ABD5",
    x"249A96A",
    x"249A700",
    x"249A497",
    x"249A22E",
    x"2499FC6",
    x"2499D5E",
    x"2499AF7",
    x"2499891",
    x"249962B",
    x"24993C5",
    x"2499161",
    x"2498EFD",
    x"2498C99",
    x"2498A36",
    x"24987D4",
    x"2498573",
    x"2498311",
    x"24980B1",
    x"2497E51",
    x"2497BF2",
    x"2497993",
    x"2497735",
    x"24974D8",
    x"249727B",
    x"249701E",
    x"2496DC3",
    x"2496B67",
    x"249690D",
    x"24966B3",
    x"249645A",
    x"2496201",
    x"2495FA9",
    x"2495D51",
    x"2495AFA",
    x"24958A3",
    x"249564E",
    x"24953F8",
    x"24951A4",
    x"2494F4F",
    x"2494CFC",
    x"2494AA9",
    x"2494857",
    x"2494605",
    x"24943B4",
    x"2494163",
    x"2493F13",
    x"2493CC3",
    x"2493A74",
    x"2493826",
    x"24935D8",
    x"249338B",
    x"249313F",
    x"2492EF3",
    x"2492CA7",
    x"2492A5C",
    x"2492812",
    x"24925C8",
    x"249237F",
    x"2492136",
    x"2491EEE",
    x"2491CA7",
    x"2491A60",
    x"249181A",
    x"24915D4",
    x"249138F",
    x"249114A",
    x"2490F06",
    x"2490CC3",
    x"2490A80",
    x"249083E",
    x"24905FC",
    x"24903BB",
    x"249017A",
    x"248FF3A",
    x"248FCFA",
    x"248FABB",
    x"248F87D",
    x"248F63F",
    x"248F402",
    x"248F1C5",
    x"248EF89",
    x"248ED4D",
    x"248EB12",
    x"248E8D8",
    x"248E69E",
    x"248E464",
    x"248E22C",
    x"248DFF3",
    x"248DDBC",
    x"248DB84",
    x"248D94E",
    x"248D718",
    x"248D4E2",
    x"248D2AD",
    x"248D079",
    x"248CE45",
    x"248CC12",
    x"248C9DF",
    x"248C7AD",
    x"248C57B",
    x"248C34A",
    x"248C11A",
    x"248BEEA",
    x"248BCBA",
    x"248BA8B",
    x"248B85D",
    x"248B62F",
    x"248B402",
    x"248B1D5",
    x"248AFA9",
    x"248AD7D",
    x"248AB52",
    x"248A928",
    x"248A6FE",
    x"248A4D4",
    x"248A2AB",
    x"248A083",
    x"2489E5B",
    x"2489C34",
    x"2489A0D",
    x"24897E7",
    x"24895C1",
    x"248939C",
    x"2489177",
    x"2488F53",
    x"2488D2F",
    x"2488B0C",
    x"24888EA",
    x"24886C8",
    x"24884A6",
    x"2488286",
    x"2488065",
    x"2487E45",
    x"2487C26",
    x"2487A07",
    x"24877E9",
    x"24875CB",
    x"24873AE",
    x"2487191",
    x"2486F75",
    x"2486D5A",
    x"2486B3F",
    x"2486924",
    x"248670A",
    x"24864F1",
    x"24862D8",
    x"24860BF",
    x"2485EA7",
    x"2485C90",
    x"2485A79",
    x"2485863",
    x"248564D",
    x"2485437",
    x"2485223",
    x"248500E",
    x"2484DFB",
    x"2484BE7",
    x"24849D5",
    x"24847C3",
    x"24845B1",
    x"24843A0",
    x"248418F",
    x"2483F7F",
    x"2483D6F",
    x"2483B60",
    x"2483952",
    x"2483744",
    x"2483536",
    x"2483329",
    x"248311C",
    x"2482F10",
    x"2482D05",
    x"2482AFA",
    x"24828EF",
    x"24826E5",
    x"24824DC",
    x"24822D3",
    x"24820CA",
    x"2481EC3",
    x"2481CBB",
    x"2481AB4",
    x"24818AE",
    x"24816A8",
    x"24814A2",
    x"248129E",
    x"2481099",
    x"2480E95",
    x"2480C92",
    x"2480A8F",
    x"248088D",
    x"248068B",
    x"2480489",
    x"2480288",
    x"2480088",
    x"247FD11",
    x"247F912",
    x"247F514",
    x"247F117",
    x"247ED1C",
    x"247E921",
    x"247E527",
    x"247E12E",
    x"247DD36",
    x"247D940",
    x"247D54A",
    x"247D155",
    x"247CD61",
    x"247C96E",
    x"247C57C",
    x"247C18C",
    x"247BD9C",
    x"247B9AD",
    x"247B5BF",
    x"247B1D2",
    x"247ADE6",
    x"247A9FB",
    x"247A611",
    x"247A228",
    x"2479E40",
    x"2479A59",
    x"2479673",
    x"247928E",
    x"2478EA9",
    x"2478AC6",
    x"24786E4",
    x"2478303",
    x"2477F23",
    x"2477B43",
    x"2477765",
    x"2477388",
    x"2476FAB",
    x"2476BD0",
    x"24767F5",
    x"247641C",
    x"2476043",
    x"2475C6C",
    x"2475895",
    x"24754BF",
    x"24750EB",
    x"2474D17",
    x"2474944",
    x"2474572",
    x"24741A1",
    x"2473DD1",
    x"2473A02",
    x"2473634",
    x"2473267",
    x"2472E9B",
    x"2472AD0",
    x"2472706",
    x"247233C",
    x"2471F74",
    x"2471BAD",
    x"24717E6",
    x"2471421",
    x"247105C",
    x"2470C99",
    x"24708D6",
    x"2470514",
    x"2470153",
    x"246FD94",
    x"246F9D5",
    x"246F617",
    x"246F25A",
    x"246EE9D",
    x"246EAE2",
    x"246E728",
    x"246E36F",
    x"246DFB6",
    x"246DBFF",
    x"246D848",
    x"246D493",
    x"246D0DE",
    x"246CD2A",
    x"246C977",
    x"246C5C5",
    x"246C215",
    x"246BE64",
    x"246BAB5",
    x"246B707",
    x"246B35A",
    x"246AFAD",
    x"246AC02",
    x"246A857",
    x"246A4AE",
    x"246A105",
    x"2469D5D",
    x"24699B6",
    x"2469610",
    x"246926B",
    x"2468EC7",
    x"2468B24",
    x"2468782",
    x"24683E0",
    x"2468040",
    x"2467CA0",
    x"2467901",
    x"2467564",
    x"24671C7",
    x"2466E2B",
    x"2466A90",
    x"24666F5",
    x"246635C",
    x"2465FC4",
    x"2465C2C",
    x"2465896",
    x"2465500",
    x"246516B",
    x"2464DD7",
    x"2464A44",
    x"24646B2",
    x"2464321",
    x"2463F91",
    x"2463C01",
    x"2463873",
    x"24634E5",
    x"2463158",
    x"2462DCC",
    x"2462A41",
    x"24626B7",
    x"246232E",
    x"2461FA5",
    x"2461C1E",
    x"2461897",
    x"2461512",
    x"246118D",
    x"2460E09",
    x"2460A86",
    x"2460704",
    x"2460382",
    x"2460002",
    x"245FC82",
    x"245F904",
    x"245F586",
    x"245F209",
    x"245EE8D",
    x"245EB12",
    x"245E797",
    x"245E41E",
    x"245E0A5",
    x"245DD2D",
    x"245D9B7",
    x"245D641",
    x"245D2CB",
    x"245CF57",
    x"245CBE4",
    x"245C871",
    x"245C500",
    x"245C18F",
    x"245BE1F",
    x"245BAB0",
    x"245B741",
    x"245B3D4",
    x"245B068",
    x"245ACFC",
    x"245A991",
    x"245A627",
    x"245A2BE",
    x"2459F56",
    x"2459BEE",
    x"2459888",
    x"2459522",
    x"24591BD",
    x"2458E59",
    x"2458AF6",
    x"2458794",
    x"2458432",
    x"24580D2",
    x"2457D72",
    x"2457A13",
    x"24576B5",
    x"2457358",
    x"2456FFB",
    x"2456CA0",
    x"2456945",
    x"24565EB",
    x"2456292",
    x"2455F3A",
    x"2455BE2",
    x"245588C",
    x"2455536",
    x"24551E1",
    x"2454E8D",
    x"2454B3A",
    x"24547E7",
    x"2454496",
    x"2454145",
    x"2453DF5",
    x"2453AA6",
    x"2453758",
    x"245340A",
    x"24530BE",
    x"2452D72",
    x"2452A27",
    x"24526DD",
    x"2452394",
    x"245204B",
    x"2451D04",
    x"24519BD",
    x"2451677",
    x"2451331",
    x"2450FED",
    x"2450CAA",
    x"2450967",
    x"2450625",
    x"24502E4",
    x"244FFA3",
    x"244FC64",
    x"244F925",
    x"244F5E7",
    x"244F2AA",
    x"244EF6E",
    x"244EC32",
    x"244E8F8",
    x"244E5BE",
    x"244E285",
    x"244DF4D",
    x"244DC15",
    x"244D8DF",
    x"244D5A9",
    x"244D274",
    x"244CF40",
    x"244CC0C",
    x"244C8DA",
    x"244C5A8",
    x"244C277",
    x"244BF47",
    x"244BC17",
    x"244B8E9",
    x"244B5BB",
    x"244B28E",
    x"244AF61",
    x"244AC36",
    x"244A90B",
    x"244A5E1",
    x"244A2B8",
    x"2449F90",
    x"2449C69",
    x"2449942",
    x"244961C",
    x"24492F7",
    x"2448FD2",
    x"2448CAF",
    x"244898C",
    x"244866A",
    x"2448349",
    x"2448029",
    x"2447D09",
    x"24479EA",
    x"24476CC",
    x"24473AF",
    x"2447092",
    x"2446D76",
    x"2446A5B",
    x"2446741",
    x"2446428",
    x"244610F",
    x"2445DF7",
    x"2445AE0",
    x"24457CA",
    x"24454B4",
    x"244519F",
    x"2444E8B",
    x"2444B78",
    x"2444866",
    x"2444554",
    x"2444243",
    x"2443F33",
    x"2443C23",
    x"2443915",
    x"2443607",
    x"24432FA",
    x"2442FED",
    x"2442CE2",
    x"24429D7",
    x"24426CD",
    x"24423C3",
    x"24420BB",
    x"2441DB3",
    x"2441AAC",
    x"24417A6",
    x"24414A0",
    x"244119B",
    x"2440E97",
    x"2440B94",
    x"2440892",
    x"2440590",
    x"244028F",
    x"243FF8F",
    x"243FC8F",
    x"243F990",
    x"243F692",
    x"243F395",
    x"243F099",
    x"243ED9D",
    x"243EAA2",
    x"243E7A7",
    x"243E4AE",
    x"243E1B5",
    x"243DEBD",
    x"243DBC6",
    x"243D8CF",
    x"243D5D9",
    x"243D2E4",
    x"243CFF0",
    x"243CCFC",
    x"243CA09",
    x"243C717",
    x"243C426",
    x"243C135",
    x"243BE45",
    x"243BB56",
    x"243B868",
    x"243B57A",
    x"243B28D",
    x"243AFA1",
    x"243ACB5",
    x"243A9CA",
    x"243A6E0",
    x"243A3F7",
    x"243A10E",
    x"2439E26",
    x"2439B3F",
    x"2439859",
    x"2439573",
    x"243928E",
    x"2438FAA",
    x"2438CC6",
    x"24389E3",
    x"2438701",
    x"2438420",
    x"243813F",
    x"2437E5F",
    x"2437B80",
    x"24378A1",
    x"24375C4",
    x"24372E6",
    x"243700A",
    x"2436D2E",
    x"2436A53",
    x"2436779",
    x"24364A0",
    x"24361C7",
    x"2435EEF",
    x"2435C17",
    x"2435941",
    x"243566B",
    x"2435396",
    x"24350C1",
    x"2434DED",
    x"2434B1A",
    x"2434848",
    x"2434576",
    x"24342A5",
    x"2433FD5",
    x"2433D05",
    x"2433A36",
    x"2433768",
    x"243349A",
    x"24331CE",
    x"2432F01",
    x"2432C36",
    x"243296B",
    x"24326A1",
    x"24323D8",
    x"243210F",
    x"2431E48",
    x"2431B80",
    x"24318BA",
    x"24315F4",
    x"243132F",
    x"243106A",
    x"2430DA7",
    x"2430AE4",
    x"2430821",
    x"243055F",
    x"243029E",
    x"242FFDE",
    x"242FD1F",
    x"242FA60",
    x"242F7A1",
    x"242F4E4",
    x"242F227",
    x"242EF6B",
    x"242ECAF",
    x"242E9F4",
    x"242E73A",
    x"242E481",
    x"242E1C8",
    x"242DF10",
    x"242DC58",
    x"242D9A2",
    x"242D6EC",
    x"242D436",
    x"242D182",
    x"242CECD",
    x"242CC1A",
    x"242C967",
    x"242C6B5",
    x"242C404",
    x"242C153",
    x"242BEA3",
    x"242BBF4",
    x"242B945",
    x"242B697",
    x"242B3EA",
    x"242B13D",
    x"242AE91",
    x"242ABE6",
    x"242A93C",
    x"242A692",
    x"242A3E8",
    x"242A140",
    x"2429E98",
    x"2429BF0",
    x"242994A",
    x"24296A4",
    x"24293FE",
    x"242915A",
    x"2428EB6",
    x"2428C12",
    x"2428970",
    x"24286CE",
    x"242842C",
    x"242818C",
    x"2427EEB",
    x"2427C4C",
    x"24279AD",
    x"242770F",
    x"2427472",
    x"24271D5",
    x"2426F39",
    x"2426C9D",
    x"2426A03",
    x"2426768",
    x"24264CF",
    x"2426236",
    x"2425F9E",
    x"2425D06",
    x"2425A6F",
    x"24257D9",
    x"2425543",
    x"24252AE",
    x"242501A",
    x"2424D86",
    x"2424AF3",
    x"2424861",
    x"24245CF",
    x"242433E",
    x"24240AD",
    x"2423E1E",
    x"2423B8E",
    x"2423900",
    x"2423672",
    x"24233E5",
    x"2423158",
    x"2422ECC",
    x"2422C40",
    x"24229B6",
    x"242272C",
    x"24224A2",
    x"2422219",
    x"2421F91",
    x"2421D0A",
    x"2421A83",
    x"24217FC",
    x"2421577",
    x"24212F2",
    x"242106D",
    x"2420DE9",
    x"2420B66",
    x"24208E4",
    x"2420662",
    x"24203E0",
    x"2420160",
    x"241FEE0",
    x"241FC60",
    x"241F9E2",
    x"241F763",
    x"241F4E6",
    x"241F269",
    x"241EFED",
    x"241ED71",
    x"241EAF6",
    x"241E87B",
    x"241E602",
    x"241E388",
    x"241E110",
    x"241DE98",
    x"241DC21",
    x"241D9AA",
    x"241D734",
    x"241D4BE",
    x"241D249",
    x"241CFD5",
    x"241CD61",
    x"241CAEE",
    x"241C87C",
    x"241C60A",
    x"241C399",
    x"241C128",
    x"241BEB8",
    x"241BC49",
    x"241B9DA",
    x"241B76C",
    x"241B4FF",
    x"241B292",
    x"241B025",
    x"241ADBA",
    x"241AB4E",
    x"241A8E4",
    x"241A67A",
    x"241A411",
    x"241A1A8",
    x"2419F40",
    x"2419CD8",
    x"2419A71",
    x"241980B",
    x"24195A5",
    x"2419340",
    x"24190DC",
    x"2418E78",
    x"2418C15",
    x"24189B2",
    x"2418750",
    x"24184EE",
    x"241828D",
    x"241802D",
    x"2417DCD",
    x"2417B6E",
    x"241790F",
    x"24176B1",
    x"2417454",
    x"24171F7",
    x"2416F9B",
    x"2416D3F",
    x"2416AE4",
    x"241688A",
    x"2416630",
    x"24163D7",
    x"241617E",
    x"2415F26",
    x"2415CCF",
    x"2415A78",
    x"2415821",
    x"24155CC",
    x"2415377",
    x"2415122",
    x"2414ECE",
    x"2414C7B",
    x"2414A28",
    x"24147D5",
    x"2414584",
    x"2414333",
    x"24140E2",
    x"2413E92",
    x"2413C43",
    x"24139F4",
    x"24137A6",
    x"2413558",
    x"241330B",
    x"24130BF",
    x"2412E73",
    x"2412C28",
    x"24129DD",
    x"2412793",
    x"2412549",
    x"2412300",
    x"24120B8",
    x"2411E70",
    x"2411C28",
    x"24119E2",
    x"241179B",
    x"2411556",
    x"2411311",
    x"24110CC",
    x"2410E88",
    x"2410C45",
    x"2410A02",
    x"24107C0",
    x"241057E",
    x"241033D",
    x"24100FD",
    x"240FEBD",
    x"240FC7D",
    x"240FA3E",
    x"240F800",
    x"240F5C2",
    x"240F385",
    x"240F149",
    x"240EF0D",
    x"240ECD1",
    x"240EA96",
    x"240E85C",
    x"240E622",
    x"240E3E9",
    x"240E1B0",
    x"240DF78",
    x"240DD40",
    x"240DB09",
    x"240D8D3",
    x"240D69D",
    x"240D468",
    x"240D233",
    x"240CFFE",
    x"240CDCB",
    x"240CB98",
    x"240C965",
    x"240C733",
    x"240C501",
    x"240C2D0",
    x"240C0A0",
    x"240BE70",
    x"240BC41",
    x"240BA12",
    x"240B7E4",
    x"240B5B6",
    x"240B389",
    x"240B15C",
    x"240AF30",
    x"240AD05",
    x"240AADA",
    x"240A8AF",
    x"240A685",
    x"240A45C",
    x"240A233",
    x"240A00B",
    x"2409DE3",
    x"2409BBC",
    x"2409995",
    x"240976F",
    x"2409549",
    x"2409324",
    x"2409100",
    x"2408EDC",
    x"2408CB8",
    x"2408A96",
    x"2408873",
    x"2408651",
    x"2408430",
    x"240820F",
    x"2407FEF",
    x"2407DCF",
    x"2407BB0",
    x"2407991",
    x"2407773",
    x"2407556",
    x"2407339",
    x"240711C",
    x"2406F00",
    x"2406CE5",
    x"2406ACA",
    x"24068AF",
    x"2406695",
    x"240647C",
    x"2406263",
    x"240604B",
    x"2405E33",
    x"2405C1C",
    x"2405A05",
    x"24057EF",
    x"24055D9",
    x"24053C4",
    x"24051AF",
    x"2404F9B",
    x"2404D87",
    x"2404B74",
    x"2404961",
    x"240474F",
    x"240453E",
    x"240432D",
    x"240411C",
    x"2403F0C",
    x"2403CFD",
    x"2403AEE",
    x"24038DF",
    x"24036D1",
    x"24034C4",
    x"24032B7",
    x"24030AA",
    x"2402E9F",
    x"2402C93",
    x"2402A88",
    x"240287E",
    x"2402674",
    x"240246B",
    x"2402262",
    x"2402059",
    x"2401E52",
    x"2401C4A",
    x"2401A43",
    x"240183D",
    x"2401637",
    x"2401432",
    x"240122D",
    x"2401029",
    x"2400E25",
    x"2400C22",
    x"2400A1F",
    x"240081D",
    x"240061B",
    x"240041A",
    x"2400219",
    x"2400019",
    x"23FFC32",
    x"23FF834",
    x"23FF436",
    x"23FF03A",
    x"23FEC3E",
    x"23FE844",
    x"23FE44A",
    x"23FE051",
    x"23FDC5A",
    x"23FD863",
    x"23FD46E",
    x"23FD079",
    x"23FCC85",
    x"23FC893",
    x"23FC4A1",
    x"23FC0B0",
    x"23FBCC1",
    x"23FB8D2",
    x"23FB4E4",
    x"23FB0F8",
    x"23FAD0C",
    x"23FA921",
    x"23FA537",
    x"23FA14F",
    x"23F9D67",
    x"23F9980",
    x"23F959A",
    x"23F91B5",
    x"23F8DD1",
    x"23F89EE",
    x"23F860C",
    x"23F822B",
    x"23F7E4B",
    x"23F7A6C",
    x"23F768E",
    x"23F72B1",
    x"23F6ED4",
    x"23F6AF9",
    x"23F671F",
    x"23F6346",
    x"23F5F6D",
    x"23F5B96",
    x"23F57C0",
    x"23F53EA",
    x"23F5016",
    x"23F4C42",
    x"23F486F",
    x"23F449E",
    x"23F40CD",
    x"23F3CFD",
    x"23F392F",
    x"23F3561",
    x"23F3194",
    x"23F2DC8",
    x"23F29FD",
    x"23F2633",
    x"23F226A",
    x"23F1EA2",
    x"23F1ADB",
    x"23F1714",
    x"23F134F",
    x"23F0F8B",
    x"23F0BC7",
    x"23F0805",
    x"23F0443",
    x"23F0083",
    x"23EFCC3",
    x"23EF904",
    x"23EF547",
    x"23EF18A",
    x"23EEDCE",
    x"23EEA13",
    x"23EE659",
    x"23EE2A0",
    x"23EDEE7",
    x"23EDB30",
    x"23ED77A",
    x"23ED3C4",
    x"23ED010",
    x"23ECC5C",
    x"23EC8AA",
    x"23EC4F8",
    x"23EC147",
    x"23EBD97",
    x"23EB9E8",
    x"23EB63A",
    x"23EB28D",
    x"23EAEE1",
    x"23EAB36",
    x"23EA78C",
    x"23EA3E2",
    x"23EA03A",
    x"23E9C92",
    x"23E98EB",
    x"23E9546",
    x"23E91A1",
    x"23E8DFD",
    x"23E8A5A",
    x"23E86B8",
    x"23E8316",
    x"23E7F76",
    x"23E7BD7",
    x"23E7838",
    x"23E749B",
    x"23E70FE",
    x"23E6D62",
    x"23E69C7",
    x"23E662D",
    x"23E6294",
    x"23E5EFC",
    x"23E5B65",
    x"23E57CE",
    x"23E5439",
    x"23E50A4",
    x"23E4D10",
    x"23E497E",
    x"23E45EC",
    x"23E425B",
    x"23E3ECA",
    x"23E3B3B",
    x"23E37AD",
    x"23E341F",
    x"23E3093",
    x"23E2D07",
    x"23E297C",
    x"23E25F2",
    x"23E2269",
    x"23E1EE1",
    x"23E1B5A",
    x"23E17D3",
    x"23E144E",
    x"23E10C9",
    x"23E0D45",
    x"23E09C3",
    x"23E0641",
    x"23E02BF",
    x"23DFF3F",
    x"23DFBC0",
    x"23DF841",
    x"23DF4C4",
    x"23DF147",
    x"23DEDCB",
    x"23DEA50",
    x"23DE6D6",
    x"23DE35D",
    x"23DDFE4",
    x"23DDC6D",
    x"23DD8F6",
    x"23DD580",
    x"23DD20B",
    x"23DCE97",
    x"23DCB24",
    x"23DC7B2",
    x"23DC440",
    x"23DC0D0",
    x"23DBD60",
    x"23DB9F1",
    x"23DB683",
    x"23DB316",
    x"23DAFA9",
    x"23DAC3E",
    x"23DA8D3",
    x"23DA569",
    x"23DA200",
    x"23D9E98",
    x"23D9B31",
    x"23D97CB",
    x"23D9465",
    x"23D9101",
    x"23D8D9D",
    x"23D8A3A",
    x"23D86D8",
    x"23D8376",
    x"23D8016",
    x"23D7CB6",
    x"23D7957",
    x"23D75FA",
    x"23D729C",
    x"23D6F40",
    x"23D6BE5",
    x"23D688A",
    x"23D6531",
    x"23D61D8",
    x"23D5E80",
    x"23D5B28",
    x"23D57D2",
    x"23D547D",
    x"23D5128",
    x"23D4DD4",
    x"23D4A81",
    x"23D472F",
    x"23D43DD",
    x"23D408D",
    x"23D3D3D",
    x"23D39EE",
    x"23D36A0",
    x"23D3353",
    x"23D3006",
    x"23D2CBB",
    x"23D2970",
    x"23D2626",
    x"23D22DD",
    x"23D1F95",
    x"23D1C4D",
    x"23D1907",
    x"23D15C1",
    x"23D127C",
    x"23D0F37",
    x"23D0BF4",
    x"23D08B1",
    x"23D0570",
    x"23D022F",
    x"23CFEEF",
    x"23CFBAF",
    x"23CF871",
    x"23CF533",
    x"23CF1F6",
    x"23CEEBA",
    x"23CEB7F",
    x"23CE844",
    x"23CE50B",
    x"23CE1D2",
    x"23CDE9A",
    x"23CDB63",
    x"23CD82C",
    x"23CD4F6",
    x"23CD1C2",
    x"23CCE8E",
    x"23CCB5A",
    x"23CC828",
    x"23CC4F6",
    x"23CC1C5",
    x"23CBE95",
    x"23CBB66",
    x"23CB838",
    x"23CB50A",
    x"23CB1DD",
    x"23CAEB1",
    x"23CAB86",
    x"23CA85B",
    x"23CA532",
    x"23CA209",
    x"23C9EE1",
    x"23C9BB9",
    x"23C9893",
    x"23C956D",
    x"23C9248",
    x"23C8F24",
    x"23C8C00",
    x"23C88DE",
    x"23C85BC",
    x"23C829B",
    x"23C7F7B",
    x"23C7C5B",
    x"23C793D",
    x"23C761F",
    x"23C7301",
    x"23C6FE5",
    x"23C6CC9",
    x"23C69AF",
    x"23C6695",
    x"23C637B",
    x"23C6063",
    x"23C5D4B",
    x"23C5A34",
    x"23C571E",
    x"23C5409",
    x"23C50F4",
    x"23C4DE0",
    x"23C4ACD",
    x"23C47BB",
    x"23C44A9",
    x"23C4198",
    x"23C3E88",
    x"23C3B79",
    x"23C386B",
    x"23C355D",
    x"23C3250",
    x"23C2F44",
    x"23C2C38",
    x"23C292E",
    x"23C2624",
    x"23C231B",
    x"23C2012",
    x"23C1D0B",
    x"23C1A04",
    x"23C16FE",
    x"23C13F8",
    x"23C10F4",
    x"23C0DF0",
    x"23C0AED",
    x"23C07EA",
    x"23C04E9",
    x"23C01E8",
    x"23BFEE8",
    x"23BFBE8",
    x"23BF8EA",
    x"23BF5EC",
    x"23BF2EF",
    x"23BEFF2",
    x"23BECF7",
    x"23BE9FC",
    x"23BE702",
    x"23BE408",
    x"23BE110",
    x"23BDE18",
    x"23BDB21",
    x"23BD82A",
    x"23BD535",
    x"23BD240",
    x"23BCF4C",
    x"23BCC58",
    x"23BC965",
    x"23BC673",
    x"23BC382",
    x"23BC092",
    x"23BBDA2",
    x"23BBAB3",
    x"23BB7C5",
    x"23BB4D7",
    x"23BB1EA",
    x"23BAEFE",
    x"23BAC13",
    x"23BA928",
    x"23BA63E",
    x"23BA355",
    x"23BA06C",
    x"23B9D85",
    x"23B9A9E",
    x"23B97B7",
    x"23B94D2",
    x"23B91ED",
    x"23B8F09",
    x"23B8C25",
    x"23B8943",
    x"23B8661",
    x"23B8380",
    x"23B809F",
    x"23B7DBF",
    x"23B7AE0",
    x"23B7802",
    x"23B7524",
    x"23B7247",
    x"23B6F6B",
    x"23B6C90",
    x"23B69B5",
    x"23B66DB",
    x"23B6401",
    x"23B6129",
    x"23B5E51",
    x"23B5B7A",
    x"23B58A3",
    x"23B55CD",
    x"23B52F8",
    x"23B5024",
    x"23B4D50",
    x"23B4A7D",
    x"23B47AB",
    x"23B44D9",
    x"23B4208",
    x"23B3F38",
    x"23B3C69",
    x"23B399A",
    x"23B36CC",
    x"23B33FF",
    x"23B3132",
    x"23B2E66",
    x"23B2B9B",
    x"23B28D0",
    x"23B2606",
    x"23B233D",
    x"23B2075",
    x"23B1DAD",
    x"23B1AE6",
    x"23B181F",
    x"23B155A",
    x"23B1295",
    x"23B0FD1",
    x"23B0D0D",
    x"23B0A4A",
    x"23B0788",
    x"23B04C6",
    x"23B0205",
    x"23AFF45",
    x"23AFC86",
    x"23AF9C7",
    x"23AF709",
    x"23AF44B",
    x"23AF18F",
    x"23AEED3",
    x"23AEC17",
    x"23AE95D",
    x"23AE6A3",
    x"23AE3E9",
    x"23AE131",
    x"23ADE79",
    x"23ADBC1",
    x"23AD90B",
    x"23AD655",
    x"23AD3A0",
    x"23AD0EB",
    x"23ACE37",
    x"23ACB84",
    x"23AC8D1",
    x"23AC620",
    x"23AC36E",
    x"23AC0BE",
    x"23ABE0E",
    x"23ABB5F",
    x"23AB8B0",
    x"23AB602",
    x"23AB355",
    x"23AB0A9",
    x"23AADFD",
    x"23AAB52",
    x"23AA8A7",
    x"23AA5FD",
    x"23AA354",
    x"23AA0AC",
    x"23A9E04",
    x"23A9B5D",
    x"23A98B6",
    x"23A9610",
    x"23A936B",
    x"23A90C7",
    x"23A8E23",
    x"23A8B80",
    x"23A88DD",
    x"23A863B",
    x"23A839A",
    x"23A80F9",
    x"23A7E5A",
    x"23A7BBA",
    x"23A791C",
    x"23A767E",
    x"23A73E0",
    x"23A7144",
    x"23A6EA8",
    x"23A6C0C",
    x"23A6972",
    x"23A66D8",
    x"23A643E",
    x"23A61A6",
    x"23A5F0D",
    x"23A5C76",
    x"23A59DF",
    x"23A5749",
    x"23A54B4",
    x"23A521F",
    x"23A4F8B",
    x"23A4CF7",
    x"23A4A64",
    x"23A47D2",
    x"23A4540",
    x"23A42AF",
    x"23A401F",
    x"23A3D8F",
    x"23A3B00",
    x"23A3872",
    x"23A35E4",
    x"23A3357",
    x"23A30CA",
    x"23A2E3E",
    x"23A2BB3",
    x"23A2928",
    x"23A269E",
    x"23A2415",
    x"23A218C",
    x"23A1F04",
    x"23A1C7D",
    x"23A19F6",
    x"23A1770",
    x"23A14EA",
    x"23A1265",
    x"23A0FE1",
    x"23A0D5E",
    x"23A0ADA",
    x"23A0858",
    x"23A05D6",
    x"23A0355",
    x"23A00D5",
    x"239FE55",
    x"239FBD5",
    x"239F957",
    x"239F6D9",
    x"239F45B",
    x"239F1DF",
    x"239EF62",
    x"239ECE7",
    x"239EA6C",
    x"239E7F2",
    x"239E578",
    x"239E2FF",
    x"239E087",
    x"239DE0F",
    x"239DB98",
    x"239D921",
    x"239D6AB",
    x"239D436",
    x"239D1C1",
    x"239CF4D",
    x"239CCD9",
    x"239CA66",
    x"239C7F4",
    x"239C582",
    x"239C311",
    x"239C0A1",
    x"239BE31",
    x"239BBC2",
    x"239B953",
    x"239B6E5",
    x"239B478",
    x"239B20B",
    x"239AF9F",
    x"239AD33",
    x"239AAC8",
    x"239A85E",
    x"239A5F4",
    x"239A38B",
    x"239A122",
    x"2399EBA",
    x"2399C53",
    x"23999EC",
    x"2399786",
    x"2399520",
    x"23992BB",
    x"2399057",
    x"2398DF3",
    x"2398B90",
    x"239892D",
    x"23986CB",
    x"239846A",
    x"2398209",
    x"2397FA9",
    x"2397D49",
    x"2397AEA",
    x"239788C",
    x"239762E",
    x"23973D1",
    x"2397174",
    x"2396F18",
    x"2396CBC",
    x"2396A61",
    x"2396807",
    x"23965AD",
    x"2396354",
    x"23960FC",
    x"2395EA4",
    x"2395C4C",
    x"23959F6",
    x"23957A0",
    x"239554A",
    x"23952F5",
    x"23950A0",
    x"2394E4D",
    x"2394BF9",
    x"23949A7",
    x"2394754",
    x"2394503",
    x"23942B2",
    x"2394062",
    x"2393E12",
    x"2393BC3",
    x"2393974",
    x"2393726",
    x"23934D8",
    x"239328B",
    x"239303F",
    x"2392DF3",
    x"2392BA8",
    x"239295D",
    x"2392713",
    x"23924CA",
    x"2392281",
    x"2392039",
    x"2391DF1",
    x"2391BAA",
    x"2391963",
    x"239171D",
    x"23914D7",
    x"2391293",
    x"239104E",
    x"2390E0A",
    x"2390BC7",
    x"2390984",
    x"2390742",
    x"2390501",
    x"23902C0",
    x"239007F",
    x"238FE40",
    x"238FC00",
    x"238F9C2",
    x"238F783",
    x"238F546",
    x"238F309",
    x"238F0CC",
    x"238EE90",
    x"238EC55",
    x"238EA1A",
    x"238E7E0",
    x"238E5A6",
    x"238E36D",
    x"238E135",
    x"238DEFD",
    x"238DCC5",
    x"238DA8E",
    x"238D858",
    x"238D622",
    x"238D3ED",
    x"238D1B8",
    x"238CF84",
    x"238CD50",
    x"238CB1D",
    x"238C8EB",
    x"238C6B9",
    x"238C487",
    x"238C257",
    x"238C026",
    x"238BDF6",
    x"238BBC7",
    x"238B999",
    x"238B76A",
    x"238B53D",
    x"238B310",
    x"238B0E3",
    x"238AEB7",
    x"238AC8C",
    x"238AA61",
    x"238A837",
    x"238A60D",
    x"238A3E4",
    x"238A1BB",
    x"2389F93",
    x"2389D6B",
    x"2389B44",
    x"238991E",
    x"23896F8",
    x"23894D2",
    x"23892AD",
    x"2389089",
    x"2388E65",
    x"2388C42",
    x"2388A1F",
    x"23887FD",
    x"23885DB",
    x"23883BA",
    x"2388199",
    x"2387F79",
    x"2387D59",
    x"2387B3A",
    x"238791C",
    x"23876FE",
    x"23874E0",
    x"23872C3",
    x"23870A7",
    x"2386E8B",
    x"2386C6F",
    x"2386A55",
    x"238683A",
    x"2386620",
    x"2386407",
    x"23861EE",
    x"2385FD6",
    x"2385DBF",
    x"2385BA7",
    x"2385991",
    x"238577B",
    x"2385565",
    x"2385350",
    x"238513B",
    x"2384F27",
    x"2384D14",
    x"2384B01",
    x"23848EE",
    x"23846DC",
    x"23844CB",
    x"23842BA",
    x"23840A9",
    x"2383E9A",
    x"2383C8A",
    x"2383A7B",
    x"238386D",
    x"238365F",
    x"2383452",
    x"2383245",
    x"2383039",
    x"2382E2D",
    x"2382C21",
    x"2382A17",
    x"238280C",
    x"2382603",
    x"23823F9",
    x"23821F1",
    x"2381FE8",
    x"2381DE1",
    x"2381BDA",
    x"23819D3",
    x"23817CD",
    x"23815C7",
    x"23813C2",
    x"23811BD",
    x"2380FB9",
    x"2380DB5",
    x"2380BB2",
    x"23809AF",
    x"23807AD",
    x"23805AB",
    x"23803AA",
    x"23801AA",
    x"237FF53",
    x"237FB54",
    x"237F756",
    x"237F358",
    x"237EF5C",
    x"237EB61",
    x"237E766",
    x"237E36D",
    x"237DF75",
    x"237DB7D",
    x"237D787",
    x"237D392",
    x"237CF9D",
    x"237CBAA",
    x"237C7B7",
    x"237C3C6",
    x"237BFD5",
    x"237BBE6",
    x"237B7F7",
    x"237B40A",
    x"237B01D",
    x"237AC32",
    x"237A847",
    x"237A45E",
    x"237A075",
    x"2379C8E",
    x"23798A7",
    x"23794C1",
    x"23790DD",
    x"2378CF9",
    x"2378916",
    x"2378534",
    x"2378153",
    x"2377D74",
    x"2377995",
    x"23775B7",
    x"23771DA",
    x"2376DFE",
    x"2376A23",
    x"2376649",
    x"2376270",
    x"2375E98",
    x"2375AC0",
    x"23756EA",
    x"2375315",
    x"2374F41",
    x"2374B6D",
    x"237479B",
    x"23743CA",
    x"2373FF9",
    x"2373C2A",
    x"237385B",
    x"237348D",
    x"23730C1",
    x"2372CF5",
    x"237292A",
    x"2372560",
    x"2372198",
    x"2371DD0",
    x"2371A09",
    x"2371643",
    x"237127D",
    x"2370EB9",
    x"2370AF6",
    x"2370734",
    x"2370373",
    x"236FFB2",
    x"236FBF3",
    x"236F834",
    x"236F477",
    x"236F0BA",
    x"236ECFE",
    x"236E943",
    x"236E58A",
    x"236E1D1",
    x"236DE19",
    x"236DA62",
    x"236D6AB",
    x"236D2F6",
    x"236CF42",
    x"236CB8F",
    x"236C7DC",
    x"236C42B",
    x"236C07A",
    x"236BCCA",
    x"236B91C",
    x"236B56E",
    x"236B1C1",
    x"236AE15",
    x"236AA6A",
    x"236A6C0",
    x"236A317",
    x"2369F6E",
    x"2369BC7",
    x"2369820",
    x"236947B",
    x"23690D6",
    x"2368D32",
    x"2368990",
    x"23685EE",
    x"236824D",
    x"2367EAC",
    x"2367B0D",
    x"236776F",
    x"23673D2",
    x"2367035",
    x"2366C99",
    x"23668FF",
    x"2366565",
    x"23661CC",
    x"2365E34",
    x"2365A9D",
    x"2365707",
    x"2365371",
    x"2364FDD",
    x"2364C49",
    x"23648B7",
    x"2364525",
    x"2364194",
    x"2363E04",
    x"2363A75",
    x"23636E7",
    x"236335A",
    x"2362FCD",
    x"2362C42",
    x"23628B7",
    x"236252E",
    x"23621A5",
    x"2361E1D",
    x"2361A96",
    x"236170F",
    x"236138A",
    x"2361006",
    x"2360C82",
    x"23608FF",
    x"236057E",
    x"23601FD",
    x"235FE7D",
    x"235FAFD",
    x"235F77F",
    x"235F402",
    x"235F085",
    x"235ED09",
    x"235E98F",
    x"235E615",
    x"235E29C",
    x"235DF23",
    x"235DBAC",
    x"235D835",
    x"235D4C0",
    x"235D14B",
    x"235CDD7",
    x"235CA64",
    x"235C6F2",
    x"235C381",
    x"235C010",
    x"235BCA1",
    x"235B932",
    x"235B5C4",
    x"235B257",
    x"235AEEB",
    x"235AB80",
    x"235A815",
    x"235A4AC",
    x"235A143",
    x"2359DDB",
    x"2359A74",
    x"235970E",
    x"23593A8",
    x"2359044",
    x"2358CE0",
    x"235897D",
    x"235861B",
    x"23582BA",
    x"2357F5A",
    x"2357BFB",
    x"235789C",
    x"235753E",
    x"23571E2",
    x"2356E85",
    x"2356B2A",
    x"23567D0",
    x"2356476",
    x"235611E",
    x"2355DC6",
    x"2355A6F",
    x"2355719",
    x"23553C3",
    x"235506F",
    x"2354D1B",
    x"23549C8",
    x"2354676",
    x"2354325",
    x"2353FD5",
    x"2353C85",
    x"2353936",
    x"23535E8",
    x"235329B",
    x"2352F4F",
    x"2352C04",
    x"23528B9",
    x"235256F",
    x"2352226",
    x"2351EDE",
    x"2351B97",
    x"2351850",
    x"235150B",
    x"23511C6",
    x"2350E82",
    x"2350B3F",
    x"23507FC",
    x"23504BB",
    x"235017A",
    x"234FE3A",
    x"234FAFB",
    x"234F7BC",
    x"234F47F",
    x"234F142",
    x"234EE06",
    x"234EACB",
    x"234E791",
    x"234E457",
    x"234E11F",
    x"234DDE7",
    x"234DAB0",
    x"234D779",
    x"234D444",
    x"234D10F",
    x"234CDDB",
    x"234CAA8",
    x"234C776",
    x"234C445",
    x"234C114",
    x"234BDE4",
    x"234BAB5",
    x"234B787",
    x"234B459",
    x"234B12D",
    x"234AE01",
    x"234AAD6",
    x"234A7AB",
    x"234A482",
    x"234A159",
    x"2349E31",
    x"2349B0A",
    x"23497E4",
    x"23494BE",
    x"2349199",
    x"2348E75",
    x"2348B52",
    x"2348830",
    x"234850E",
    x"23481ED",
    x"2347ECD",
    x"2347BAE",
    x"234788F",
    x"2347571",
    x"2347254",
    x"2346F38",
    x"2346C1D",
    x"2346902",
    x"23465E8",
    x"23462CF",
    x"2345FB7",
    x"2345C9F",
    x"2345989",
    x"2345673",
    x"234535D",
    x"2345049",
    x"2344D35",
    x"2344A22",
    x"2344710",
    x"23443FF",
    x"23440EE",
    x"2343DDE",
    x"2343ACF",
    x"23437C1",
    x"23434B3",
    x"23431A6",
    x"2342E9A",
    x"2342B8F",
    x"2342885",
    x"234257B",
    x"2342272",
    x"2341F6A",
    x"2341C62",
    x"234195B",
    x"2341656",
    x"2341350",
    x"234104C",
    x"2340D48",
    x"2340A45",
    x"2340743",
    x"2340442",
    x"2340141",
    x"233FE41",
    x"233FB42",
    x"233F843",
    x"233F546",
    x"233F249",
    x"233EF4C",
    x"233EC51",
    x"233E956",
    x"233E65C",
    x"233E363",
    x"233E06B",
    x"233DD73",
    x"233DA7C",
    x"233D786",
    x"233D490",
    x"233D19B",
    x"233CEA7",
    x"233CBB4",
    x"233C8C2",
    x"233C5D0",
    x"233C2DF",
    x"233BFEE",
    x"233BCFF",
    x"233BA10",
    x"233B722",
    x"233B434",
    x"233B148",
    x"233AE5C",
    x"233AB70",
    x"233A886",
    x"233A59C",
    x"233A2B3",
    x"2339FCB",
    x"2339CE3",
    x"23399FC",
    x"2339716",
    x"2339431",
    x"233914C",
    x"2338E68",
    x"2338B85",
    x"23388A2",
    x"23385C1",
    x"23382DF",
    x"2337FFF",
    x"2337D1F",
    x"2337A41",
    x"2337762",
    x"2337485",
    x"23371A8",
    x"2336ECC",
    x"2336BF1",
    x"2336916",
    x"233663C",
    x"2336363",
    x"233608A",
    x"2335DB3",
    x"2335ADC",
    x"2335805",
    x"2335530",
    x"233525B",
    x"2334F86",
    x"2334CB3",
    x"23349E0",
    x"233470E",
    x"233443D",
    x"233416C",
    x"2333E9C",
    x"2333BCC",
    x"23338FE",
    x"2333630",
    x"2333363",
    x"2333096",
    x"2332DCB",
    x"2332AFF",
    x"2332835",
    x"233256B",
    x"23322A2",
    x"2331FDA",
    x"2331D12",
    x"2331A4B",
    x"2331785",
    x"23314C0",
    x"23311FB",
    x"2330F37",
    x"2330C73",
    x"23309B0",
    x"23306EE",
    x"233042D",
    x"233016C",
    x"232FEAC",
    x"232FBED",
    x"232F92E",
    x"232F670",
    x"232F3B3",
    x"232F0F7",
    x"232EE3B",
    x"232EB7F",
    x"232E8C5",
    x"232E60B",
    x"232E352",
    x"232E099",
    x"232DDE2",
    x"232DB2A",
    x"232D874",
    x"232D5BE",
    x"232D309",
    x"232D055",
    x"232CDA1",
    x"232CAEE",
    x"232C83B",
    x"232C58A",
    x"232C2D9",
    x"232C028",
    x"232BD79",
    x"232BACA",
    x"232B81B",
    x"232B56E",
    x"232B2C1",
    x"232B014",
    x"232AD68",
    x"232AABD",
    x"232A813",
    x"232A569",
    x"232A2C0",
    x"232A018",
    x"2329D70",
    x"2329AC9",
    x"2329823",
    x"232957D",
    x"23292D8",
    x"2329034",
    x"2328D90",
    x"2328AED",
    x"232884B",
    x"23285A9",
    x"2328308",
    x"2328067",
    x"2327DC8",
    x"2327B28",
    x"232788A",
    x"23275EC",
    x"232734F",
    x"23270B3",
    x"2326E17",
    x"2326B7C",
    x"23268E1",
    x"2326647",
    x"23263AE",
    x"2326115",
    x"2325E7D",
    x"2325BE6",
    x"232594F",
    x"23256B9",
    x"2325424",
    x"232518F",
    x"2324EFB",
    x"2324C68",
    x"23249D5",
    x"2324743",
    x"23244B1",
    x"2324220",
    x"2323F90",
    x"2323D01",
    x"2323A72",
    x"23237E3",
    x"2323556",
    x"23232C9",
    x"232303C",
    x"2322DB1",
    x"2322B26",
    x"232289B",
    x"2322611",
    x"2322388",
    x"2322100",
    x"2321E78",
    x"2321BF0",
    x"232196A",
    x"23216E4",
    x"232145E",
    x"23211D9",
    x"2320F55",
    x"2320CD2",
    x"2320A4F",
    x"23207CD",
    x"232054B",
    x"23202CA",
    x"232004A",
    x"231FDCA",
    x"231FB4B",
    x"231F8CC",
    x"231F64E",
    x"231F3D1",
    x"231F154",
    x"231EED8",
    x"231EC5D",
    x"231E9E2",
    x"231E768",
    x"231E4EE",
    x"231E276",
    x"231DFFD",
    x"231DD86",
    x"231DB0E",
    x"231D898",
    x"231D622",
    x"231D3AD",
    x"231D138",
    x"231CEC4",
    x"231CC51",
    x"231C9DE",
    x"231C76C",
    x"231C4FA",
    x"231C289",
    x"231C019",
    x"231BDA9",
    x"231BB3A",
    x"231B8CC",
    x"231B65E",
    x"231B3F1",
    x"231B184",
    x"231AF18",
    x"231ACAC",
    x"231AA42",
    x"231A7D7",
    x"231A56E",
    x"231A305",
    x"231A09C",
    x"2319E34",
    x"2319BCD",
    x"2319966",
    x"2319700",
    x"231949B",
    x"2319236",
    x"2318FD2",
    x"2318D6E",
    x"2318B0B",
    x"23188A9",
    x"2318647",
    x"23183E5",
    x"2318185",
    x"2317F25",
    x"2317CC5",
    x"2317A66",
    x"2317808",
    x"23175AA",
    x"231734D",
    x"23170F1",
    x"2316E95",
    x"2316C39",
    x"23169DF",
    x"2316784",
    x"231652B",
    x"23162D2",
    x"2316079",
    x"2315E22",
    x"2315BCA",
    x"2315974",
    x"231571E",
    x"23154C8",
    x"2315273",
    x"231501F",
    x"2314DCB",
    x"2314B78",
    x"2314925",
    x"23146D3",
    x"2314482",
    x"2314231",
    x"2313FE1",
    x"2313D91",
    x"2313B42",
    x"23138F4",
    x"23136A6",
    x"2313458",
    x"231320B",
    x"2312FBF",
    x"2312D74",
    x"2312B29",
    x"23128DE",
    x"2312694",
    x"231244B",
    x"2312202",
    x"2311FBA",
    x"2311D72",
    x"2311B2B",
    x"23118E4",
    x"231169F",
    x"2311459",
    x"2311214",
    x"2310FD0",
    x"2310D8C",
    x"2310B49",
    x"2310907",
    x"23106C5",
    x"2310483",
    x"2310243",
    x"2310002",
    x"230FDC3",
    x"230FB83",
    x"230F945",
    x"230F707",
    x"230F4C9",
    x"230F28C",
    x"230F050",
    x"230EE14",
    x"230EBD9",
    x"230E99E",
    x"230E764",
    x"230E52B",
    x"230E2F2",
    x"230E0B9",
    x"230DE81",
    x"230DC4A",
    x"230DA13",
    x"230D7DD",
    x"230D5A7",
    x"230D372",
    x"230D13D",
    x"230CF09",
    x"230CCD6",
    x"230CAA3",
    x"230C871",
    x"230C63F",
    x"230C40D",
    x"230C1DD",
    x"230BFAD",
    x"230BD7D",
    x"230BB4E",
    x"230B91F",
    x"230B6F1",
    x"230B4C4",
    x"230B297",
    x"230B06A",
    x"230AE3F",
    x"230AC13",
    x"230A9E9",
    x"230A7BE",
    x"230A595",
    x"230A36C",
    x"230A143",
    x"2309F1B",
    x"2309CF3",
    x"2309ACC",
    x"23098A6",
    x"2309680",
    x"230945B",
    x"2309236",
    x"2309012",
    x"2308DEE",
    x"2308BCB",
    x"23089A8",
    x"2308786",
    x"2308564",
    x"2308343",
    x"2308123",
    x"2307F03",
    x"2307CE3",
    x"2307AC4",
    x"23078A6",
    x"2307688",
    x"230746B",
    x"230724E",
    x"2307031",
    x"2306E16",
    x"2306BFA",
    x"23069E0",
    x"23067C5",
    x"23065AC",
    x"2306393",
    x"230617A",
    x"2305F62",
    x"2305D4A",
    x"2305B33",
    x"230591D",
    x"2305707",
    x"23054F1",
    x"23052DC",
    x"23050C8",
    x"2304EB4",
    x"2304CA0",
    x"2304A8D",
    x"230487B",
    x"2304669",
    x"2304458",
    x"2304247",
    x"2304037",
    x"2303E27",
    x"2303C18",
    x"2303A09",
    x"23037FB",
    x"23035ED",
    x"23033E0",
    x"23031D3",
    x"2302FC7",
    x"2302DBB",
    x"2302BB0",
    x"23029A5",
    x"230279B",
    x"2302591",
    x"2302388",
    x"2302180",
    x"2301F77",
    x"2301D70",
    x"2301B69",
    x"2301962",
    x"230175C",
    x"2301556",
    x"2301351",
    x"230114D",
    x"2300F49",
    x"2300D45",
    x"2300B42",
    x"2300940",
    x"230073D",
    x"230053C",
    x"230033B",
    x"230013A",
    x"22FFE75",
    x"22FFA76",
    x"22FF678",
    x"22FF27B",
    x"22FEE7F",
    x"22FEA83",
    x"22FE689",
    x"22FE290",
    x"22FDE98",
    x"22FDAA1",
    x"22FD6AB",
    x"22FD2B5",
    x"22FCEC1",
    x"22FCACE",
    x"22FC6DC",
    x"22FC2EB",
    x"22FBEFA",
    x"22FBB0B",
    x"22FB71D",
    x"22FB330",
    x"22FAF43",
    x"22FAB58",
    x"22FA76E",
    x"22FA384",
    x"22F9F9C",
    x"22F9BB4",
    x"22F97CE",
    x"22F93E9",
    x"22F9004",
    x"22F8C21",
    x"22F883E",
    x"22F845C",
    x"22F807C",
    x"22F7C9C",
    x"22F78BE",
    x"22F74E0",
    x"22F7103",
    x"22F6D27",
    x"22F694D",
    x"22F6573",
    x"22F619A",
    x"22F5DC2",
    x"22F59EB",
    x"22F5615",
    x"22F5240",
    x"22F4E6C",
    x"22F4A99",
    x"22F46C6",
    x"22F42F5",
    x"22F3F25",
    x"22F3B56",
    x"22F3787",
    x"22F33BA",
    x"22F2FED",
    x"22F2C22",
    x"22F2857",
    x"22F248E",
    x"22F20C5",
    x"22F1CFD",
    x"22F1937",
    x"22F1571",
    x"22F11AC",
    x"22F0DE8",
    x"22F0A25",
    x"22F0663",
    x"22F02A2",
    x"22EFEE2",
    x"22EFB22",
    x"22EF764",
    x"22EF3A7",
    x"22EEFEA",
    x"22EEC2F",
    x"22EE874",
    x"22EE4BA",
    x"22EE102",
    x"22EDD4A",
    x"22ED993",
    x"22ED5DD",
    x"22ED228",
    x"22ECE74",
    x"22ECAC1",
    x"22EC70F",
    x"22EC35D",
    x"22EBFAD",
    x"22EBBFE",
    x"22EB84F",
    x"22EB4A1",
    x"22EB0F5",
    x"22EAD49",
    x"22EA99E",
    x"22EA5F4",
    x"22EA24B",
    x"22E9EA3",
    x"22E9AFC",
    x"22E9755",
    x"22E93B0",
    x"22E900C",
    x"22E8C68",
    x"22E88C5",
    x"22E8524",
    x"22E8183",
    x"22E7DE3",
    x"22E7A44",
    x"22E76A6",
    x"22E7309",
    x"22E6F6C",
    x"22E6BD1",
    x"22E6836",
    x"22E649D",
    x"22E6104",
    x"22E5D6C",
    x"22E59D5",
    x"22E563F",
    x"22E52AA",
    x"22E4F16",
    x"22E4B83",
    x"22E47F0",
    x"22E445F",
    x"22E40CE",
    x"22E3D3E",
    x"22E39AF",
    x"22E3621",
    x"22E3294",
    x"22E2F08",
    x"22E2B7D",
    x"22E27F2",
    x"22E2469",
    x"22E20E0",
    x"22E1D58",
    x"22E19D2",
    x"22E164C",
    x"22E12C6",
    x"22E0F42",
    x"22E0BBF",
    x"22E083C",
    x"22E04BB",
    x"22E013A",
    x"22DFDBA",
    x"22DFA3B",
    x"22DF6BD",
    x"22DF340",
    x"22DEFC3",
    x"22DEC48",
    x"22DE8CD",
    x"22DE553",
    x"22DE1DA",
    x"22DDE62",
    x"22DDAEB",
    x"22DD775",
    x"22DD400",
    x"22DD08B",
    x"22DCD17",
    x"22DC9A4",
    x"22DC632",
    x"22DC2C1",
    x"22DBF51",
    x"22DBBE2",
    x"22DB873",
    x"22DB505",
    x"22DB199",
    x"22DAE2D",
    x"22DAAC2",
    x"22DA757",
    x"22DA3EE",
    x"22DA085",
    x"22D9D1E",
    x"22D99B7",
    x"22D9651",
    x"22D92EC",
    x"22D8F87",
    x"22D8C24",
    x"22D88C1",
    x"22D855F",
    x"22D81FF",
    x"22D7E9E",
    x"22D7B3F",
    x"22D77E1",
    x"22D7483",
    x"22D7127",
    x"22D6DCB",
    x"22D6A70",
    x"22D6715",
    x"22D63BC",
    x"22D6064",
    x"22D5D0C",
    x"22D59B5",
    x"22D565F",
    x"22D530A",
    x"22D4FB6",
    x"22D4C62",
    x"22D490F",
    x"22D45BE",
    x"22D426C",
    x"22D3F1C",
    x"22D3BCD",
    x"22D387E",
    x"22D3531",
    x"22D31E4",
    x"22D2E98",
    x"22D2B4C",
    x"22D2802",
    x"22D24B8",
    x"22D2170",
    x"22D1E28",
    x"22D1AE1",
    x"22D179A",
    x"22D1455",
    x"22D1110",
    x"22D0DCC",
    x"22D0A89",
    x"22D0747",
    x"22D0406",
    x"22D00C5",
    x"22CFD85",
    x"22CFA46",
    x"22CF708",
    x"22CF3CB",
    x"22CF08E",
    x"22CED52",
    x"22CEA18",
    x"22CE6DD",
    x"22CE3A4",
    x"22CE06C",
    x"22CDD34",
    x"22CD9FD",
    x"22CD6C7",
    x"22CD392",
    x"22CD05D",
    x"22CCD29",
    x"22CC9F7",
    x"22CC6C4",
    x"22CC393",
    x"22CC063",
    x"22CBD33",
    x"22CBA04",
    x"22CB6D6",
    x"22CB3A9",
    x"22CB07C",
    x"22CAD50",
    x"22CAA25",
    x"22CA6FB",
    x"22CA3D2",
    x"22CA0A9",
    x"22C9D82",
    x"22C9A5B",
    x"22C9734",
    x"22C940F",
    x"22C90EA",
    x"22C8DC7",
    x"22C8AA4",
    x"22C8781",
    x"22C8460",
    x"22C813F",
    x"22C7E1F",
    x"22C7B00",
    x"22C77E2",
    x"22C74C4",
    x"22C71A7",
    x"22C6E8B",
    x"22C6B70",
    x"22C6856",
    x"22C653C",
    x"22C6223",
    x"22C5F0B",
    x"22C5BF3",
    x"22C58DD",
    x"22C55C7",
    x"22C52B2",
    x"22C4F9E",
    x"22C4C8A",
    x"22C4977",
    x"22C4665",
    x"22C4354",
    x"22C4044",
    x"22C3D34",
    x"22C3A25",
    x"22C3717",
    x"22C340A",
    x"22C30FD",
    x"22C2DF1",
    x"22C2AE6",
    x"22C27DC",
    x"22C24D2",
    x"22C21C9",
    x"22C1EC1",
    x"22C1BBA",
    x"22C18B3",
    x"22C15AD",
    x"22C12A8",
    x"22C0FA4",
    x"22C0CA1",
    x"22C099E",
    x"22C069C",
    x"22C039A",
    x"22C009A",
    x"22BFD9A",
    x"22BFA9B",
    x"22BF79D",
    x"22BF49F",
    x"22BF1A3",
    x"22BEEA7",
    x"22BEBAB",
    x"22BE8B1",
    x"22BE5B7",
    x"22BE2BE",
    x"22BDFC6",
    x"22BDCCE",
    x"22BD9D7",
    x"22BD6E1",
    x"22BD3EC",
    x"22BD0F7",
    x"22BCE03",
    x"22BCB10",
    x"22BC81E",
    x"22BC52C",
    x"22BC23B",
    x"22BBF4B",
    x"22BBC5B",
    x"22BB96D",
    x"22BB67F",
    x"22BB391",
    x"22BB0A5",
    x"22BADB9",
    x"22BAACE",
    x"22BA7E4",
    x"22BA4FA",
    x"22BA211",
    x"22B9F29",
    x"22B9C42",
    x"22B995B",
    x"22B9675",
    x"22B9390",
    x"22B90AB",
    x"22B8DC7",
    x"22B8AE4",
    x"22B8802",
    x"22B8520",
    x"22B823F",
    x"22B7F5F",
    x"22B7C80",
    x"22B79A1",
    x"22B76C3",
    x"22B73E6",
    x"22B7109",
    x"22B6E2D",
    x"22B6B52",
    x"22B6877",
    x"22B659E",
    x"22B62C5",
    x"22B5FEC",
    x"22B5D15",
    x"22B5A3E",
    x"22B5767",
    x"22B5492",
    x"22B51BD",
    x"22B4EE9",
    x"22B4C16",
    x"22B4943",
    x"22B4671",
    x"22B43A0",
    x"22B40CF",
    x"22B3DFF",
    x"22B3B30",
    x"22B3862",
    x"22B3594",
    x"22B32C7",
    x"22B2FFB",
    x"22B2D2F",
    x"22B2A64",
    x"22B279A",
    x"22B24D0",
    x"22B2207",
    x"22B1F3F",
    x"22B1C78",
    x"22B19B1",
    x"22B16EB",
    x"22B1426",
    x"22B1161",
    x"22B0E9D",
    x"22B0BDA",
    x"22B0917",
    x"22B0655",
    x"22B0394",
    x"22B00D3",
    x"22AFE13",
    x"22AFB54",
    x"22AF896",
    x"22AF5D8",
    x"22AF31B",
    x"22AF05E",
    x"22AEDA3",
    x"22AEAE8",
    x"22AE82D",
    x"22AE573",
    x"22AE2BA",
    x"22AE002",
    x"22ADD4A",
    x"22ADA93",
    x"22AD7DD",
    x"22AD528",
    x"22AD273",
    x"22ACFBE",
    x"22ACD0B",
    x"22ACA58",
    x"22AC7A6",
    x"22AC4F4",
    x"22AC243",
    x"22ABF93",
    x"22ABCE3",
    x"22ABA34",
    x"22AB786",
    x"22AB4D9",
    x"22AB22C",
    x"22AAF80",
    x"22AACD4",
    x"22AAA29",
    x"22AA77F",
    x"22AA4D5",
    x"22AA22C",
    x"22A9F84",
    x"22A9CDD",
    x"22A9A36",
    x"22A9790",
    x"22A94EA",
    x"22A9245",
    x"22A8FA1",
    x"22A8CFD",
    x"22A8A5A",
    x"22A87B8",
    x"22A8517",
    x"22A8276",
    x"22A7FD5",
    x"22A7D36",
    x"22A7A97",
    x"22A77F8",
    x"22A755B",
    x"22A72BE",
    x"22A7021",
    x"22A6D86",
    x"22A6AEB",
    x"22A6850",
    x"22A65B6",
    x"22A631D",
    x"22A6085",
    x"22A5DED",
    x"22A5B56",
    x"22A58BF",
    x"22A562A",
    x"22A5394",
    x"22A5100",
    x"22A4E6C",
    x"22A4BD9",
    x"22A4946",
    x"22A46B4",
    x"22A4423",
    x"22A4192",
    x"22A3F02",
    x"22A3C72",
    x"22A39E4",
    x"22A3755",
    x"22A34C8",
    x"22A323B",
    x"22A2FAF",
    x"22A2D23",
    x"22A2A98",
    x"22A280E",
    x"22A2584",
    x"22A22FB",
    x"22A2073",
    x"22A1DEB",
    x"22A1B64",
    x"22A18DD",
    x"22A1657",
    x"22A13D2",
    x"22A114D",
    x"22A0EC9",
    x"22A0C46",
    x"22A09C3",
    x"22A0741",
    x"22A04C0",
    x"22A023F",
    x"229FFBE",
    x"229FD3F",
    x"229FAC0",
    x"229F841",
    x"229F5C4",
    x"229F347",
    x"229F0CA",
    x"229EE4E",
    x"229EBD3",
    x"229E958",
    x"229E6DE",
    x"229E465",
    x"229E1EC",
    x"229DF74",
    x"229DCFC",
    x"229DA85",
    x"229D80F",
    x"229D599",
    x"229D324",
    x"229D0B0",
    x"229CE3C",
    x"229CBC9",
    x"229C956",
    x"229C6E4",
    x"229C473",
    x"229C202",
    x"229BF92",
    x"229BD22",
    x"229BAB3",
    x"229B845",
    x"229B5D7",
    x"229B36A",
    x"229B0FD",
    x"229AE91",
    x"229AC26",
    x"229A9BB",
    x"229A751",
    x"229A4E7",
    x"229A27F",
    x"229A016",
    x"2299DAF",
    x"2299B47",
    x"22998E1",
    x"229967B",
    x"2299416",
    x"22991B1",
    x"2298F4D",
    x"2298CE9",
    x"2298A86",
    x"2298824",
    x"22985C2",
    x"2298361",
    x"2298101",
    x"2297EA1",
    x"2297C41",
    x"22979E2",
    x"2297784",
    x"2297527",
    x"22972CA",
    x"229706D",
    x"2296E12",
    x"2296BB6",
    x"229695C",
    x"2296702",
    x"22964A8",
    x"229624F",
    x"2295FF7",
    x"2295D9F",
    x"2295B48",
    x"22958F2",
    x"229569C",
    x"2295446",
    x"22951F2",
    x"2294F9D",
    x"2294D4A",
    x"2294AF7",
    x"22948A4",
    x"2294652",
    x"2294401",
    x"22941B0",
    x"2293F60",
    x"2293D11",
    x"2293AC2",
    x"2293873",
    x"2293626",
    x"22933D8",
    x"229318C",
    x"2292F40",
    x"2292CF4",
    x"2292AA9",
    x"229285F",
    x"2292615",
    x"22923CC",
    x"2292183",
    x"2291F3B",
    x"2291CF3",
    x"2291AAC",
    x"2291866",
    x"2291620",
    x"22913DB",
    x"2291196",
    x"2290F52",
    x"2290D0F",
    x"2290ACC",
    x"2290889",
    x"2290647",
    x"2290406",
    x"22901C5",
    x"228FF85",
    x"228FD46",
    x"228FB07",
    x"228F8C8",
    x"228F68A",
    x"228F44D",
    x"228F210",
    x"228EFD4",
    x"228ED98",
    x"228EB5D",
    x"228E922",
    x"228E6E8",
    x"228E4AF",
    x"228E276",
    x"228E03E",
    x"228DE06",
    x"228DBCF",
    x"228D998",
    x"228D762",
    x"228D52C",
    x"228D2F7",
    x"228D0C3",
    x"228CE8F",
    x"228CC5C",
    x"228CA29",
    x"228C7F6",
    x"228C5C5",
    x"228C394",
    x"228C163",
    x"228BF33",
    x"228BD03",
    x"228BAD4",
    x"228B8A6",
    x"228B678",
    x"228B44B",
    x"228B21E",
    x"228AFF2",
    x"228ADC6",
    x"228AB9B",
    x"228A970",
    x"228A746",
    x"228A51C",
    x"228A2F3",
    x"228A0CB",
    x"2289EA3",
    x"2289C7C",
    x"2289A55",
    x"228982F",
    x"2289609",
    x"22893E4",
    x"22891BF",
    x"2288F9B",
    x"2288D77",
    x"2288B54",
    x"2288931",
    x"228870F",
    x"22884EE",
    x"22882CD",
    x"22880AC",
    x"2287E8D",
    x"2287C6D",
    x"2287A4E",
    x"2287830",
    x"2287612",
    x"22873F5",
    x"22871D8",
    x"2286FBC",
    x"2286DA0",
    x"2286B85",
    x"228696B",
    x"2286750",
    x"2286537",
    x"228631E",
    x"2286105",
    x"2285EED",
    x"2285CD6",
    x"2285ABF",
    x"22858A9",
    x"2285693",
    x"228547D",
    x"2285268",
    x"2285054",
    x"2284E40",
    x"2284C2D",
    x"2284A1A",
    x"2284808",
    x"22845F6",
    x"22843E5",
    x"22841D4",
    x"2283FC4",
    x"2283DB4",
    x"2283BA5",
    x"2283996",
    x"2283788",
    x"228357B",
    x"228336E",
    x"2283161",
    x"2282F55",
    x"2282D49",
    x"2282B3E",
    x"2282934",
    x"228272A",
    x"2282520",
    x"2282317",
    x"228210F",
    x"2281F07",
    x"2281CFF",
    x"2281AF8",
    x"22818F2",
    x"22816EC",
    x"22814E6",
    x"22812E1",
    x"22810DD",
    x"2280ED9",
    x"2280CD5",
    x"2280AD2",
    x"22808D0",
    x"22806CE",
    x"22804CC",
    x"22802CB",
    x"22800CB",
    x"227FD97",
    x"227F998",
    x"227F59A",
    x"227F19D",
    x"227EDA1",
    x"227E9A6",
    x"227E5AC",
    x"227E1B3",
    x"227DDBB",
    x"227D9C4",
    x"227D5CE",
    x"227D1D9",
    x"227CDE6",
    x"227C9F3",
    x"227C601",
    x"227C210",
    x"227BE1F",
    x"227BA30",
    x"227B642",
    x"227B255",
    x"227AE69",
    x"227AA7E",
    x"227A694",
    x"227A2AB",
    x"2279EC3",
    x"2279ADB",
    x"22796F5",
    x"2279310",
    x"2278F2C",
    x"2278B48",
    x"2278766",
    x"2278385",
    x"2277FA4",
    x"2277BC5",
    x"22777E6",
    x"2277409",
    x"227702C",
    x"2276C51",
    x"2276876",
    x"227649D",
    x"22760C4",
    x"2275CEC",
    x"2275915",
    x"2275540",
    x"227516B",
    x"2274D97",
    x"22749C4",
    x"22745F2",
    x"2274221",
    x"2273E51",
    x"2273A82",
    x"22736B4",
    x"22732E7",
    x"2272F1A",
    x"2272B4F",
    x"2272785",
    x"22723BB",
    x"2271FF3",
    x"2271C2B",
    x"2271865",
    x"227149F",
    x"22710DA",
    x"2270D17",
    x"2270954",
    x"2270592",
    x"22701D1",
    x"226FE11",
    x"226FA52",
    x"226F694",
    x"226F2D7",
    x"226EF1A",
    x"226EB5F",
    x"226E7A5",
    x"226E3EB",
    x"226E033",
    x"226DC7B",
    x"226D8C5",
    x"226D50F",
    x"226D15A",
    x"226CDA6",
    x"226C9F3",
    x"226C641",
    x"226C290",
    x"226BEE0",
    x"226BB31",
    x"226B782",
    x"226B3D5",
    x"226B028",
    x"226AC7D",
    x"226A8D2",
    x"226A528",
    x"226A180",
    x"2269DD8",
    x"2269A31",
    x"226968B",
    x"22692E5",
    x"2268F41",
    x"2268B9E",
    x"22687FB",
    x"226845A",
    x"22680B9",
    x"2267D19",
    x"226797B",
    x"22675DD",
    x"2267240",
    x"2266EA4",
    x"2266B08",
    x"226676E",
    x"22663D5",
    x"226603C",
    x"2265CA4",
    x"226590E",
    x"2265578",
    x"22651E3",
    x"2264E4F",
    x"2264ABC",
    x"226472A",
    x"2264398",
    x"2264008",
    x"2263C78",
    x"22638EA",
    x"226355C",
    x"22631CF",
    x"2262E43",
    x"2262AB8",
    x"226272E",
    x"22623A4",
    x"226201C",
    x"2261C94",
    x"226190D",
    x"2261588",
    x"2261203",
    x"2260E7F",
    x"2260AFB",
    x"2260779",
    x"22603F8",
    x"2260077",
    x"225FCF7",
    x"225F979",
    x"225F5FB",
    x"225F27E",
    x"225EF01",
    x"225EB86",
    x"225E80C",
    x"225E492",
    x"225E119",
    x"225DDA2",
    x"225DA2B",
    x"225D6B5",
    x"225D33F",
    x"225CFCB",
    x"225CC57",
    x"225C8E5",
    x"225C573",
    x"225C202",
    x"225BE92",
    x"225BB23",
    x"225B7B4",
    x"225B447",
    x"225B0DA",
    x"225AD6E",
    x"225AA03",
    x"225A699",
    x"225A330",
    x"2259FC8",
    x"2259C60",
    x"22598FA",
    x"2259594",
    x"225922F",
    x"2258ECB",
    x"2258B67",
    x"2258805",
    x"22584A3",
    x"2258143",
    x"2257DE3",
    x"2257A84",
    x"2257726",
    x"22573C8",
    x"225706C",
    x"2256D10",
    x"22569B5",
    x"225665B",
    x"2256302",
    x"2255FAA",
    x"2255C52",
    x"22558FB",
    x"22555A6",
    x"2255251",
    x"2254EFC",
    x"2254BA9",
    x"2254857",
    x"2254505",
    x"22541B4",
    x"2253E64",
    x"2253B15",
    x"22537C7",
    x"2253479",
    x"225312C",
    x"2252DE0",
    x"2252A95",
    x"225274B",
    x"2252402",
    x"22520B9",
    x"2251D71",
    x"2251A2A",
    x"22516E4",
    x"225139F",
    x"225105A",
    x"2250D17",
    x"22509D4",
    x"2250692",
    x"2250351",
    x"2250010",
    x"224FCD1",
    x"224F992",
    x"224F654",
    x"224F317",
    x"224EFDA",
    x"224EC9F",
    x"224E964",
    x"224E62A",
    x"224E2F1",
    x"224DFB9",
    x"224DC81",
    x"224D94A",
    x"224D614",
    x"224D2DF",
    x"224CFAB",
    x"224CC77",
    x"224C945",
    x"224C613",
    x"224C2E2",
    x"224BFB1",
    x"224BC82",
    x"224B953",
    x"224B625",
    x"224B2F8",
    x"224AFCC",
    x"224ACA0",
    x"224A975",
    x"224A64B",
    x"224A322",
    x"2249FFA",
    x"2249CD2",
    x"22499AB",
    x"2249685",
    x"2249360",
    x"224903C",
    x"2248D18",
    x"22489F5",
    x"22486D3",
    x"22483B2",
    x"2248091",
    x"2247D71",
    x"2247A52",
    x"2247734",
    x"2247417",
    x"22470FA",
    x"2246DDE",
    x"2246AC3",
    x"22467A9",
    x"224648F",
    x"2246177",
    x"2245E5F",
    x"2245B48",
    x"2245831",
    x"224551B",
    x"2245207",
    x"2244EF2",
    x"2244BDF",
    x"22448CC",
    x"22445BB",
    x"22442AA",
    x"2243F99",
    x"2243C8A",
    x"224397B",
    x"224366D",
    x"2243360",
    x"2243053",
    x"2242D48",
    x"2242A3D",
    x"2242733",
    x"2242429",
    x"2242120",
    x"2241E19",
    x"2241B11",
    x"224180B",
    x"2241505",
    x"2241201",
    x"2240EFC",
    x"2240BF9",
    x"22408F6",
    x"22405F5",
    x"22402F3",
    x"223FFF3",
    x"223FCF3",
    x"223F9F5",
    x"223F6F6",
    x"223F3F9",
    x"223F0FD",
    x"223EE01",
    x"223EB06",
    x"223E80B",
    x"223E511",
    x"223E219",
    x"223DF20",
    x"223DC29",
    x"223D932",
    x"223D63C",
    x"223D347",
    x"223D053",
    x"223CD5F",
    x"223CA6C",
    x"223C77A",
    x"223C488",
    x"223C198",
    x"223BEA8",
    x"223BBB8",
    x"223B8CA",
    x"223B5DC",
    x"223B2EF",
    x"223B002",
    x"223AD17",
    x"223AA2C",
    x"223A742",
    x"223A458",
    x"223A16F",
    x"2239E88",
    x"2239BA0",
    x"22398BA",
    x"22395D4",
    x"22392EF",
    x"223900A",
    x"2238D27",
    x"2238A44",
    x"2238762",
    x"2238480",
    x"223819F",
    x"2237EBF",
    x"2237BE0",
    x"2237901",
    x"2237623",
    x"2237346",
    x"223706A",
    x"2236D8E",
    x"2236AB3",
    x"22367D9",
    x"22364FF",
    x"2236226",
    x"2235F4E",
    x"2235C77",
    x"22359A0",
    x"22356CA",
    x"22353F4",
    x"2235120",
    x"2234E4C",
    x"2234B79",
    x"22348A6",
    x"22345D4",
    x"2234303",
    x"2234033",
    x"2233D63",
    x"2233A94",
    x"22337C6",
    x"22334F8",
    x"223322B",
    x"2232F5F",
    x"2232C94",
    x"22329C9",
    x"22326FF",
    x"2232435",
    x"223216D",
    x"2231EA5",
    x"2231BDD",
    x"2231917",
    x"2231651",
    x"223138C",
    x"22310C7",
    x"2230E03",
    x"2230B40",
    x"223087E",
    x"22305BC",
    x"22302FB",
    x"223003A",
    x"222FD7B",
    x"222FABC",
    x"222F7FD",
    x"222F540",
    x"222F283",
    x"222EFC6",
    x"222ED0B",
    x"222EA50",
    x"222E796",
    x"222E4DC",
    x"222E223",
    x"222DF6B",
    x"222DCB3",
    x"222D9FD",
    x"222D746",
    x"222D491",
    x"222D1DC",
    x"222CF28",
    x"222CC75",
    x"222C9C2",
    x"222C710",
    x"222C45E",
    x"222C1AD",
    x"222BEFD",
    x"222BC4E",
    x"222B99F",
    x"222B6F1",
    x"222B444",
    x"222B197",
    x"222AEEB",
    x"222AC40",
    x"222A995",
    x"222A6EB",
    x"222A441",
    x"222A199",
    x"2229EF1",
    x"2229C49",
    x"22299A2",
    x"22296FC",
    x"2229457",
    x"22291B2",
    x"2228F0E",
    x"2228C6B",
    x"22289C8",
    x"2228726",
    x"2228484",
    x"22281E3",
    x"2227F43",
    x"2227CA4",
    x"2227A05",
    x"2227767",
    x"22274C9",
    x"222722C",
    x"2226F90",
    x"2226CF5",
    x"2226A5A",
    x"22267C0",
    x"2226526",
    x"222628D",
    x"2225FF5",
    x"2225D5D",
    x"2225AC6",
    x"2225830",
    x"222559A",
    x"2225305",
    x"2225070",
    x"2224DDD",
    x"2224B49",
    x"22248B7",
    x"2224625",
    x"2224394",
    x"2224103",
    x"2223E73",
    x"2223BE4",
    x"2223955",
    x"22236C7",
    x"222343A",
    x"22231AD",
    x"2222F21",
    x"2222C96",
    x"2222A0B",
    x"2222781",
    x"22224F7",
    x"222226E",
    x"2221FE6",
    x"2221D5E",
    x"2221AD7",
    x"2221851",
    x"22215CB",
    x"2221346",
    x"22210C1",
    x"2220E3E",
    x"2220BBA",
    x"2220938",
    x"22206B6",
    x"2220434",
    x"22201B4",
    x"221FF33",
    x"221FCB4",
    x"221FA35",
    x"221F7B7",
    x"221F539",
    x"221F2BC",
    x"221F040",
    x"221EDC4",
    x"221EB49",
    x"221E8CE",
    x"221E655",
    x"221E3DB",
    x"221E163",
    x"221DEEB",
    x"221DC73",
    x"221D9FC",
    x"221D786",
    x"221D511",
    x"221D29C",
    x"221D027",
    x"221CDB4",
    x"221CB40",
    x"221C8CE",
    x"221C65C",
    x"221C3EB",
    x"221C17A",
    x"221BF0A",
    x"221BC9B",
    x"221BA2C",
    x"221B7BD",
    x"221B550",
    x"221B2E3",
    x"221B076",
    x"221AE0B",
    x"221AB9F",
    x"221A935",
    x"221A6CB",
    x"221A461",
    x"221A1F9",
    x"2219F90",
    x"2219D29",
    x"2219AC2",
    x"221985B",
    x"22195F6",
    x"2219390",
    x"221912C",
    x"2218EC8",
    x"2218C64",
    x"2218A02",
    x"221879F",
    x"221853E",
    x"22182DD",
    x"221807C",
    x"2217E1D",
    x"2217BBD",
    x"221795F",
    x"2217701",
    x"22174A3",
    x"2217246",
    x"2216FEA",
    x"2216D8E",
    x"2216B33",
    x"22168D9",
    x"221667F",
    x"2216426",
    x"22161CD",
    x"2215F75",
    x"2215D1D",
    x"2215AC6",
    x"2215870",
    x"221561A",
    x"22153C5",
    x"2215170",
    x"2214F1C",
    x"2214CC8",
    x"2214A76",
    x"2214823",
    x"22145D1",
    x"2214380",
    x"2214130",
    x"2213EE0",
    x"2213C90",
    x"2213A41",
    x"22137F3",
    x"22135A5",
    x"2213358",
    x"221310C",
    x"2212EC0",
    x"2212C74",
    x"2212A2A",
    x"22127DF",
    x"2212596",
    x"221234D",
    x"2212104",
    x"2211EBC",
    x"2211C75",
    x"2211A2E",
    x"22117E8",
    x"22115A2",
    x"221135D",
    x"2211118",
    x"2210ED4",
    x"2210C91",
    x"2210A4E",
    x"221080C",
    x"22105CA",
    x"2210389",
    x"2210148",
    x"220FF08",
    x"220FCC9",
    x"220FA8A",
    x"220F84B",
    x"220F60D",
    x"220F3D0",
    x"220F194",
    x"220EF57",
    x"220ED1C",
    x"220EAE1",
    x"220E8A6",
    x"220E66D",
    x"220E433",
    x"220E1FA",
    x"220DFC2",
    x"220DD8B",
    x"220DB54",
    x"220D91D",
    x"220D6E7",
    x"220D4B1",
    x"220D27D",
    x"220D048",
    x"220CE14",
    x"220CBE1",
    x"220C9AF",
    x"220C77C",
    x"220C54B",
    x"220C31A",
    x"220C0E9",
    x"220BEB9",
    x"220BC8A",
    x"220BA5B",
    x"220B82D",
    x"220B5FF",
    x"220B3D2",
    x"220B1A5",
    x"220AF79",
    x"220AD4D",
    x"220AB22",
    x"220A8F8",
    x"220A6CE",
    x"220A4A4",
    x"220A27B",
    x"220A053",
    x"2209E2B",
    x"2209C04",
    x"22099DD",
    x"22097B7",
    x"2209591",
    x"220936C",
    x"2209148",
    x"2208F24",
    x"2208D00",
    x"2208ADD",
    x"22088BB",
    x"2208699",
    x"2208477",
    x"2208256",
    x"2208036",
    x"2207E16",
    x"2207BF7",
    x"22079D8",
    x"22077BA",
    x"220759D",
    x"220737F",
    x"2207163",
    x"2206F47",
    x"2206D2B",
    x"2206B10",
    x"22068F6",
    x"22066DC",
    x"22064C2",
    x"22062A9",
    x"2206091",
    x"2205E79",
    x"2205C62",
    x"2205A4B",
    x"2205834",
    x"220561F",
    x"2205409",
    x"22051F5",
    x"2204FE0",
    x"2204DCD",
    x"2204BBA",
    x"22049A7",
    x"2204795",
    x"2204583",
    x"2204372",
    x"2204161",
    x"2203F51",
    x"2203D42",
    x"2203B33",
    x"2203924",
    x"2203716",
    x"2203509",
    x"22032FC",
    x"22030EF",
    x"2202EE3",
    x"2202CD8",
    x"2202ACD",
    x"22028C2",
    x"22026B8",
    x"22024AF",
    x"22022A6",
    x"220209E",
    x"2201E96",
    x"2201C8E",
    x"2201A87",
    x"2201881",
    x"220167B",
    x"2201476",
    x"2201271",
    x"220106C",
    x"2200E69",
    x"2200C65",
    x"2200A62",
    x"2200860",
    x"220065E",
    x"220045D",
    x"220025C",
    x"220005C",
    x"21FFCB8",
    x"21FF8BA",
    x"21FF4BC",
    x"21FF0BF",
    x"21FECC4",
    x"21FE8C9",
    x"21FE4CF",
    x"21FE0D6",
    x"21FDCDF",
    x"21FD8E8",
    x"21FD4F2",
    x"21FD0FE",
    x"21FCD0A",
    x"21FC917",
    x"21FC525",
    x"21FC134",
    x"21FBD45",
    x"21FB956",
    x"21FB568",
    x"21FB17B",
    x"21FAD8F",
    x"21FA9A4",
    x"21FA5BA",
    x"21FA1D1",
    x"21F9DE9",
    x"21F9A02",
    x"21F961C",
    x"21F9237",
    x"21F8E53",
    x"21F8A70",
    x"21F868E",
    x"21F82AD",
    x"21F7ECD",
    x"21F7AEE",
    x"21F770F",
    x"21F7332",
    x"21F6F56",
    x"21F6B7A",
    x"21F67A0",
    x"21F63C7",
    x"21F5FEE",
    x"21F5C17",
    x"21F5840",
    x"21F546A",
    x"21F5096",
    x"21F4CC2",
    x"21F48EF",
    x"21F451E",
    x"21F414D",
    x"21F3D7D",
    x"21F39AE",
    x"21F35E0",
    x"21F3213",
    x"21F2E47",
    x"21F2A7C",
    x"21F26B2",
    x"21F22E9",
    x"21F1F20",
    x"21F1B59",
    x"21F1793",
    x"21F13CD",
    x"21F1009",
    x"21F0C45",
    x"21F0883",
    x"21F04C1",
    x"21F0100",
    x"21EFD41",
    x"21EF982",
    x"21EF5C4",
    x"21EF207",
    x"21EEE4B",
    x"21EEA90",
    x"21EE6D6",
    x"21EE31C",
    x"21EDF64",
    x"21EDBAD",
    x"21ED7F6",
    x"21ED441",
    x"21ED08C",
    x"21ECCD8",
    x"21EC926",
    x"21EC574",
    x"21EC1C3",
    x"21EBE13",
    x"21EBA64",
    x"21EB6B6",
    x"21EB308",
    x"21EAF5C",
    x"21EABB1",
    x"21EA806",
    x"21EA45D",
    x"21EA0B4",
    x"21E9D0C",
    x"21E9966",
    x"21E95C0",
    x"21E921B",
    x"21E8E77",
    x"21E8AD4",
    x"21E8731",
    x"21E8390",
    x"21E7FEF",
    x"21E7C50",
    x"21E78B1",
    x"21E7514",
    x"21E7177",
    x"21E6DDB",
    x"21E6A40",
    x"21E66A6",
    x"21E630D",
    x"21E5F74",
    x"21E5BDD",
    x"21E5846",
    x"21E54B1",
    x"21E511C",
    x"21E4D88",
    x"21E49F5",
    x"21E4663",
    x"21E42D2",
    x"21E3F42",
    x"21E3BB2",
    x"21E3824",
    x"21E3496",
    x"21E310A",
    x"21E2D7E",
    x"21E29F3",
    x"21E2669",
    x"21E22E0",
    x"21E1F57",
    x"21E1BD0",
    x"21E1849",
    x"21E14C4",
    x"21E113F",
    x"21E0DBB",
    x"21E0A38",
    x"21E06B6",
    x"21E0335",
    x"21DFFB4",
    x"21DFC35",
    x"21DF8B6",
    x"21DF539",
    x"21DF1BC",
    x"21DEE40",
    x"21DEAC5",
    x"21DE74A",
    x"21DE3D1",
    x"21DE058",
    x"21DDCE1",
    x"21DD96A",
    x"21DD5F4",
    x"21DD27F",
    x"21DCF0B",
    x"21DCB98",
    x"21DC825",
    x"21DC4B3",
    x"21DC143",
    x"21DBDD3",
    x"21DBA64",
    x"21DB6F6",
    x"21DB388",
    x"21DB01C",
    x"21DACB0",
    x"21DA945",
    x"21DA5DC",
    x"21DA273",
    x"21D9F0A",
    x"21D9BA3",
    x"21D983D",
    x"21D94D7",
    x"21D9172",
    x"21D8E0E",
    x"21D8AAB",
    x"21D8749",
    x"21D83E7",
    x"21D8087",
    x"21D7D27",
    x"21D79C8",
    x"21D766A",
    x"21D730D",
    x"21D6FB1",
    x"21D6C55",
    x"21D68FB",
    x"21D65A1",
    x"21D6248",
    x"21D5EF0",
    x"21D5B98",
    x"21D5842",
    x"21D54EC",
    x"21D5197",
    x"21D4E43",
    x"21D4AF0",
    x"21D479E",
    x"21D444C",
    x"21D40FC",
    x"21D3DAC",
    x"21D3A5D",
    x"21D370F",
    x"21D33C1",
    x"21D3075",
    x"21D2D29",
    x"21D29DE",
    x"21D2694",
    x"21D234B",
    x"21D2003",
    x"21D1CBB",
    x"21D1974",
    x"21D162E",
    x"21D12E9",
    x"21D0FA5",
    x"21D0C61",
    x"21D091F",
    x"21D05DD",
    x"21D029C",
    x"21CFF5B",
    x"21CFC1C",
    x"21CF8DD",
    x"21CF5A0",
    x"21CF263",
    x"21CEF26",
    x"21CEBEB",
    x"21CE8B0",
    x"21CE577",
    x"21CE23E",
    x"21CDF06",
    x"21CDBCE",
    x"21CD898",
    x"21CD562",
    x"21CD22D",
    x"21CCEF9",
    x"21CCBC5",
    x"21CC893",
    x"21CC561",
    x"21CC230",
    x"21CBF00",
    x"21CBBD1",
    x"21CB8A2",
    x"21CB574",
    x"21CB247",
    x"21CAF1B",
    x"21CABF0",
    x"21CA8C5",
    x"21CA59B",
    x"21CA272",
    x"21C9F4A",
    x"21C9C23",
    x"21C98FC",
    x"21C95D6",
    x"21C92B1",
    x"21C8F8D",
    x"21C8C6A",
    x"21C8947",
    x"21C8625",
    x"21C8304",
    x"21C7FE3",
    x"21C7CC4",
    x"21C79A5",
    x"21C7687",
    x"21C736A",
    x"21C704D",
    x"21C6D32",
    x"21C6A17",
    x"21C66FD",
    x"21C63E3",
    x"21C60CB",
    x"21C5DB3",
    x"21C5A9C",
    x"21C5785",
    x"21C5470",
    x"21C515B",
    x"21C4E47",
    x"21C4B34",
    x"21C4822",
    x"21C4510",
    x"21C41FF",
    x"21C3EEF",
    x"21C3BE0",
    x"21C38D1",
    x"21C35C3",
    x"21C32B6",
    x"21C2FAA",
    x"21C2C9E",
    x"21C2994",
    x"21C268A",
    x"21C2380",
    x"21C2078",
    x"21C1D70",
    x"21C1A69",
    x"21C1763",
    x"21C145D",
    x"21C1159",
    x"21C0E55",
    x"21C0B52",
    x"21C084F",
    x"21C054D",
    x"21C024C",
    x"21BFF4C",
    x"21BFC4D",
    x"21BF94E",
    x"21BF650",
    x"21BF353",
    x"21BF056",
    x"21BED5B",
    x"21BEA60",
    x"21BE766",
    x"21BE46C",
    x"21BE173",
    x"21BDE7B",
    x"21BDB84",
    x"21BD88E",
    x"21BD598",
    x"21BD2A3",
    x"21BCFAF",
    x"21BCCBB",
    x"21BC9C8",
    x"21BC6D6",
    x"21BC3E5",
    x"21BC0F4",
    x"21BBE04",
    x"21BBB15",
    x"21BB827",
    x"21BB539",
    x"21BB24C",
    x"21BAF60",
    x"21BAC74",
    x"21BA98A",
    x"21BA6A0",
    x"21BA3B6",
    x"21BA0CE",
    x"21B9DE6",
    x"21B9AFF",
    x"21B9818",
    x"21B9533",
    x"21B924E",
    x"21B8F6A",
    x"21B8C86",
    x"21B89A3",
    x"21B86C1",
    x"21B83E0",
    x"21B80FF",
    x"21B7E1F",
    x"21B7B40",
    x"21B7862",
    x"21B7584",
    x"21B72A7",
    x"21B6FCB",
    x"21B6CEF",
    x"21B6A14",
    x"21B673A",
    x"21B6461",
    x"21B6188",
    x"21B5EB0",
    x"21B5BD9",
    x"21B5902",
    x"21B562C",
    x"21B5357",
    x"21B5082",
    x"21B4DAF",
    x"21B4ADC",
    x"21B4809",
    x"21B4538",
    x"21B4267",
    x"21B3F96",
    x"21B3CC7",
    x"21B39F8",
    x"21B372A",
    x"21B345C",
    x"21B3190",
    x"21B2EC4",
    x"21B2BF8",
    x"21B292E",
    x"21B2664",
    x"21B239A",
    x"21B20D2",
    x"21B1E0A",
    x"21B1B43",
    x"21B187C",
    x"21B15B7",
    x"21B12F2",
    x"21B102D",
    x"21B0D69",
    x"21B0AA6",
    x"21B07E4",
    x"21B0523",
    x"21B0262",
    x"21AFFA1",
    x"21AFCE2",
    x"21AFA23",
    x"21AF765",
    x"21AF4A7",
    x"21AF1EA",
    x"21AEF2E",
    x"21AEC73",
    x"21AE9B8",
    x"21AE6FE",
    x"21AE444",
    x"21AE18C",
    x"21ADED4",
    x"21ADC1C",
    x"21AD966",
    x"21AD6B0",
    x"21AD3FA",
    x"21AD146",
    x"21ACE92",
    x"21ACBDE",
    x"21AC92C",
    x"21AC67A",
    x"21AC3C9",
    x"21AC118",
    x"21ABE68",
    x"21ABBB9",
    x"21AB90A",
    x"21AB65C",
    x"21AB3AF",
    x"21AB102",
    x"21AAE56",
    x"21AABAB",
    x"21AA901",
    x"21AA657",
    x"21AA3AD",
    x"21AA105",
    x"21A9E5D",
    x"21A9BB6",
    x"21A990F",
    x"21A9669",
    x"21A93C4",
    x"21A911F",
    x"21A8E7B",
    x"21A8BD8",
    x"21A8935",
    x"21A8693",
    x"21A83F2",
    x"21A8151",
    x"21A7EB1",
    x"21A7C12",
    x"21A7973",
    x"21A76D5",
    x"21A7438",
    x"21A719B",
    x"21A6EFF",
    x"21A6C64",
    x"21A69C9",
    x"21A672F",
    x"21A6495",
    x"21A61FD",
    x"21A5F64",
    x"21A5CCD",
    x"21A5A36",
    x"21A57A0",
    x"21A550A",
    x"21A5275",
    x"21A4FE1",
    x"21A4D4D",
    x"21A4ABA",
    x"21A4828",
    x"21A4596",
    x"21A4305",
    x"21A4075",
    x"21A3DE5",
    x"21A3B56",
    x"21A38C7",
    x"21A3639",
    x"21A33AC",
    x"21A311F",
    x"21A2E94",
    x"21A2C08",
    x"21A297E",
    x"21A26F3",
    x"21A246A",
    x"21A21E1",
    x"21A1F59",
    x"21A1CD2",
    x"21A1A4B",
    x"21A17C4",
    x"21A153F",
    x"21A12BA",
    x"21A1035",
    x"21A0DB2",
    x"21A0B2F",
    x"21A08AC",
    x"21A062A",
    x"21A03A9",
    x"21A0128",
    x"219FEA8",
    x"219FC29",
    x"219F9AA",
    x"219F72C",
    x"219F4AF",
    x"219F232",
    x"219EFB6",
    x"219ED3A",
    x"219EABF",
    x"219E845",
    x"219E5CB",
    x"219E352",
    x"219E0D9",
    x"219DE61",
    x"219DBEA",
    x"219D973",
    x"219D6FD",
    x"219D488",
    x"219D213",
    x"219CF9F",
    x"219CD2B",
    x"219CAB8",
    x"219C846",
    x"219C5D4",
    x"219C363",
    x"219C0F2",
    x"219BE83",
    x"219BC13",
    x"219B9A4",
    x"219B736",
    x"219B4C9",
    x"219B25C",
    x"219AFF0",
    x"219AD84",
    x"219AB19",
    x"219A8AE",
    x"219A645",
    x"219A3DB",
    x"219A173",
    x"2199F0B",
    x"2199CA3",
    x"2199A3C",
    x"21997D6",
    x"2199570",
    x"219930B",
    x"21990A7",
    x"2198E43",
    x"2198BE0",
    x"219897D",
    x"219871B",
    x"21984B9",
    x"2198259",
    x"2197FF8",
    x"2197D99",
    x"2197B3A",
    x"21978DB",
    x"219767D",
    x"2197420",
    x"21971C3",
    x"2196F67",
    x"2196D0B",
    x"2196AB0",
    x"2196856",
    x"21965FC",
    x"21963A3",
    x"219614A",
    x"2195EF2",
    x"2195C9B",
    x"2195A44",
    x"21957EE",
    x"2195598",
    x"2195343",
    x"21950EE",
    x"2194E9A",
    x"2194C47",
    x"21949F4",
    x"21947A2",
    x"2194551",
    x"21942FF",
    x"21940AF",
    x"2193E5F",
    x"2193C10",
    x"21939C1",
    x"2193773",
    x"2193525",
    x"21932D8",
    x"219308C",
    x"2192E40",
    x"2192BF5",
    x"21929AA",
    x"2192760",
    x"2192516",
    x"21922CD",
    x"2192085",
    x"2191E3D",
    x"2191BF6",
    x"21919AF",
    x"2191769",
    x"2191524",
    x"21912DF",
    x"219109A",
    x"2190E56",
    x"2190C13",
    x"21909D0",
    x"219078E",
    x"219054C",
    x"219030B",
    x"21900CB",
    x"218FE8B",
    x"218FC4C",
    x"218FA0D",
    x"218F7CF",
    x"218F591",
    x"218F354",
    x"218F117",
    x"218EEDB",
    x"218ECA0",
    x"218EA65",
    x"218E82B",
    x"218E5F1",
    x"218E3B8",
    x"218E17F",
    x"218DF47",
    x"218DD0F",
    x"218DAD8",
    x"218D8A2",
    x"218D66C",
    x"218D437",
    x"218D202",
    x"218CFCE",
    x"218CD9A",
    x"218CB67",
    x"218C934",
    x"218C702",
    x"218C4D1",
    x"218C2A0",
    x"218C06F",
    x"218BE40",
    x"218BC10",
    x"218B9E2",
    x"218B7B3",
    x"218B586",
    x"218B359",
    x"218B12C",
    x"218AF00",
    x"218ACD5",
    x"218AAAA",
    x"218A87F",
    x"218A655",
    x"218A42C",
    x"218A203",
    x"2189FDB",
    x"2189DB3",
    x"2189B8C",
    x"2189966",
    x"2189740",
    x"218951A",
    x"21892F5",
    x"21890D1",
    x"2188EAD",
    x"2188C89",
    x"2188A66",
    x"2188844",
    x"2188622",
    x"2188401",
    x"21881E0",
    x"2187FC0",
    x"2187DA0",
    x"2187B81",
    x"2187963",
    x"2187744",
    x"2187527",
    x"218730A",
    x"21870ED",
    x"2186ED1",
    x"2186CB6",
    x"2186A9B",
    x"2186881",
    x"2186667",
    x"218644D",
    x"2186235",
    x"218601C",
    x"2185E05",
    x"2185BED",
    x"21859D7",
    x"21857C0",
    x"21855AB",
    x"2185396",
    x"2185181",
    x"2184F6D",
    x"2184D59",
    x"2184B46",
    x"2184934",
    x"2184722",
    x"2184510",
    x"21842FF",
    x"21840EF",
    x"2183EDF",
    x"2183CCF",
    x"2183AC0",
    x"21838B2",
    x"21836A4",
    x"2183496",
    x"218328A",
    x"218307D",
    x"2182E71",
    x"2182C66",
    x"2182A5B",
    x"2182851",
    x"2182647",
    x"218243E",
    x"2182235",
    x"218202D",
    x"2181E25",
    x"2181C1D",
    x"2181A17",
    x"2181810",
    x"218160B",
    x"2181405",
    x"2181201",
    x"2180FFC",
    x"2180DF9",
    x"2180BF5",
    x"21809F3",
    x"21807F0",
    x"21805EF",
    x"21803ED",
    x"21801ED",
    x"217FFD9",
    x"217FBDA",
    x"217F7DB",
    x"217F3DE",
    x"217EFE2",
    x"217EBE6",
    x"217E7EC",
    x"217E3F2",
    x"217DFFA",
    x"217DC02",
    x"217D80C",
    x"217D416",
    x"217D022",
    x"217CC2E",
    x"217C83B",
    x"217C44A",
    x"217C059",
    x"217BC6A",
    x"217B87B",
    x"217B48E",
    x"217B0A1",
    x"217ACB5",
    x"217A8CA",
    x"217A4E1",
    x"217A0F8",
    x"2179D10",
    x"217992A",
    x"2179544",
    x"217915F",
    x"2178D7B",
    x"2178998",
    x"21785B6",
    x"21781D5",
    x"2177DF5",
    x"2177A16",
    x"2177638",
    x"217725B",
    x"2176E7F",
    x"2176AA4",
    x"21766CA",
    x"21762F1",
    x"2175F18",
    x"2175B41",
    x"217576B",
    x"2175395",
    x"2174FC1",
    x"2174BED",
    x"217481B",
    x"2174449",
    x"2174079",
    x"2173CA9",
    x"21738DA",
    x"217350D",
    x"2173140",
    x"2172D74",
    x"21729A9",
    x"21725DF",
    x"2172216",
    x"2171E4E",
    x"2171A87",
    x"21716C1",
    x"21712FC",
    x"2170F37",
    x"2170B74",
    x"21707B2",
    x"21703F0",
    x"2170030",
    x"216FC70",
    x"216F8B2",
    x"216F4F4",
    x"216F137",
    x"216ED7B",
    x"216E9C0",
    x"216E606",
    x"216E24D",
    x"216DE95",
    x"216DADE",
    x"216D728",
    x"216D372",
    x"216CFBE",
    x"216CC0B",
    x"216C858",
    x"216C4A6",
    x"216C0F6",
    x"216BD46",
    x"216B997",
    x"216B5E9",
    x"216B23C",
    x"216AE90",
    x"216AAE5",
    x"216A73B",
    x"216A391",
    x"2169FE9",
    x"2169C41",
    x"216989B",
    x"21694F5",
    x"2169150",
    x"2168DAC",
    x"2168A09",
    x"2168667",
    x"21682C6",
    x"2167F26",
    x"2167B87",
    x"21677E8",
    x"216744B",
    x"21670AE",
    x"2166D12",
    x"2166977",
    x"21665DD",
    x"2166244",
    x"2165EAC",
    x"2165B15",
    x"216577F",
    x"21653E9",
    x"2165055",
    x"2164CC1",
    x"216492E",
    x"216459D",
    x"216420C",
    x"2163E7C",
    x"2163AEC",
    x"216375E",
    x"21633D1",
    x"2163044",
    x"2162CB9",
    x"216292E",
    x"21625A4",
    x"216221B",
    x"2161E93",
    x"2161B0C",
    x"2161785",
    x"2161400",
    x"216107B",
    x"2160CF8",
    x"2160975",
    x"21605F3",
    x"2160272",
    x"215FEF2",
    x"215FB73",
    x"215F7F4",
    x"215F477",
    x"215F0FA",
    x"215ED7E",
    x"215EA03",
    x"215E689",
    x"215E310",
    x"215DF97",
    x"215DC20",
    x"215D8A9",
    x"215D534",
    x"215D1BF",
    x"215CE4B",
    x"215CAD8",
    x"215C765",
    x"215C3F4",
    x"215C083",
    x"215BD14",
    x"215B9A5",
    x"215B637",
    x"215B2CA",
    x"215AF5E",
    x"215ABF2",
    x"215A888",
    x"215A51E",
    x"215A1B5",
    x"2159E4D",
    x"2159AE6",
    x"2159780",
    x"215941A",
    x"21590B5",
    x"2158D52",
    x"21589EF",
    x"215868D",
    x"215832C",
    x"2157FCB",
    x"2157C6C",
    x"215790D",
    x"21575AF",
    x"2157252",
    x"2156EF6",
    x"2156B9B",
    x"2156840",
    x"21564E7",
    x"215618E",
    x"2155E36",
    x"2155ADF",
    x"2155788",
    x"2155433",
    x"21550DE",
    x"2154D8A",
    x"2154A37",
    x"21546E5",
    x"2154394",
    x"2154043",
    x"2153CF4",
    x"21539A5",
    x"2153657",
    x"215330A",
    x"2152FBD",
    x"2152C72",
    x"2152927",
    x"21525DD",
    x"2152294",
    x"2151F4C",
    x"2151C05",
    x"21518BE",
    x"2151578",
    x"2151233",
    x"2150EEF",
    x"2150BAC",
    x"2150869",
    x"2150528",
    x"21501E7",
    x"214FEA7",
    x"214FB67",
    x"214F829",
    x"214F4EB",
    x"214F1AF",
    x"214EE73",
    x"214EB37",
    x"214E7FD",
    x"214E4C3",
    x"214E18B",
    x"214DE53",
    x"214DB1B",
    x"214D7E5",
    x"214D4AF",
    x"214D17B",
    x"214CE47",
    x"214CB14",
    x"214C7E1",
    x"214C4B0",
    x"214C17F",
    x"214BE4F",
    x"214BB20",
    x"214B7F1",
    x"214B4C4",
    x"214B197",
    x"214AE6B",
    x"214AB40",
    x"214A815",
    x"214A4EC",
    x"214A1C3",
    x"2149E9B",
    x"2149B74",
    x"214984D",
    x"2149527",
    x"2149202",
    x"2148EDE",
    x"2148BBB",
    x"2148898",
    x"2148577",
    x"2148256",
    x"2147F36",
    x"2147C16",
    x"21478F8",
    x"21475DA",
    x"21472BD",
    x"2146FA0",
    x"2146C85",
    x"214696A",
    x"2146650",
    x"2146337",
    x"214601E",
    x"2145D07",
    x"21459F0",
    x"21456DA",
    x"21453C5",
    x"21450B0",
    x"2144D9C",
    x"2144A89",
    x"2144777",
    x"2144465",
    x"2144155",
    x"2143E45",
    x"2143B36",
    x"2143827",
    x"2143519",
    x"214320D",
    x"2142F00",
    x"2142BF5",
    x"21428EA",
    x"21425E1",
    x"21422D8",
    x"2141FCF",
    x"2141CC8",
    x"21419C1",
    x"21416BB",
    x"21413B5",
    x"21410B1",
    x"2140DAD",
    x"2140AAA",
    x"21407A8",
    x"21404A6",
    x"21401A5",
    x"213FEA5",
    x"213FBA6",
    x"213F8A8",
    x"213F5AA",
    x"213F2AD",
    x"213EFB0",
    x"213ECB5",
    x"213E9BA",
    x"213E6C0",
    x"213E3C7",
    x"213E0CE",
    x"213DDD6",
    x"213DADF",
    x"213D7E9",
    x"213D4F3",
    x"213D1FE",
    x"213CF0A",
    x"213CC17",
    x"213C924",
    x"213C632",
    x"213C341",
    x"213C051",
    x"213BD61",
    x"213BA72",
    x"213B784",
    x"213B496",
    x"213B1A9",
    x"213AEBD",
    x"213ABD2",
    x"213A8E7",
    x"213A5FE",
    x"213A314",
    x"213A02C",
    x"2139D44",
    x"2139A5D",
    x"2139777",
    x"2139492",
    x"21391AD",
    x"2138EC9",
    x"2138BE6",
    x"2138903",
    x"2138621",
    x"2138340",
    x"213805F",
    x"2137D80",
    x"2137AA1",
    x"21377C2",
    x"21374E5",
    x"2137208",
    x"2136F2C",
    x"2136C50",
    x"2136976",
    x"213669C",
    x"21363C2",
    x"21360EA",
    x"2135E12",
    x"2135B3B",
    x"2135864",
    x"213558E",
    x"21352B9",
    x"2134FE5",
    x"2134D11",
    x"2134A3F",
    x"213476C",
    x"213449B",
    x"21341CA",
    x"2133EFA",
    x"2133C2B",
    x"213395C",
    x"213368E",
    x"21333C1",
    x"21330F4",
    x"2132E28",
    x"2132B5D",
    x"2132892",
    x"21325C9",
    x"2132300",
    x"2132037",
    x"2131D6F",
    x"2131AA8",
    x"21317E2",
    x"213151C",
    x"2131258",
    x"2130F93",
    x"2130CD0",
    x"2130A0D",
    x"213074B",
    x"2130489",
    x"21301C8",
    x"212FF08",
    x"212FC49",
    x"212F98A",
    x"212F6CC",
    x"212F40F",
    x"212F152",
    x"212EE96",
    x"212EBDB",
    x"212E920",
    x"212E666",
    x"212E3AD",
    x"212E0F4",
    x"212DE3D",
    x"212DB85",
    x"212D8CF",
    x"212D619",
    x"212D364",
    x"212D0AF",
    x"212CDFB",
    x"212CB48",
    x"212C896",
    x"212C5E4",
    x"212C333",
    x"212C082",
    x"212BDD3",
    x"212BB23",
    x"212B875",
    x"212B5C7",
    x"212B31A",
    x"212B06E",
    x"212ADC2",
    x"212AB17",
    x"212A86C",
    x"212A5C3",
    x"212A319",
    x"212A071",
    x"2129DC9",
    x"2129B22",
    x"212987C",
    x"21295D6",
    x"2129331",
    x"212908C",
    x"2128DE8",
    x"2128B45",
    x"21288A3",
    x"2128601",
    x"2128360",
    x"21280BF",
    x"2127E1F",
    x"2127B80",
    x"21278E2",
    x"2127644",
    x"21273A7",
    x"212710A",
    x"2126E6E",
    x"2126BD3",
    x"2126938",
    x"212669E",
    x"2126405",
    x"212616C",
    x"2125ED4",
    x"2125C3D",
    x"21259A6",
    x"2125710",
    x"212547A",
    x"21251E6",
    x"2124F52",
    x"2124CBE",
    x"2124A2B",
    x"2124799",
    x"2124507",
    x"2124276",
    x"2123FE6",
    x"2123D56",
    x"2123AC7",
    x"2123839",
    x"21235AB",
    x"212331E",
    x"2123092",
    x"2122E06",
    x"2122B7B",
    x"21228F0",
    x"2122666",
    x"21223DD",
    x"2122154",
    x"2121ECC",
    x"2121C45",
    x"21219BE",
    x"2121738",
    x"21214B3",
    x"212122E",
    x"2120FAA",
    x"2120D26",
    x"2120AA3",
    x"2120821",
    x"212059F",
    x"212031E",
    x"212009D",
    x"211FE1D",
    x"211FB9E",
    x"211F920",
    x"211F6A2",
    x"211F424",
    x"211F1A8",
    x"211EF2C",
    x"211ECB0",
    x"211EA35",
    x"211E7BB",
    x"211E541",
    x"211E2C8",
    x"211E050",
    x"211DDD8",
    x"211DB61",
    x"211D8EA",
    x"211D675",
    x"211D3FF",
    x"211D18B",
    x"211CF16",
    x"211CCA3",
    x"211CA30",
    x"211C7BE",
    x"211C54C",
    x"211C2DB",
    x"211C06B",
    x"211BDFB",
    x"211BB8C",
    x"211B91D",
    x"211B6AF",
    x"211B442",
    x"211B1D5",
    x"211AF69",
    x"211ACFD",
    x"211AA92",
    x"211A828",
    x"211A5BE",
    x"211A355",
    x"211A0ED",
    x"2119E85",
    x"2119C1D",
    x"21199B7",
    x"2119751",
    x"21194EB",
    x"2119286",
    x"2119022",
    x"2118DBE",
    x"2118B5B",
    x"21188F8",
    x"2118696",
    x"2118435",
    x"21181D4",
    x"2117F74",
    x"2117D15",
    x"2117AB6",
    x"2117857",
    x"21175F9",
    x"211739C",
    x"2117140",
    x"2116EE4",
    x"2116C88",
    x"2116A2D",
    x"21167D3",
    x"2116579",
    x"2116320",
    x"21160C8",
    x"2115E70",
    x"2115C19",
    x"21159C2",
    x"211576C",
    x"2115516",
    x"21152C1",
    x"211506D",
    x"2114E19",
    x"2114BC6",
    x"2114973",
    x"2114721",
    x"21144D0",
    x"211427F",
    x"211402E",
    x"2113DDF",
    x"2113B8F",
    x"2113941",
    x"21136F3",
    x"21134A5",
    x"2113258",
    x"211300C",
    x"2112DC0",
    x"2112B75",
    x"211292B",
    x"21126E1",
    x"2112497",
    x"211224E",
    x"2112006",
    x"2111DBE",
    x"2111B77",
    x"2111931",
    x"21116EB",
    x"21114A5",
    x"2111260",
    x"211101C",
    x"2110DD8",
    x"2110B95",
    x"2110952",
    x"2110710",
    x"21104CF",
    x"211028E",
    x"211004E",
    x"210FE0E",
    x"210FBCF",
    x"210F990",
    x"210F752",
    x"210F514",
    x"210F2D7",
    x"210F09B",
    x"210EE5F",
    x"210EC24",
    x"210E9E9",
    x"210E7AF",
    x"210E575",
    x"210E33C",
    x"210E103",
    x"210DECC",
    x"210DC94",
    x"210DA5D",
    x"210D827",
    x"210D5F1",
    x"210D3BC",
    x"210D187",
    x"210CF53",
    x"210CD20",
    x"210CAED",
    x"210C8BA",
    x"210C688",
    x"210C457",
    x"210C226",
    x"210BFF6",
    x"210BDC6",
    x"210BB97",
    x"210B968",
    x"210B73A",
    x"210B50D",
    x"210B2E0",
    x"210B0B3",
    x"210AE87",
    x"210AC5C",
    x"210AA31",
    x"210A807",
    x"210A5DD",
    x"210A3B4",
    x"210A18B",
    x"2109F63",
    x"2109D3C",
    x"2109B15",
    x"21098EE",
    x"21096C8",
    x"21094A3",
    x"210927E",
    x"2109059",
    x"2108E36",
    x"2108C12",
    x"21089F0",
    x"21087CD",
    x"21085AC",
    x"210838B",
    x"210816A",
    x"2107F4A",
    x"2107D2A",
    x"2107B0B",
    x"21078ED",
    x"21076CF",
    x"21074B1",
    x"2107294",
    x"2107078",
    x"2106E5C",
    x"2106C41",
    x"2106A26",
    x"210680C",
    x"21065F2",
    x"21063D9",
    x"21061C0",
    x"2105FA8",
    x"2105D90",
    x"2105B79",
    x"2105963",
    x"210574C",
    x"2105537",
    x"2105322",
    x"210510D",
    x"2104EF9",
    x"2104CE6",
    x"2104AD3",
    x"21048C0",
    x"21046AE",
    x"210449D",
    x"210428C",
    x"210407C",
    x"2103E6C",
    x"2103C5D",
    x"2103A4E",
    x"210383F",
    x"2103632",
    x"2103424",
    x"2103218",
    x"210300B",
    x"2102E00",
    x"2102BF4",
    x"21029EA",
    x"21027DF",
    x"21025D6",
    x"21023CC",
    x"21021C4",
    x"2101FBC",
    x"2101DB4",
    x"2101BAD",
    x"21019A6",
    x"21017A0",
    x"210159A",
    x"2101395",
    x"2101190",
    x"2100F8C",
    x"2100D89",
    x"2100B85",
    x"2100983",
    x"2100781",
    x"210057F",
    x"210037E",
    x"210017D",
    x"20FFEFB",
    x"20FFAFC",
    x"20FF6FD",
    x"20FF300",
    x"20FEF04",
    x"20FEB09",
    x"20FE70E",
    x"20FE315",
    x"20FDF1D",
    x"20FDB26",
    x"20FD72F",
    x"20FD33A",
    x"20FCF46",
    x"20FCB52",
    x"20FC760",
    x"20FC36F",
    x"20FBF7E",
    x"20FBB8F",
    x"20FB7A1",
    x"20FB3B3",
    x"20FAFC7",
    x"20FABDB",
    x"20FA7F1",
    x"20FA407",
    x"20FA01F",
    x"20F9C37",
    x"20F9851",
    x"20F946B",
    x"20F9086",
    x"20F8CA3",
    x"20F88C0",
    x"20F84DE",
    x"20F80FE",
    x"20F7D1E",
    x"20F793F",
    x"20F7561",
    x"20F7184",
    x"20F6DA9",
    x"20F69CE",
    x"20F65F4",
    x"20F621B",
    x"20F5E43",
    x"20F5A6B",
    x"20F5695",
    x"20F52C0",
    x"20F4EEC",
    x"20F4B19",
    x"20F4746",
    x"20F4375",
    x"20F3FA5",
    x"20F3BD5",
    x"20F3807",
    x"20F3439",
    x"20F306D",
    x"20F2CA1",
    x"20F28D6",
    x"20F250D",
    x"20F2144",
    x"20F1D7C",
    x"20F19B5",
    x"20F15EF",
    x"20F122A",
    x"20F0E66",
    x"20F0AA3",
    x"20F06E1",
    x"20F031F",
    x"20EFF5F",
    x"20EFBA0",
    x"20EF7E1",
    x"20EF424",
    x"20EF067",
    x"20EECAC",
    x"20EE8F1",
    x"20EE537",
    x"20EE17E",
    x"20EDDC6",
    x"20EDA0F",
    x"20ED659",
    x"20ED2A4",
    x"20ECEF0",
    x"20ECB3D",
    x"20EC78A",
    x"20EC3D9",
    x"20EC029",
    x"20EBC79",
    x"20EB8CA",
    x"20EB51D",
    x"20EB170",
    x"20EADC4",
    x"20EAA19",
    x"20EA66F",
    x"20EA2C6",
    x"20E9F1D",
    x"20E9B76",
    x"20E97D0",
    x"20E942A",
    x"20E9086",
    x"20E8CE2",
    x"20E893F",
    x"20E859D",
    x"20E81FC",
    x"20E7E5C",
    x"20E7ABD",
    x"20E771F",
    x"20E7382",
    x"20E6FE5",
    x"20E6C4A",
    x"20E68AF",
    x"20E6515",
    x"20E617C",
    x"20E5DE5",
    x"20E5A4E",
    x"20E56B7",
    x"20E5322",
    x"20E4F8E",
    x"20E4BFA",
    x"20E4868",
    x"20E44D6",
    x"20E4145",
    x"20E3DB6",
    x"20E3A27",
    x"20E3698",
    x"20E330B",
    x"20E2F7F",
    x"20E2BF4",
    x"20E2869",
    x"20E24DF",
    x"20E2157",
    x"20E1DCF",
    x"20E1A48",
    x"20E16C1",
    x"20E133C",
    x"20E0FB8",
    x"20E0C34",
    x"20E08B2",
    x"20E0530",
    x"20E01AF",
    x"20DFE2F",
    x"20DFAB0",
    x"20DF732",
    x"20DF3B4",
    x"20DF038",
    x"20DECBC",
    x"20DE942",
    x"20DE5C8",
    x"20DE24F",
    x"20DDED7",
    x"20DDB5F",
    x"20DD7E9",
    x"20DD473",
    x"20DD0FF",
    x"20DCD8B",
    x"20DCA18",
    x"20DC6A6",
    x"20DC335",
    x"20DBFC4",
    x"20DBC55",
    x"20DB8E6",
    x"20DB578",
    x"20DB20B",
    x"20DAE9F",
    x"20DAB34",
    x"20DA7CA",
    x"20DA460",
    x"20DA0F7",
    x"20D9D90",
    x"20D9A29",
    x"20D96C3",
    x"20D935D",
    x"20D8FF9",
    x"20D8C95",
    x"20D8933",
    x"20D85D1",
    x"20D8270",
    x"20D7F0F",
    x"20D7BB0",
    x"20D7852",
    x"20D74F4",
    x"20D7197",
    x"20D6E3B",
    x"20D6AE0",
    x"20D6786",
    x"20D642C",
    x"20D60D4",
    x"20D5D7C",
    x"20D5A25",
    x"20D56CF",
    x"20D5379",
    x"20D5025",
    x"20D4CD1",
    x"20D497F",
    x"20D462D",
    x"20D42DC",
    x"20D3F8B",
    x"20D3C3C",
    x"20D38ED",
    x"20D359F",
    x"20D3252",
    x"20D2F06",
    x"20D2BBB",
    x"20D2870",
    x"20D2527",
    x"20D21DE",
    x"20D1E96",
    x"20D1B4E",
    x"20D1808",
    x"20D14C2",
    x"20D117E",
    x"20D0E3A",
    x"20D0AF6",
    x"20D07B4",
    x"20D0473",
    x"20D0132",
    x"20CFDF2",
    x"20CFAB3",
    x"20CF775",
    x"20CF437",
    x"20CF0FB",
    x"20CEDBF",
    x"20CEA84",
    x"20CE749",
    x"20CE410",
    x"20CE0D7",
    x"20CDDA0",
    x"20CDA69",
    x"20CD732",
    x"20CD3FD",
    x"20CD0C8",
    x"20CCD95",
    x"20CCA62",
    x"20CC72F",
    x"20CC3FE",
    x"20CC0CD",
    x"20CBD9E",
    x"20CBA6F",
    x"20CB740",
    x"20CB413",
    x"20CB0E6",
    x"20CADBB",
    x"20CAA90",
    x"20CA765",
    x"20CA43C",
    x"20CA113",
    x"20C9DEB",
    x"20C9AC4",
    x"20C979E",
    x"20C9478",
    x"20C9154",
    x"20C8E30",
    x"20C8B0D",
    x"20C87EA",
    x"20C84C9",
    x"20C81A8",
    x"20C7E88",
    x"20C7B69",
    x"20C784A",
    x"20C752C",
    x"20C720F",
    x"20C6EF3",
    x"20C6BD8",
    x"20C68BD",
    x"20C65A4",
    x"20C628B",
    x"20C5F72",
    x"20C5C5B",
    x"20C5944",
    x"20C562E",
    x"20C5319",
    x"20C5005",
    x"20C4CF1",
    x"20C49DE",
    x"20C46CC",
    x"20C43BB",
    x"20C40AA",
    x"20C3D9B",
    x"20C3A8B",
    x"20C377D",
    x"20C3470",
    x"20C3163",
    x"20C2E57",
    x"20C2B4C",
    x"20C2841",
    x"20C2538",
    x"20C222F",
    x"20C1F27",
    x"20C1C1F",
    x"20C1919",
    x"20C1613",
    x"20C130E",
    x"20C1009",
    x"20C0D05",
    x"20C0A03",
    x"20C0700",
    x"20C03FF",
    x"20C00FE",
    x"20BFDFF",
    x"20BFAFF",
    x"20BF801",
    x"20BF503",
    x"20BF207",
    x"20BEF0A",
    x"20BEC0F",
    x"20BE914",
    x"20BE61B",
    x"20BE321",
    x"20BE029",
    x"20BDD31",
    x"20BDA3A",
    x"20BD744",
    x"20BD44F",
    x"20BD15A",
    x"20BCE66",
    x"20BCB73",
    x"20BC880",
    x"20BC58F",
    x"20BC29E",
    x"20BBFAD",
    x"20BBCBE",
    x"20BB9CF",
    x"20BB6E1",
    x"20BB3F3",
    x"20BB107",
    x"20BAE1B",
    x"20BAB30",
    x"20BA845",
    x"20BA55C",
    x"20BA273",
    x"20B9F8A",
    x"20B9CA3",
    x"20B99BC",
    x"20B96D6",
    x"20B93F1",
    x"20B910C",
    x"20B8E28",
    x"20B8B45",
    x"20B8863",
    x"20B8581",
    x"20B82A0",
    x"20B7FBF",
    x"20B7CE0",
    x"20B7A01",
    x"20B7723",
    x"20B7445",
    x"20B7169",
    x"20B6E8D",
    x"20B6BB1",
    x"20B68D7",
    x"20B65FD",
    x"20B6324",
    x"20B604B",
    x"20B5D74",
    x"20B5A9D",
    x"20B57C6",
    x"20B54F1",
    x"20B521C",
    x"20B4F48",
    x"20B4C74",
    x"20B49A2",
    x"20B46D0",
    x"20B43FE",
    x"20B412E",
    x"20B3E5E",
    x"20B3B8E",
    x"20B38C0",
    x"20B35F2",
    x"20B3325",
    x"20B3058",
    x"20B2D8D",
    x"20B2AC2",
    x"20B27F7",
    x"20B252E",
    x"20B2265",
    x"20B1F9C",
    x"20B1CD5",
    x"20B1A0E",
    x"20B1748",
    x"20B1482",
    x"20B11BE",
    x"20B0EFA",
    x"20B0C36",
    x"20B0973",
    x"20B06B1",
    x"20B03F0",
    x"20B012F",
    x"20AFE6F",
    x"20AFBB0",
    x"20AF8F2",
    x"20AF634",
    x"20AF377",
    x"20AF0BA",
    x"20AEDFE",
    x"20AEB43",
    x"20AE889",
    x"20AE5CF",
    x"20AE316",
    x"20AE05D",
    x"20ADDA5",
    x"20ADAEE",
    x"20AD838",
    x"20AD582",
    x"20AD2CD",
    x"20AD019",
    x"20ACD65",
    x"20ACAB2",
    x"20AC800",
    x"20AC54E",
    x"20AC29D",
    x"20ABFED",
    x"20ABD3D",
    x"20ABA8E",
    x"20AB7E0",
    x"20AB532",
    x"20AB285",
    x"20AAFD9",
    x"20AAD2D",
    x"20AAA82",
    x"20AA7D8",
    x"20AA52F",
    x"20AA286",
    x"20A9FDD",
    x"20A9D36",
    x"20A9A8F",
    x"20A97E8",
    x"20A9543",
    x"20A929E",
    x"20A8FF9",
    x"20A8D56",
    x"20A8AB3",
    x"20A8810",
    x"20A856F",
    x"20A82CE",
    x"20A802D",
    x"20A7D8E",
    x"20A7AEF",
    x"20A7850",
    x"20A75B2",
    x"20A7315",
    x"20A7079",
    x"20A6DDD",
    x"20A6B42",
    x"20A68A7",
    x"20A660E",
    x"20A6374",
    x"20A60DC",
    x"20A5E44",
    x"20A5BAD",
    x"20A5916",
    x"20A5680",
    x"20A53EB",
    x"20A5156",
    x"20A4EC2",
    x"20A4C2F",
    x"20A499C",
    x"20A470A",
    x"20A4479",
    x"20A41E8",
    x"20A3F58",
    x"20A3CC8",
    x"20A3A39",
    x"20A37AB",
    x"20A351D",
    x"20A3290",
    x"20A3004",
    x"20A2D78",
    x"20A2AED",
    x"20A2863",
    x"20A25D9",
    x"20A2350",
    x"20A20C7",
    x"20A1E40",
    x"20A1BB8",
    x"20A1932",
    x"20A16AC",
    x"20A1426",
    x"20A11A2",
    x"20A0F1E",
    x"20A0C9A",
    x"20A0A17",
    x"20A0795",
    x"20A0514",
    x"20A0293",
    x"20A0012",
    x"209FD93",
    x"209FB13",
    x"209F895",
    x"209F617",
    x"209F39A",
    x"209F11D",
    x"209EEA1",
    x"209EC26",
    x"209E9AB",
    x"209E731",
    x"209E4B8",
    x"209E23F",
    x"209DFC7",
    x"209DD4F",
    x"209DAD8",
    x"209D862",
    x"209D5EC",
    x"209D377",
    x"209D102",
    x"209CE8E",
    x"209CC1B",
    x"209C9A8",
    x"209C736",
    x"209C4C4",
    x"209C254",
    x"209BFE3",
    x"209BD74",
    x"209BB04",
    x"209B896",
    x"209B628",
    x"209B3BB",
    x"209B14E",
    x"209AEE2",
    x"209AC77",
    x"209AA0C",
    x"209A7A2",
    x"209A538",
    x"209A2CF",
    x"209A067",
    x"2099DFF",
    x"2099B98",
    x"2099931",
    x"20996CB",
    x"2099466",
    x"2099201",
    x"2098F9D",
    x"2098D39",
    x"2098AD6",
    x"2098874",
    x"2098612",
    x"20983B1",
    x"2098150",
    x"2097EF0",
    x"2097C91",
    x"2097A32",
    x"20977D4",
    x"2097576",
    x"2097319",
    x"20970BC",
    x"2096E61",
    x"2096C05",
    x"20969AA",
    x"2096750",
    x"20964F7",
    x"209629E",
    x"2096046",
    x"2095DEE",
    x"2095B97",
    x"2095940",
    x"20956EA",
    x"2095494",
    x"2095240",
    x"2094FEB",
    x"2094D98",
    x"2094B45",
    x"20948F2",
    x"20946A0",
    x"209444F",
    x"20941FE",
    x"2093FAE",
    x"2093D5E",
    x"2093B0F",
    x"20938C1",
    x"2093673",
    x"2093425",
    x"20931D9",
    x"2092F8C",
    x"2092D41",
    x"2092AF6",
    x"20928AB",
    x"2092661",
    x"2092418",
    x"20921CF",
    x"2091F87",
    x"2091D40",
    x"2091AF9",
    x"20918B2",
    x"209166C",
    x"2091427",
    x"20911E2",
    x"2090F9E",
    x"2090D5A",
    x"2090B17",
    x"20908D5",
    x"2090693",
    x"2090452",
    x"2090211",
    x"208FFD1",
    x"208FD91",
    x"208FB52",
    x"208F913",
    x"208F6D5",
    x"208F498",
    x"208F25B",
    x"208F01F",
    x"208EDE3",
    x"208EBA8",
    x"208E96D",
    x"208E733",
    x"208E4F9",
    x"208E2C0",
    x"208E088",
    x"208DE50",
    x"208DC19",
    x"208D9E2",
    x"208D7AC",
    x"208D576",
    x"208D341",
    x"208D10D",
    x"208CED9",
    x"208CCA5",
    x"208CA72",
    x"208C840",
    x"208C60E",
    x"208C3DD",
    x"208C1AC",
    x"208BF7C",
    x"208BD4D",
    x"208BB1D",
    x"208B8EF",
    x"208B6C1",
    x"208B494",
    x"208B267",
    x"208B03A",
    x"208AE0F",
    x"208ABE3",
    x"208A9B9",
    x"208A78F",
    x"208A565",
    x"208A33C",
    x"208A113",
    x"2089EEB",
    x"2089CC4",
    x"2089A9D",
    x"2089877",
    x"2089651",
    x"208942B",
    x"2089207",
    x"2088FE2",
    x"2088DBF",
    x"2088B9B",
    x"2088979",
    x"2088757",
    x"2088535",
    x"2088314",
    x"20880F4",
    x"2087ED4",
    x"2087CB4",
    x"2087A95",
    x"2087877",
    x"2087659",
    x"208743C",
    x"208721F",
    x"2087003",
    x"2086DE7",
    x"2086BCC",
    x"20869B1",
    x"2086797",
    x"208657D",
    x"2086364",
    x"208614C",
    x"2085F33",
    x"2085D1C",
    x"2085B05",
    x"20858EE",
    x"20856D8",
    x"20854C3",
    x"20852AE",
    x"208509A",
    x"2084E86",
    x"2084C72",
    x"2084A60",
    x"208484D",
    x"208463B",
    x"208442A",
    x"2084219",
    x"2084009",
    x"2083DF9",
    x"2083BEA",
    x"20839DB",
    x"20837CD",
    x"20835BF",
    x"20833B2",
    x"20831A6",
    x"2082F99",
    x"2082D8E",
    x"2082B83",
    x"2082978",
    x"208276E",
    x"2082564",
    x"208235B",
    x"2082153",
    x"2081F4B",
    x"2081D43",
    x"2081B3C",
    x"2081935",
    x"208172F",
    x"208152A",
    x"2081325",
    x"2081120",
    x"2080F1C",
    x"2080D19",
    x"2080B16",
    x"2080913",
    x"2080711",
    x"2080510",
    x"208030F",
    x"208010E",
    x"207FE1D",
    x"207FA1D",
    x"207F61F",
    x"207F222",
    x"207EE26",
    x"207EA2B",
    x"207E631",
    x"207E238",
    x"207DE40",
    x"207DA49",
    x"207D653",
    x"207D25E",
    x"207CE6A",
    x"207CA77",
    x"207C685",
    x"207C293",
    x"207BEA3",
    x"207BAB4",
    x"207B6C6",
    x"207B2D9",
    x"207AEED",
    x"207AB01",
    x"207A717",
    x"207A32E",
    x"2079F45",
    x"2079B5E",
    x"2079778",
    x"2079392",
    x"2078FAE",
    x"2078BCB",
    x"20787E8",
    x"2078407",
    x"2078026",
    x"2077C47",
    x"2077868",
    x"207748A",
    x"20770AE",
    x"2076CD2",
    x"20768F7",
    x"207651E",
    x"2076145",
    x"2075D6D",
    x"2075996",
    x"20755C0",
    x"20751EB",
    x"2074E17",
    x"2074A44",
    x"2074672",
    x"20742A1",
    x"2073ED1",
    x"2073B01",
    x"2073733",
    x"2073366",
    x"2072F99",
    x"2072BCE",
    x"2072804",
    x"207243A",
    x"2072071",
    x"2071CAA",
    x"20718E3",
    x"207151D",
    x"2071159",
    x"2070D95",
    x"20709D2",
    x"2070610",
    x"207024F",
    x"206FE8F",
    x"206FACF",
    x"206F711",
    x"206F354",
    x"206EF98",
    x"206EBDC",
    x"206E822",
    x"206E468",
    x"206E0AF",
    x"206DCF8",
    x"206D941",
    x"206D58B",
    x"206D1D6",
    x"206CE22",
    x"206CA6F",
    x"206C6BD",
    x"206C30C",
    x"206BF5B",
    x"206BBAC",
    x"206B7FE",
    x"206B450",
    x"206B0A3",
    x"206ACF8",
    x"206A94D",
    x"206A5A3",
    x"206A1FA",
    x"2069E52",
    x"2069AAB",
    x"2069705",
    x"206935F",
    x"2068FBB",
    x"2068C18",
    x"2068875",
    x"20684D3",
    x"2068133",
    x"2067D93",
    x"20679F4",
    x"2067656",
    x"20672B9",
    x"2066F1C",
    x"2066B81",
    x"20667E7",
    x"206644D",
    x"20660B5",
    x"2065D1D",
    x"2065986",
    x"20655F0",
    x"206525B",
    x"2064EC7",
    x"2064B34",
    x"20647A1",
    x"2064410",
    x"206407F",
    x"2063CF0",
    x"2063961",
    x"20635D3",
    x"2063246",
    x"2062EBA",
    x"2062B2E",
    x"20627A4",
    x"206241B",
    x"2062092",
    x"2061D0A",
    x"2061984",
    x"20615FE",
    x"2061279",
    x"2060EF4",
    x"2060B71",
    x"20607EF",
    x"206046D",
    x"20600EC",
    x"205FD6D",
    x"205F9EE",
    x"205F670",
    x"205F2F2",
    x"205EF76",
    x"205EBFB",
    x"205E880",
    x"205E506",
    x"205E18E",
    x"205DE16",
    x"205DA9F",
    x"205D728",
    x"205D3B3",
    x"205D03F",
    x"205CCCB",
    x"205C958",
    x"205C5E6",
    x"205C275",
    x"205BF05",
    x"205BB96",
    x"205B827",
    x"205B4BA",
    x"205B14D",
    x"205ADE1",
    x"205AA76",
    x"205A70C",
    x"205A3A2",
    x"205A03A",
    x"2059CD2",
    x"205996C",
    x"2059606",
    x"20592A0",
    x"2058F3C",
    x"2058BD9",
    x"2058876",
    x"2058515",
    x"20581B4",
    x"2057E54",
    x"2057AF5",
    x"2057796",
    x"2057439",
    x"20570DC",
    x"2056D80",
    x"2056A25",
    x"20566CB",
    x"2056372",
    x"205601A",
    x"2055CC2",
    x"205596B",
    x"2055615",
    x"20552C0",
    x"2054F6C",
    x"2054C18",
    x"20548C6",
    x"2054574",
    x"2054223",
    x"2053ED3",
    x"2053B84",
    x"2053835",
    x"20534E8",
    x"205319B",
    x"2052E4F",
    x"2052B04",
    x"20527B9",
    x"2052470",
    x"2052127",
    x"2051DDF",
    x"2051A98",
    x"2051752",
    x"205140C",
    x"20510C8",
    x"2050D84",
    x"2050A41",
    x"20506FF",
    x"20503BE",
    x"205007D",
    x"204FD3D",
    x"204F9FE",
    x"204F6C0",
    x"204F383",
    x"204F047",
    x"204ED0B",
    x"204E9D0",
    x"204E696",
    x"204E35D",
    x"204E024",
    x"204DCED",
    x"204D9B6",
    x"204D680",
    x"204D34B",
    x"204D016",
    x"204CCE3",
    x"204C9B0",
    x"204C67E",
    x"204C34D",
    x"204C01C",
    x"204BCEC",
    x"204B9BE",
    x"204B690",
    x"204B362",
    x"204B036",
    x"204AD0A",
    x"204A9DF",
    x"204A6B5",
    x"204A38C",
    x"204A064",
    x"2049D3C",
    x"2049A15",
    x"20496EF",
    x"20493C9",
    x"20490A5",
    x"2048D81",
    x"2048A5E",
    x"204873C",
    x"204841B",
    x"20480FA",
    x"2047DDA",
    x"2047ABB",
    x"204779D",
    x"204747F",
    x"2047162",
    x"2046E46",
    x"2046B2B",
    x"2046811",
    x"20464F7",
    x"20461DE",
    x"2045EC6",
    x"2045BAF",
    x"2045898",
    x"2045583",
    x"204526E",
    x"2044F5A",
    x"2044C46",
    x"2044933",
    x"2044621",
    x"2044310",
    x"2044000",
    x"2043CF0",
    x"20439E1",
    x"20436D3",
    x"20433C6",
    x"20430B9",
    x"2042DAE",
    x"2042AA3",
    x"2042798",
    x"204248F",
    x"2042186",
    x"2041E7E",
    x"2041B77",
    x"2041870",
    x"204156B",
    x"2041266",
    x"2040F61",
    x"2040C5E",
    x"204095B",
    x"2040659",
    x"2040358",
    x"2040058",
    x"203FD58",
    x"203FA59",
    x"203F75B",
    x"203F45D",
    x"203F161",
    x"203EE65",
    x"203EB69",
    x"203E86F",
    x"203E575",
    x"203E27C",
    x"203DF84",
    x"203DC8C",
    x"203D996",
    x"203D6A0",
    x"203D3AA",
    x"203D0B6",
    x"203CDC2",
    x"203CACF",
    x"203C7DD",
    x"203C4EB",
    x"203C1FA",
    x"203BF0A",
    x"203BC1B",
    x"203B92C",
    x"203B63E",
    x"203B351",
    x"203B064",
    x"203AD79",
    x"203AA8E",
    x"203A7A3",
    x"203A4BA",
    x"203A1D1",
    x"2039EE9",
    x"2039C01",
    x"203991B",
    x"2039635",
    x"2039350",
    x"203906B",
    x"2038D87",
    x"2038AA4",
    x"20387C2",
    x"20384E1",
    x"2038200",
    x"2037F20",
    x"2037C40",
    x"2037961",
    x"2037683",
    x"20373A6",
    x"20370CA",
    x"2036DEE",
    x"2036B13",
    x"2036838",
    x"203655F",
    x"2036286",
    x"2035FAD",
    x"2035CD6",
    x"20359FF",
    x"2035729",
    x"2035453",
    x"203517F",
    x"2034EAB",
    x"2034BD7",
    x"2034905",
    x"2034633",
    x"2034362",
    x"2034091",
    x"2033DC1",
    x"2033AF2",
    x"2033824",
    x"2033556",
    x"2033289",
    x"2032FBD",
    x"2032CF1",
    x"2032A26",
    x"203275C",
    x"2032493",
    x"20321CA",
    x"2031F02",
    x"2031C3A",
    x"2031974",
    x"20316AE",
    x"20313E8",
    x"2031124",
    x"2030E60",
    x"2030B9D",
    x"20308DA",
    x"2030618",
    x"2030357",
    x"2030096",
    x"202FDD7",
    x"202FB17",
    x"202F859",
    x"202F59B",
    x"202F2DE",
    x"202F022",
    x"202ED66",
    x"202EAAB",
    x"202E7F1",
    x"202E537",
    x"202E27E",
    x"202DFC6",
    x"202DD0E",
    x"202DA57",
    x"202D7A1",
    x"202D4EC",
    x"202D237",
    x"202CF83",
    x"202CCCF",
    x"202CA1C",
    x"202C76A",
    x"202C4B8",
    x"202C208",
    x"202BF57",
    x"202BCA8",
    x"202B9F9",
    x"202B74B",
    x"202B49D",
    x"202B1F1",
    x"202AF44",
    x"202AC99",
    x"202A9EE",
    x"202A744",
    x"202A49A",
    x"202A1F2",
    x"2029F4A",
    x"2029CA2",
    x"20299FB",
    x"2029755",
    x"20294B0",
    x"202920B",
    x"2028F67",
    x"2028CC3",
    x"2028A20",
    x"202877E",
    x"20284DC",
    x"202823B",
    x"2027F9B",
    x"2027CFC",
    x"2027A5D",
    x"20277BF",
    x"2027521",
    x"2027284",
    x"2026FE8",
    x"2026D4C",
    x"2026AB1",
    x"2026817",
    x"202657D",
    x"20262E4",
    x"202604C",
    x"2025DB4",
    x"2025B1D",
    x"2025886",
    x"20255F0",
    x"202535B",
    x"20250C7",
    x"2024E33",
    x"2024BA0",
    x"202490D",
    x"202467B",
    x"20243EA",
    x"2024159",
    x"2023EC9",
    x"2023C3A",
    x"20239AB",
    x"202371D",
    x"202348F",
    x"2023203",
    x"2022F76",
    x"2022CEB",
    x"2022A60",
    x"20227D6",
    x"202254C",
    x"20222C3",
    x"202203B",
    x"2021DB3",
    x"2021B2C",
    x"20218A5",
    x"202161F",
    x"202139A",
    x"2021116",
    x"2020E92",
    x"2020C0E",
    x"202098C",
    x"202070A",
    x"2020488",
    x"2020207",
    x"201FF87",
    x"201FD08",
    x"201FA89",
    x"201F80A",
    x"201F58D",
    x"201F310",
    x"201F093",
    x"201EE17",
    x"201EB9C",
    x"201E921",
    x"201E6A7",
    x"201E42E",
    x"201E1B5",
    x"201DF3D",
    x"201DCC6",
    x"201DA4F",
    x"201D7D9",
    x"201D563",
    x"201D2EE",
    x"201D079",
    x"201CE06",
    x"201CB92",
    x"201C920",
    x"201C6AE",
    x"201C43D",
    x"201C1CC",
    x"201BF5C",
    x"201BCEC",
    x"201BA7D",
    x"201B80F",
    x"201B5A1",
    x"201B334",
    x"201B0C8",
    x"201AE5C",
    x"201ABF0",
    x"201A986",
    x"201A71C",
    x"201A4B2",
    x"201A249",
    x"2019FE1",
    x"2019D79",
    x"2019B12",
    x"20198AC",
    x"2019646",
    x"20193E1",
    x"201917C",
    x"2018F18",
    x"2018CB4",
    x"2018A52",
    x"20187EF",
    x"201858E",
    x"201832D",
    x"20180CC",
    x"2017E6C",
    x"2017C0D",
    x"20179AE",
    x"2017750",
    x"20174F2",
    x"2017295",
    x"2017039",
    x"2016DDD",
    x"2016B82",
    x"2016928",
    x"20166CE",
    x"2016474",
    x"201621B",
    x"2015FC3",
    x"2015D6C",
    x"2015B14",
    x"20158BE",
    x"2015668",
    x"2015413",
    x"20151BE",
    x"2014F6A",
    x"2014D16",
    x"2014AC3",
    x"2014871",
    x"201461F",
    x"20143CE",
    x"201417D",
    x"2013F2D",
    x"2013CDE",
    x"2013A8F",
    x"2013840",
    x"20135F3",
    x"20133A5",
    x"2013159",
    x"2012F0D",
    x"2012CC1",
    x"2012A76",
    x"201282C",
    x"20125E2",
    x"2012399",
    x"2012150",
    x"2011F08",
    x"2011CC1",
    x"2011A7A",
    x"2011834",
    x"20115EE",
    x"20113A9",
    x"2011164",
    x"2010F20",
    x"2010CDD",
    x"2010A9A",
    x"2010857",
    x"2010615",
    x"20103D4",
    x"2010193",
    x"200FF53",
    x"200FD14",
    x"200FAD5",
    x"200F896",
    x"200F659",
    x"200F41B",
    x"200F1DE",
    x"200EFA2",
    x"200ED67",
    x"200EB2C",
    x"200E8F1",
    x"200E6B7",
    x"200E47E",
    x"200E245",
    x"200E00D",
    x"200DDD5",
    x"200DB9E",
    x"200D967",
    x"200D731",
    x"200D4FB",
    x"200D2C6",
    x"200D092",
    x"200CE5E",
    x"200CC2B",
    x"200C9F8",
    x"200C7C6",
    x"200C594",
    x"200C363",
    x"200C133",
    x"200BF03",
    x"200BCD3",
    x"200BAA4",
    x"200B876",
    x"200B648",
    x"200B41B",
    x"200B1EE",
    x"200AFC2",
    x"200AD96",
    x"200AB6B",
    x"200A940",
    x"200A716",
    x"200A4ED",
    x"200A2C4",
    x"200A09B",
    x"2009E73",
    x"2009C4C",
    x"2009A25",
    x"20097FF",
    x"20095D9",
    x"20093B4",
    x"200918F",
    x"2008F6B",
    x"2008D48",
    x"2008B25",
    x"2008902",
    x"20086E0",
    x"20084BF",
    x"200829E",
    x"200807D",
    x"2007E5E",
    x"2007C3E",
    x"2007A1F",
    x"2007801",
    x"20075E3",
    x"20073C6",
    x"20071AA",
    x"2006F8D",
    x"2006D72",
    x"2006B57",
    x"200693C",
    x"2006722",
    x"2006508",
    x"20062EF",
    x"20060D7",
    x"2005EBF",
    x"2005CA8",
    x"2005A91",
    x"200587A",
    x"2005665",
    x"200544F",
    x"200523A",
    x"2005026",
    x"2004E12",
    x"2004BFF",
    x"20049EC",
    x"20047DA",
    x"20045C8",
    x"20043B7",
    x"20041A6",
    x"2003F96",
    x"2003D87",
    x"2003B78",
    x"2003969",
    x"200375B",
    x"200354D",
    x"2003340",
    x"2003134",
    x"2002F28",
    x"2002D1C",
    x"2002B11",
    x"2002907",
    x"20026FD",
    x"20024F3",
    x"20022EA",
    x"20020E2",
    x"2001EDA",
    x"2001CD2",
    x"2001ACB",
    x"20018C5",
    x"20016BF",
    x"20014B9",
    x"20012B4",
    x"20010B0",
    x"2000EAC",
    x"2000CA9",
    x"2000AA6",
    x"20008A3",
    x"20006A1",
    x"20004A0",
    x"200029F",
    x"200009F",
    x"1FFFD3E",
    x"1FFF93F",
    x"1FFF542",
    x"1FFF145",
    x"1FFED49",
    x"1FFE94E",
    x"1FFE554",
    x"1FFE15B",
    x"1FFDD64",
    x"1FFD96D",
    x"1FFD577",
    x"1FFD182",
    x"1FFCD8E",
    x"1FFC99B",
    x"1FFC5A9",
    x"1FFC1B8",
    x"1FFBDC8",
    x"1FFB9D9",
    x"1FFB5EB",
    x"1FFB1FE",
    x"1FFAE12",
    x"1FFAA27",
    x"1FFA63D",
    x"1FFA254",
    x"1FF9E6C",
    x"1FF9A85",
    x"1FF969F",
    x"1FF92BA",
    x"1FF8ED6",
    x"1FF8AF2",
    x"1FF8710",
    x"1FF832F",
    x"1FF7F4F",
    x"1FF7B6F",
    x"1FF7791",
    x"1FF73B3",
    x"1FF6FD7",
    x"1FF6BFC",
    x"1FF6821",
    x"1FF6447",
    x"1FF606F",
    x"1FF5C97",
    x"1FF58C1",
    x"1FF54EB",
    x"1FF5116",
    x"1FF4D42",
    x"1FF496F",
    x"1FF459E",
    x"1FF41CD",
    x"1FF3DFD",
    x"1FF3A2E",
    x"1FF3660",
    x"1FF3292",
    x"1FF2EC6",
    x"1FF2AFB",
    x"1FF2731",
    x"1FF2367",
    x"1FF1F9F",
    x"1FF1BD8",
    x"1FF1811",
    x"1FF144C",
    x"1FF1087",
    x"1FF0CC3",
    x"1FF0901",
    x"1FF053F",
    x"1FF017E",
    x"1FEFDBE",
    x"1FEF9FF",
    x"1FEF641",
    x"1FEF284",
    x"1FEEEC8",
    x"1FEEB0D",
    x"1FEE752",
    x"1FEE399",
    x"1FEDFE1",
    x"1FEDC29",
    x"1FED872",
    x"1FED4BD",
    x"1FED108",
    x"1FECD54",
    x"1FEC9A1",
    x"1FEC5EF",
    x"1FEC23E",
    x"1FEBE8E",
    x"1FEBADF",
    x"1FEB731",
    x"1FEB384",
    x"1FEAFD7",
    x"1FEAC2C",
    x"1FEA881",
    x"1FEA4D7",
    x"1FEA12F",
    x"1FE9D87",
    x"1FE99E0",
    x"1FE963A",
    x"1FE9295",
    x"1FE8EF1",
    x"1FE8B4D",
    x"1FE87AB",
    x"1FE8409",
    x"1FE8069",
    x"1FE7CC9",
    x"1FE792B",
    x"1FE758D",
    x"1FE71F0",
    x"1FE6E54",
    x"1FE6AB9",
    x"1FE671E",
    x"1FE6385",
    x"1FE5FED",
    x"1FE5C55",
    x"1FE58BE",
    x"1FE5529",
    x"1FE5194",
    x"1FE4E00",
    x"1FE4A6D",
    x"1FE46DB",
    x"1FE4349",
    x"1FE3FB9",
    x"1FE3C2A",
    x"1FE389B",
    x"1FE350D",
    x"1FE3180",
    x"1FE2DF4",
    x"1FE2A69",
    x"1FE26DF",
    x"1FE2356",
    x"1FE1FCE",
    x"1FE1C46",
    x"1FE18BF",
    x"1FE153A",
    x"1FE11B5",
    x"1FE0E31",
    x"1FE0AAE",
    x"1FE072C",
    x"1FE03AA",
    x"1FE002A",
    x"1FDFCAA",
    x"1FDF92B",
    x"1FDF5AE",
    x"1FDF231",
    x"1FDEEB4",
    x"1FDEB39",
    x"1FDE7BF",
    x"1FDE445",
    x"1FDE0CD",
    x"1FDDD55",
    x"1FDD9DE",
    x"1FDD668",
    x"1FDD2F3",
    x"1FDCF7E",
    x"1FDCC0B",
    x"1FDC898",
    x"1FDC527",
    x"1FDC1B6",
    x"1FDBE46",
    x"1FDBAD7",
    x"1FDB768",
    x"1FDB3FB",
    x"1FDB08E",
    x"1FDAD23",
    x"1FDA9B8",
    x"1FDA64E",
    x"1FDA2E5",
    x"1FD9F7C",
    x"1FD9C15",
    x"1FD98AE",
    x"1FD9549",
    x"1FD91E4",
    x"1FD8E80",
    x"1FD8B1D",
    x"1FD87BA",
    x"1FD8459",
    x"1FD80F8",
    x"1FD7D98",
    x"1FD7A39",
    x"1FD76DB",
    x"1FD737E",
    x"1FD7021",
    x"1FD6CC6",
    x"1FD696B",
    x"1FD6611",
    x"1FD62B8",
    x"1FD5F60",
    x"1FD5C08",
    x"1FD58B2",
    x"1FD555C",
    x"1FD5207",
    x"1FD4EB3",
    x"1FD4B60",
    x"1FD480D",
    x"1FD44BC",
    x"1FD416B",
    x"1FD3E1B",
    x"1FD3ACC",
    x"1FD377D",
    x"1FD3430",
    x"1FD30E3",
    x"1FD2D98",
    x"1FD2A4D",
    x"1FD2702",
    x"1FD23B9",
    x"1FD2071",
    x"1FD1D29",
    x"1FD19E2",
    x"1FD169C",
    x"1FD1357",
    x"1FD1012",
    x"1FD0CCF",
    x"1FD098C",
    x"1FD064A",
    x"1FD0309",
    x"1FCFFC8",
    x"1FCFC89",
    x"1FCF94A",
    x"1FCF60C",
    x"1FCF2CF",
    x"1FCEF93",
    x"1FCEC57",
    x"1FCE91D",
    x"1FCE5E3",
    x"1FCE2AA",
    x"1FCDF71",
    x"1FCDC3A",
    x"1FCD903",
    x"1FCD5CD",
    x"1FCD298",
    x"1FCCF64",
    x"1FCCC31",
    x"1FCC8FE",
    x"1FCC5CC",
    x"1FCC29B",
    x"1FCBF6B",
    x"1FCBC3B",
    x"1FCB90D",
    x"1FCB5DF",
    x"1FCB2B2",
    x"1FCAF85",
    x"1FCAC5A",
    x"1FCA92F",
    x"1FCA605",
    x"1FCA2DC",
    x"1FC9FB4",
    x"1FC9C8C",
    x"1FC9966",
    x"1FC9640",
    x"1FC931B",
    x"1FC8FF6",
    x"1FC8CD3",
    x"1FC89B0",
    x"1FC868E",
    x"1FC836D",
    x"1FC804C",
    x"1FC7D2C",
    x"1FC7A0D",
    x"1FC76EF",
    x"1FC73D2",
    x"1FC70B5",
    x"1FC6D9A",
    x"1FC6A7F",
    x"1FC6764",
    x"1FC644B",
    x"1FC6132",
    x"1FC5E1A",
    x"1FC5B03",
    x"1FC57ED",
    x"1FC54D7",
    x"1FC51C2",
    x"1FC4EAE",
    x"1FC4B9B",
    x"1FC4889",
    x"1FC4577",
    x"1FC4266",
    x"1FC3F56",
    x"1FC3C46",
    x"1FC3937",
    x"1FC362A",
    x"1FC331C",
    x"1FC3010",
    x"1FC2D04",
    x"1FC29F9",
    x"1FC26EF",
    x"1FC23E6",
    x"1FC20DD",
    x"1FC1DD6",
    x"1FC1ACE",
    x"1FC17C8",
    x"1FC14C3",
    x"1FC11BE",
    x"1FC0EBA",
    x"1FC0BB6",
    x"1FC08B4",
    x"1FC05B2",
    x"1FC02B1",
    x"1FBFFB1",
    x"1FBFCB1",
    x"1FBF9B2",
    x"1FBF6B4",
    x"1FBF3B7",
    x"1FBF0BA",
    x"1FBEDBF",
    x"1FBEAC4",
    x"1FBE7C9",
    x"1FBE4D0",
    x"1FBE1D7",
    x"1FBDEDF",
    x"1FBDBE7",
    x"1FBD8F1",
    x"1FBD5FB",
    x"1FBD306",
    x"1FBD011",
    x"1FBCD1E",
    x"1FBCA2B",
    x"1FBC739",
    x"1FBC447",
    x"1FBC157",
    x"1FBBE67",
    x"1FBBB77",
    x"1FBB889",
    x"1FBB59B",
    x"1FBB2AE",
    x"1FBAFC2",
    x"1FBACD6",
    x"1FBA9EB",
    x"1FBA701",
    x"1FBA418",
    x"1FBA12F",
    x"1FB9E47",
    x"1FB9B60",
    x"1FB987A",
    x"1FB9594",
    x"1FB92AF",
    x"1FB8FCA",
    x"1FB8CE7",
    x"1FB8A04",
    x"1FB8722",
    x"1FB8440",
    x"1FB8160",
    x"1FB7E80",
    x"1FB7BA0",
    x"1FB78C2",
    x"1FB75E4",
    x"1FB7307",
    x"1FB702B",
    x"1FB6D4F",
    x"1FB6A74",
    x"1FB679A",
    x"1FB64C0",
    x"1FB61E7",
    x"1FB5F0F",
    x"1FB5C38",
    x"1FB5961",
    x"1FB568B",
    x"1FB53B6",
    x"1FB50E1",
    x"1FB4E0D",
    x"1FB4B3A",
    x"1FB4868",
    x"1FB4596",
    x"1FB42C5",
    x"1FB3FF5",
    x"1FB3D25",
    x"1FB3A56",
    x"1FB3788",
    x"1FB34BA",
    x"1FB31ED",
    x"1FB2F21",
    x"1FB2C56",
    x"1FB298B",
    x"1FB26C1",
    x"1FB23F8",
    x"1FB212F",
    x"1FB1E67",
    x"1FB1BA0",
    x"1FB18D9",
    x"1FB1613",
    x"1FB134E",
    x"1FB108A",
    x"1FB0DC6",
    x"1FB0B03",
    x"1FB0841",
    x"1FB057F",
    x"1FB02BE",
    x"1FAFFFD",
    x"1FAFD3E",
    x"1FAFA7F",
    x"1FAF7C1",
    x"1FAF503",
    x"1FAF246",
    x"1FAEF8A",
    x"1FAECCE",
    x"1FAEA13",
    x"1FAE759",
    x"1FAE4A0",
    x"1FAE1E7",
    x"1FADF2F",
    x"1FADC77",
    x"1FAD9C1",
    x"1FAD70A",
    x"1FAD455",
    x"1FAD1A0",
    x"1FACEEC",
    x"1FACC39",
    x"1FAC986",
    x"1FAC6D4",
    x"1FAC423",
    x"1FAC172",
    x"1FABEC2",
    x"1FABC13",
    x"1FAB964",
    x"1FAB6B6",
    x"1FAB409",
    x"1FAB15C",
    x"1FAAEB0",
    x"1FAAC05",
    x"1FAA95A",
    x"1FAA6B0",
    x"1FAA407",
    x"1FAA15E",
    x"1FA9EB6",
    x"1FA9C0E",
    x"1FA9968",
    x"1FA96C2",
    x"1FA941C",
    x"1FA9178",
    x"1FA8ED4",
    x"1FA8C30",
    x"1FA898E",
    x"1FA86EC",
    x"1FA844A",
    x"1FA81A9",
    x"1FA7F09",
    x"1FA7C6A",
    x"1FA79CB",
    x"1FA772D",
    x"1FA748F",
    x"1FA71F3",
    x"1FA6F57",
    x"1FA6CBB",
    x"1FA6A20",
    x"1FA6786",
    x"1FA64EC",
    x"1FA6253",
    x"1FA5FBB",
    x"1FA5D24",
    x"1FA5A8D",
    x"1FA57F6",
    x"1FA5561",
    x"1FA52CC",
    x"1FA5037",
    x"1FA4DA4",
    x"1FA4B10",
    x"1FA487E",
    x"1FA45EC",
    x"1FA435B",
    x"1FA40CB",
    x"1FA3E3B",
    x"1FA3BAB",
    x"1FA391D",
    x"1FA368F",
    x"1FA3402",
    x"1FA3175",
    x"1FA2EE9",
    x"1FA2C5D",
    x"1FA29D3",
    x"1FA2748",
    x"1FA24BF",
    x"1FA2236",
    x"1FA1FAE",
    x"1FA1D26",
    x"1FA1A9F",
    x"1FA1819",
    x"1FA1593",
    x"1FA130E",
    x"1FA108A",
    x"1FA0E06",
    x"1FA0B83",
    x"1FA0900",
    x"1FA067E",
    x"1FA03FD",
    x"1FA017C",
    x"1F9FEFC",
    x"1F9FC7D",
    x"1F9F9FE",
    x"1F9F780",
    x"1F9F502",
    x"1F9F285",
    x"1F9F009",
    x"1F9ED8D",
    x"1F9EB12",
    x"1F9E898",
    x"1F9E61E",
    x"1F9E3A5",
    x"1F9E12C",
    x"1F9DEB4",
    x"1F9DC3D",
    x"1F9D9C6",
    x"1F9D750",
    x"1F9D4DA",
    x"1F9D265",
    x"1F9CFF1",
    x"1F9CD7D",
    x"1F9CB0A",
    x"1F9C898",
    x"1F9C626",
    x"1F9C3B5",
    x"1F9C144",
    x"1F9BED4",
    x"1F9BC65",
    x"1F9B9F6",
    x"1F9B788",
    x"1F9B51A",
    x"1F9B2AD",
    x"1F9B041",
    x"1F9ADD5",
    x"1F9AB6A",
    x"1F9A8FF",
    x"1F9A695",
    x"1F9A42C",
    x"1F9A1C3",
    x"1F99F5B",
    x"1F99CF4",
    x"1F99A8D",
    x"1F99826",
    x"1F995C1",
    x"1F9935B",
    x"1F990F7",
    x"1F98E93",
    x"1F98C30",
    x"1F989CD",
    x"1F9876B",
    x"1F98509",
    x"1F982A8",
    x"1F98048",
    x"1F97DE8",
    x"1F97B89",
    x"1F9792A",
    x"1F976CC",
    x"1F9746F",
    x"1F97212",
    x"1F96FB6",
    x"1F96D5A",
    x"1F96AFF",
    x"1F968A5",
    x"1F9664B",
    x"1F963F2",
    x"1F96199",
    x"1F95F41",
    x"1F95CE9",
    x"1F95A92",
    x"1F9583C",
    x"1F955E6",
    x"1F95391",
    x"1F9513C",
    x"1F94EE8",
    x"1F94C95",
    x"1F94A42",
    x"1F947F0",
    x"1F9459E",
    x"1F9434D",
    x"1F940FD",
    x"1F93EAD",
    x"1F93C5D",
    x"1F93A0E",
    x"1F937C0",
    x"1F93572",
    x"1F93325",
    x"1F930D9",
    x"1F92E8D",
    x"1F92C42",
    x"1F929F7",
    x"1F927AD",
    x"1F92563",
    x"1F9231A",
    x"1F920D1",
    x"1F91E8A",
    x"1F91C42",
    x"1F919FB",
    x"1F917B5",
    x"1F91570",
    x"1F9132A",
    x"1F910E6",
    x"1F90EA2",
    x"1F90C5F",
    x"1F90A1C",
    x"1F907DA",
    x"1F90598",
    x"1F90357",
    x"1F90116",
    x"1F8FED6",
    x"1F8FC97",
    x"1F8FA58",
    x"1F8F81A",
    x"1F8F5DC",
    x"1F8F39F",
    x"1F8F162",
    x"1F8EF26",
    x"1F8ECEB",
    x"1F8EAB0",
    x"1F8E875",
    x"1F8E63B",
    x"1F8E402",
    x"1F8E1C9",
    x"1F8DF91",
    x"1F8DD5A",
    x"1F8DB23",
    x"1F8D8EC",
    x"1F8D6B6",
    x"1F8D481",
    x"1F8D24C",
    x"1F8D017",
    x"1F8CDE4",
    x"1F8CBB1",
    x"1F8C97E",
    x"1F8C74C",
    x"1F8C51A",
    x"1F8C2E9",
    x"1F8C0B9",
    x"1F8BE89",
    x"1F8BC5A",
    x"1F8BA2B",
    x"1F8B7FC",
    x"1F8B5CF",
    x"1F8B3A2",
    x"1F8B175",
    x"1F8AF49",
    x"1F8AD1D",
    x"1F8AAF2",
    x"1F8A8C8",
    x"1F8A69E",
    x"1F8A474",
    x"1F8A24C",
    x"1F8A023",
    x"1F89DFC",
    x"1F89BD4",
    x"1F899AE",
    x"1F89787",
    x"1F89562",
    x"1F8933D",
    x"1F89118",
    x"1F88EF4",
    x"1F88CD1",
    x"1F88AAE",
    x"1F8888B",
    x"1F8866A",
    x"1F88448",
    x"1F88227",
    x"1F88007",
    x"1F87DE7",
    x"1F87BC8",
    x"1F879AA",
    x"1F8778B",
    x"1F8756E",
    x"1F87351",
    x"1F87134",
    x"1F86F18",
    x"1F86CFD",
    x"1F86AE2",
    x"1F868C7",
    x"1F866AD",
    x"1F86494",
    x"1F8627B",
    x"1F86063",
    x"1F85E4B",
    x"1F85C33",
    x"1F85A1D",
    x"1F85806",
    x"1F855F1",
    x"1F853DB",
    x"1F851C7",
    x"1F84FB2",
    x"1F84D9F",
    x"1F84B8C",
    x"1F84979",
    x"1F84767",
    x"1F84555",
    x"1F84344",
    x"1F84134",
    x"1F83F24",
    x"1F83D14",
    x"1F83B05",
    x"1F838F7",
    x"1F836E9",
    x"1F834DB",
    x"1F832CE",
    x"1F830C2",
    x"1F82EB6",
    x"1F82CAA",
    x"1F82A9F",
    x"1F82895",
    x"1F8268B",
    x"1F82482",
    x"1F82279",
    x"1F82071",
    x"1F81E69",
    x"1F81C61",
    x"1F81A5B",
    x"1F81854",
    x"1F8164E",
    x"1F81449",
    x"1F81244",
    x"1F81040",
    x"1F80E3C",
    x"1F80C39",
    x"1F80A36",
    x"1F80834",
    x"1F80632",
    x"1F80431",
    x"1F80230",
    x"1F8002F",
    x"1F7FC60",
    x"1F7F861",
    x"1F7F464",
    x"1F7F067",
    x"1F7EC6B",
    x"1F7E871",
    x"1F7E477",
    x"1F7E07F",
    x"1F7DC87",
    x"1F7D890",
    x"1F7D49B",
    x"1F7D0A6",
    x"1F7CCB2",
    x"1F7C8C0",
    x"1F7C4CE",
    x"1F7C0DD",
    x"1F7BCEE",
    x"1F7B8FF",
    x"1F7B511",
    x"1F7B124",
    x"1F7AD38",
    x"1F7A94E",
    x"1F7A564",
    x"1F7A17B",
    x"1F79D93",
    x"1F799AC",
    x"1F795C6",
    x"1F791E1",
    x"1F78DFD",
    x"1F78A1A",
    x"1F78638",
    x"1F78257",
    x"1F77E77",
    x"1F77A98",
    x"1F776BA",
    x"1F772DD",
    x"1F76F00",
    x"1F76B25",
    x"1F7674B",
    x"1F76371",
    x"1F75F99",
    x"1F75BC2",
    x"1F757EB",
    x"1F75416",
    x"1F75041",
    x"1F74C6E",
    x"1F7489B",
    x"1F744C9",
    x"1F740F9",
    x"1F73D29",
    x"1F7395A",
    x"1F7358C",
    x"1F731BF",
    x"1F72DF3",
    x"1F72A28",
    x"1F7265E",
    x"1F72295",
    x"1F71ECD",
    x"1F71B06",
    x"1F7173F",
    x"1F7137A",
    x"1F70FB6",
    x"1F70BF2",
    x"1F70830",
    x"1F7046E",
    x"1F700AD",
    x"1F6FCEE",
    x"1F6F92F",
    x"1F6F571",
    x"1F6F1B4",
    x"1F6EDF8",
    x"1F6EA3D",
    x"1F6E683",
    x"1F6E2CA",
    x"1F6DF12",
    x"1F6DB5A",
    x"1F6D7A4",
    x"1F6D3EF",
    x"1F6D03A",
    x"1F6CC86",
    x"1F6C8D4",
    x"1F6C522",
    x"1F6C171",
    x"1F6BDC1",
    x"1F6BA12",
    x"1F6B664",
    x"1F6B2B7",
    x"1F6AF0B",
    x"1F6AB60",
    x"1F6A7B5",
    x"1F6A40C",
    x"1F6A063",
    x"1F69CBC",
    x"1F69915",
    x"1F6956F",
    x"1F691CA",
    x"1F68E26",
    x"1F68A83",
    x"1F686E1",
    x"1F68340",
    x"1F67F9F",
    x"1F67C00",
    x"1F67861",
    x"1F674C4",
    x"1F67127",
    x"1F66D8B",
    x"1F669F0",
    x"1F66656",
    x"1F662BD",
    x"1F65F25",
    x"1F65B8D",
    x"1F657F7",
    x"1F65461",
    x"1F650CD",
    x"1F64D39",
    x"1F649A6",
    x"1F64614",
    x"1F64283",
    x"1F63EF3",
    x"1F63B64",
    x"1F637D5",
    x"1F63448",
    x"1F630BB",
    x"1F62D2F",
    x"1F629A4",
    x"1F6261A",
    x"1F62291",
    x"1F61F09",
    x"1F61B82",
    x"1F617FB",
    x"1F61476",
    x"1F610F1",
    x"1F60D6D",
    x"1F609EB",
    x"1F60668",
    x"1F602E7",
    x"1F5FF67",
    x"1F5FBE8",
    x"1F5F869",
    x"1F5F4EB",
    x"1F5F16F",
    x"1F5EDF3",
    x"1F5EA78",
    x"1F5E6FD",
    x"1F5E384",
    x"1F5E00C",
    x"1F5DC94",
    x"1F5D91D",
    x"1F5D5A8",
    x"1F5D233",
    x"1F5CEBE",
    x"1F5CB4B",
    x"1F5C7D9",
    x"1F5C467",
    x"1F5C0F7",
    x"1F5BD87",
    x"1F5BA18",
    x"1F5B6AA",
    x"1F5B33D",
    x"1F5AFD0",
    x"1F5AC65",
    x"1F5A8FA",
    x"1F5A590",
    x"1F5A227",
    x"1F59EBF",
    x"1F59B58",
    x"1F597F1",
    x"1F5948C",
    x"1F59127",
    x"1F58DC3",
    x"1F58A60",
    x"1F586FE",
    x"1F5839D",
    x"1F5803C",
    x"1F57CDD",
    x"1F5797E",
    x"1F57620",
    x"1F572C3",
    x"1F56F66",
    x"1F56C0B",
    x"1F568B0",
    x"1F56557",
    x"1F561FE",
    x"1F55EA6",
    x"1F55B4E",
    x"1F557F8",
    x"1F554A2",
    x"1F5514E",
    x"1F54DFA",
    x"1F54AA7",
    x"1F54754",
    x"1F54403",
    x"1F540B2",
    x"1F53D63",
    x"1F53A14",
    x"1F536C6",
    x"1F53378",
    x"1F5302C",
    x"1F52CE0",
    x"1F52995",
    x"1F5264C",
    x"1F52302",
    x"1F51FBA",
    x"1F51C72",
    x"1F5192C",
    x"1F515E6",
    x"1F512A1",
    x"1F50F5D",
    x"1F50C19",
    x"1F508D7",
    x"1F50595",
    x"1F50254",
    x"1F4FF14",
    x"1F4FBD4",
    x"1F4F896",
    x"1F4F558",
    x"1F4F21B",
    x"1F4EEDF",
    x"1F4EBA4",
    x"1F4E869",
    x"1F4E52F",
    x"1F4E1F6",
    x"1F4DEBE",
    x"1F4DB87",
    x"1F4D851",
    x"1F4D51B",
    x"1F4D1E6",
    x"1F4CEB2",
    x"1F4CB7F",
    x"1F4C84C",
    x"1F4C51B",
    x"1F4C1EA",
    x"1F4BEBA",
    x"1F4BB8A",
    x"1F4B85C",
    x"1F4B52E",
    x"1F4B201",
    x"1F4AED5",
    x"1F4ABAA",
    x"1F4A87F",
    x"1F4A556",
    x"1F4A22D",
    x"1F49F04",
    x"1F49BDD",
    x"1F498B7",
    x"1F49591",
    x"1F4926C",
    x"1F48F48",
    x"1F48C24",
    x"1F48901",
    x"1F485E0",
    x"1F482BF",
    x"1F47F9E",
    x"1F47C7F",
    x"1F47960",
    x"1F47642",
    x"1F47325",
    x"1F47008",
    x"1F46CED",
    x"1F469D2",
    x"1F466B8",
    x"1F4639F",
    x"1F46086",
    x"1F45D6E",
    x"1F45A57",
    x"1F45741",
    x"1F4542C",
    x"1F45117",
    x"1F44E03",
    x"1F44AF0",
    x"1F447DE",
    x"1F444CC",
    x"1F441BB",
    x"1F43EAB",
    x"1F43B9C",
    x"1F4388D",
    x"1F43580",
    x"1F43273",
    x"1F42F66",
    x"1F42C5B",
    x"1F42950",
    x"1F42646",
    x"1F4233D",
    x"1F42035",
    x"1F41D2D",
    x"1F41A26",
    x"1F41720",
    x"1F4141B",
    x"1F41116",
    x"1F40E12",
    x"1F40B0F",
    x"1F4080D",
    x"1F4050B",
    x"1F4020A",
    x"1F3FF0A",
    x"1F3FC0A",
    x"1F3F90C",
    x"1F3F60E",
    x"1F3F311",
    x"1F3F014",
    x"1F3ED19",
    x"1F3EA1E",
    x"1F3E724",
    x"1F3E42A",
    x"1F3E132",
    x"1F3DE3A",
    x"1F3DB43",
    x"1F3D84C",
    x"1F3D556",
    x"1F3D261",
    x"1F3CF6D",
    x"1F3CC7A",
    x"1F3C987",
    x"1F3C695",
    x"1F3C3A4",
    x"1F3C0B3",
    x"1F3BDC3",
    x"1F3BAD4",
    x"1F3B7E6",
    x"1F3B4F8",
    x"1F3B20B",
    x"1F3AF1F",
    x"1F3AC34",
    x"1F3A949",
    x"1F3A65F",
    x"1F3A376",
    x"1F3A08D",
    x"1F39DA6",
    x"1F39ABF",
    x"1F397D8",
    x"1F394F3",
    x"1F3920E",
    x"1F38F2A",
    x"1F38C46",
    x"1F38964",
    x"1F38682",
    x"1F383A0",
    x"1F380C0",
    x"1F37DE0",
    x"1F37B01",
    x"1F37822",
    x"1F37545",
    x"1F37268",
    x"1F36F8C",
    x"1F36CB0",
    x"1F369D5",
    x"1F366FB",
    x"1F36422",
    x"1F36149",
    x"1F35E71",
    x"1F35B9A",
    x"1F358C3",
    x"1F355ED",
    x"1F35318",
    x"1F35044",
    x"1F34D70",
    x"1F34A9D",
    x"1F347CB",
    x"1F344F9",
    x"1F34228",
    x"1F33F58",
    x"1F33C89",
    x"1F339BA",
    x"1F336EC",
    x"1F3341E",
    x"1F33152",
    x"1F32E86",
    x"1F32BBA",
    x"1F328F0",
    x"1F32626",
    x"1F3235D",
    x"1F32094",
    x"1F31DCD",
    x"1F31B05",
    x"1F3183F",
    x"1F31579",
    x"1F312B4",
    x"1F30FF0",
    x"1F30D2C",
    x"1F30A69",
    x"1F307A7",
    x"1F304E6",
    x"1F30225",
    x"1F2FF64",
    x"1F2FCA5",
    x"1F2F9E6",
    x"1F2F728",
    x"1F2F46B",
    x"1F2F1AE",
    x"1F2EEF2",
    x"1F2EC36",
    x"1F2E97C",
    x"1F2E6C2",
    x"1F2E408",
    x"1F2E150",
    x"1F2DE98",
    x"1F2DBE0",
    x"1F2D92A",
    x"1F2D674",
    x"1F2D3BE",
    x"1F2D10A",
    x"1F2CE56",
    x"1F2CBA3",
    x"1F2C8F0",
    x"1F2C63E",
    x"1F2C38D",
    x"1F2C0DC",
    x"1F2BE2D",
    x"1F2BB7D",
    x"1F2B8CF",
    x"1F2B621",
    x"1F2B374",
    x"1F2B0C7",
    x"1F2AE1B",
    x"1F2AB70",
    x"1F2A8C6",
    x"1F2A61C",
    x"1F2A373",
    x"1F2A0CA",
    x"1F29E22",
    x"1F29B7B",
    x"1F298D4",
    x"1F2962F",
    x"1F29389",
    x"1F290E5",
    x"1F28E41",
    x"1F28B9E",
    x"1F288FB",
    x"1F28659",
    x"1F283B8",
    x"1F28117",
    x"1F27E77",
    x"1F27BD8",
    x"1F27939",
    x"1F2769B",
    x"1F273FE",
    x"1F27161",
    x"1F26EC5",
    x"1F26C2A",
    x"1F2698F",
    x"1F266F5",
    x"1F2645C",
    x"1F261C3",
    x"1F25F2B",
    x"1F25C94",
    x"1F259FD",
    x"1F25767",
    x"1F254D1",
    x"1F2523C",
    x"1F24FA8",
    x"1F24D14",
    x"1F24A81",
    x"1F247EF",
    x"1F2455D",
    x"1F242CC",
    x"1F2403C",
    x"1F23DAC",
    x"1F23B1D",
    x"1F2388F",
    x"1F23601",
    x"1F23374",
    x"1F230E7",
    x"1F22E5B",
    x"1F22BD0",
    x"1F22945",
    x"1F226BB",
    x"1F22432",
    x"1F221A9",
    x"1F21F21",
    x"1F21C9A",
    x"1F21A13",
    x"1F2178D",
    x"1F21507",
    x"1F21282",
    x"1F20FFE",
    x"1F20D7A",
    x"1F20AF7",
    x"1F20875",
    x"1F205F3",
    x"1F20372",
    x"1F200F1",
    x"1F1FE71",
    x"1F1FBF2",
    x"1F1F973",
    x"1F1F6F5",
    x"1F1F478",
    x"1F1F1FB",
    x"1F1EF7F",
    x"1F1ED03",
    x"1F1EA88",
    x"1F1E80E",
    x"1F1E594",
    x"1F1E31B",
    x"1F1E0A3",
    x"1F1DE2B",
    x"1F1DBB4",
    x"1F1D93D",
    x"1F1D6C7",
    x"1F1D452",
    x"1F1D1DD",
    x"1F1CF69",
    x"1F1CCF5",
    x"1F1CA82",
    x"1F1C810",
    x"1F1C59E",
    x"1F1C32D",
    x"1F1C0BC",
    x"1F1BE4D",
    x"1F1BBDD",
    x"1F1B96F",
    x"1F1B701",
    x"1F1B493",
    x"1F1B226",
    x"1F1AFBA",
    x"1F1AD4E",
    x"1F1AAE3",
    x"1F1A879",
    x"1F1A60F",
    x"1F1A3A6",
    x"1F1A13D",
    x"1F19ED5",
    x"1F19C6E",
    x"1F19A07",
    x"1F197A1",
    x"1F1953B",
    x"1F192D6",
    x"1F19072",
    x"1F18E0E",
    x"1F18BAB",
    x"1F18948",
    x"1F186E6",
    x"1F18485",
    x"1F18224",
    x"1F17FC4",
    x"1F17D64",
    x"1F17B05",
    x"1F178A7",
    x"1F17649",
    x"1F173EB",
    x"1F1718F",
    x"1F16F33",
    x"1F16CD7",
    x"1F16A7C",
    x"1F16822",
    x"1F165C8",
    x"1F1636F",
    x"1F16116",
    x"1F15EBE",
    x"1F15C67",
    x"1F15A10",
    x"1F157BA",
    x"1F15564",
    x"1F1530F",
    x"1F150BB",
    x"1F14E67",
    x"1F14C14",
    x"1F149C1",
    x"1F1476F",
    x"1F1451D",
    x"1F142CC",
    x"1F1407C",
    x"1F13E2C",
    x"1F13BDD",
    x"1F1398E",
    x"1F13740",
    x"1F134F2",
    x"1F132A6",
    x"1F13059",
    x"1F12E0D",
    x"1F12BC2",
    x"1F12977",
    x"1F1272D",
    x"1F124E4",
    x"1F1229B",
    x"1F12053",
    x"1F11E0B",
    x"1F11BC4",
    x"1F1197D",
    x"1F11737",
    x"1F114F1",
    x"1F112AC",
    x"1F11068",
    x"1F10E24",
    x"1F10BE1",
    x"1F1099E",
    x"1F1075C",
    x"1F1051A",
    x"1F102D9",
    x"1F10099",
    x"1F0FE59",
    x"1F0FC1A",
    x"1F0F9DB",
    x"1F0F79D",
    x"1F0F55F",
    x"1F0F322",
    x"1F0F0E6",
    x"1F0EEAA",
    x"1F0EC6E",
    x"1F0EA34",
    x"1F0E7F9",
    x"1F0E5C0",
    x"1F0E386",
    x"1F0E14E",
    x"1F0DF16",
    x"1F0DCDE",
    x"1F0DAA7",
    x"1F0D871",
    x"1F0D63B",
    x"1F0D406",
    x"1F0D1D1",
    x"1F0CF9D",
    x"1F0CD69",
    x"1F0CB36",
    x"1F0C904",
    x"1F0C6D2",
    x"1F0C4A0",
    x"1F0C26F",
    x"1F0C03F",
    x"1F0BE0F",
    x"1F0BBE0",
    x"1F0B9B1",
    x"1F0B783",
    x"1F0B556",
    x"1F0B329",
    x"1F0B0FC",
    x"1F0AED0",
    x"1F0ACA5",
    x"1F0AA7A",
    x"1F0A84F",
    x"1F0A626",
    x"1F0A3FC",
    x"1F0A1D4",
    x"1F09FAB",
    x"1F09D84",
    x"1F09B5D",
    x"1F09936",
    x"1F09710",
    x"1F094EB",
    x"1F092C6",
    x"1F090A1",
    x"1F08E7D",
    x"1F08C5A",
    x"1F08A37",
    x"1F08815",
    x"1F085F3",
    x"1F083D2",
    x"1F081B1",
    x"1F07F91",
    x"1F07D71",
    x"1F07B52",
    x"1F07934",
    x"1F07716",
    x"1F074F8",
    x"1F072DB",
    x"1F070BF",
    x"1F06EA3",
    x"1F06C87",
    x"1F06A6D",
    x"1F06852",
    x"1F06638",
    x"1F0641F",
    x"1F06206",
    x"1F05FEE",
    x"1F05DD6",
    x"1F05BBF",
    x"1F059A8",
    x"1F05792",
    x"1F0557D",
    x"1F05368",
    x"1F05153",
    x"1F04F3F",
    x"1F04D2B",
    x"1F04B18",
    x"1F04906",
    x"1F046F4",
    x"1F044E2",
    x"1F042D1",
    x"1F040C1",
    x"1F03EB1",
    x"1F03CA2",
    x"1F03A93",
    x"1F03884",
    x"1F03676",
    x"1F03469",
    x"1F0325C",
    x"1F03050",
    x"1F02E44",
    x"1F02C39",
    x"1F02A2E",
    x"1F02824",
    x"1F0261A",
    x"1F02411",
    x"1F02208",
    x"1F02000",
    x"1F01DF8",
    x"1F01BF1",
    x"1F019EA",
    x"1F017E4",
    x"1F015DE",
    x"1F013D9",
    x"1F011D4",
    x"1F00FD0",
    x"1F00DCC",
    x"1F00BC9",
    x"1F009C6",
    x"1F007C4",
    x"1F005C2",
    x"1F003C1",
    x"1F001C0",
    x"1EFFF81",
    x"1EFFB82",
    x"1EFF783",
    x"1EFF386",
    x"1EFEF89",
    x"1EFEB8E",
    x"1EFE794",
    x"1EFE39A",
    x"1EFDFA2",
    x"1EFDBAA",
    x"1EFD7B4",
    x"1EFD3BF",
    x"1EFCFCA",
    x"1EFCBD7",
    x"1EFC7E4",
    x"1EFC3F3",
    x"1EFC002",
    x"1EFBC13",
    x"1EFB824",
    x"1EFB437",
    x"1EFB04A",
    x"1EFAC5E",
    x"1EFA874",
    x"1EFA48A",
    x"1EFA0A2",
    x"1EF9CBA",
    x"1EF98D3",
    x"1EF94EE",
    x"1EF9109",
    x"1EF8D25",
    x"1EF8942",
    x"1EF8560",
    x"1EF8180",
    x"1EF7DA0",
    x"1EF79C1",
    x"1EF75E3",
    x"1EF7206",
    x"1EF6E2A",
    x"1EF6A4F",
    x"1EF6675",
    x"1EF629B",
    x"1EF5EC3",
    x"1EF5AEC",
    x"1EF5716",
    x"1EF5341",
    x"1EF4F6C",
    x"1EF4B99",
    x"1EF47C6",
    x"1EF43F5",
    x"1EF4024",
    x"1EF3C55",
    x"1EF3886",
    x"1EF34B9",
    x"1EF30EC",
    x"1EF2D20",
    x"1EF2955",
    x"1EF258B",
    x"1EF21C3",
    x"1EF1DFB",
    x"1EF1A34",
    x"1EF166D",
    x"1EF12A8",
    x"1EF0EE4",
    x"1EF0B21",
    x"1EF075F",
    x"1EF039D",
    x"1EEFFDD",
    x"1EEFC1D",
    x"1EEF85F",
    x"1EEF4A1",
    x"1EEF0E4",
    x"1EEED29",
    x"1EEE96E",
    x"1EEE5B4",
    x"1EEE1FB",
    x"1EEDE43",
    x"1EEDA8C",
    x"1EED6D6",
    x"1EED320",
    x"1EECF6C",
    x"1EECBB9",
    x"1EEC806",
    x"1EEC455",
    x"1EEC0A4",
    x"1EEBCF4",
    x"1EEB946",
    x"1EEB598",
    x"1EEB1EB",
    x"1EEAE3F",
    x"1EEAA94",
    x"1EEA6E9",
    x"1EEA340",
    x"1EE9F98",
    x"1EE9BF0",
    x"1EE984A",
    x"1EE94A4",
    x"1EE9100",
    x"1EE8D5C",
    x"1EE89B9",
    x"1EE8617",
    x"1EE8276",
    x"1EE7ED6",
    x"1EE7B36",
    x"1EE7798",
    x"1EE73FB",
    x"1EE705E",
    x"1EE6CC2",
    x"1EE6928",
    x"1EE658E",
    x"1EE61F5",
    x"1EE5E5D",
    x"1EE5AC6",
    x"1EE572F",
    x"1EE539A",
    x"1EE5006",
    x"1EE4C72",
    x"1EE48DF",
    x"1EE454E",
    x"1EE41BD",
    x"1EE3E2D",
    x"1EE3A9E",
    x"1EE3710",
    x"1EE3382",
    x"1EE2FF6",
    x"1EE2C6A",
    x"1EE28E0",
    x"1EE2556",
    x"1EE21CD",
    x"1EE1E45",
    x"1EE1ABE",
    x"1EE1737",
    x"1EE13B2",
    x"1EE102E",
    x"1EE0CAA",
    x"1EE0927",
    x"1EE05A5",
    x"1EE0224",
    x"1EDFEA4",
    x"1EDFB25",
    x"1EDF7A7",
    x"1EDF429",
    x"1EDF0AD",
    x"1EDED31",
    x"1EDE9B6",
    x"1EDE63C",
    x"1EDE2C3",
    x"1EDDF4B",
    x"1EDDBD3",
    x"1EDD85D",
    x"1EDD4E7",
    x"1EDD172",
    x"1EDCDFE",
    x"1EDCA8B",
    x"1EDC719",
    x"1EDC3A8",
    x"1EDC037",
    x"1EDBCC8",
    x"1EDB959",
    x"1EDB5EB",
    x"1EDB27E",
    x"1EDAF12",
    x"1EDABA6",
    x"1EDA83C",
    x"1EDA4D2",
    x"1EDA16A",
    x"1ED9E02",
    x"1ED9A9B",
    x"1ED9734",
    x"1ED93CF",
    x"1ED906A",
    x"1ED8D07",
    x"1ED89A4",
    x"1ED8642",
    x"1ED82E1",
    x"1ED7F80",
    x"1ED7C21",
    x"1ED78C2",
    x"1ED7565",
    x"1ED7208",
    x"1ED6EAC",
    x"1ED6B50",
    x"1ED67F6",
    x"1ED649C",
    x"1ED6144",
    x"1ED5DEC",
    x"1ED5A95",
    x"1ED573E",
    x"1ED53E9",
    x"1ED5095",
    x"1ED4D41",
    x"1ED49EE",
    x"1ED469C",
    x"1ED434B",
    x"1ED3FFA",
    x"1ED3CAB",
    x"1ED395C",
    x"1ED360E",
    x"1ED32C1",
    x"1ED2F75",
    x"1ED2C29",
    x"1ED28DE",
    x"1ED2595",
    x"1ED224C",
    x"1ED1F04",
    x"1ED1BBC",
    x"1ED1876",
    x"1ED1530",
    x"1ED11EB",
    x"1ED0EA7",
    x"1ED0B64",
    x"1ED0821",
    x"1ED04E0",
    x"1ED019F",
    x"1ECFE5F",
    x"1ECFB20",
    x"1ECF7E1",
    x"1ECF4A4",
    x"1ECF167",
    x"1ECEE2B",
    x"1ECEAF0",
    x"1ECE7B6",
    x"1ECE47C",
    x"1ECE143",
    x"1ECDE0B",
    x"1ECDAD4",
    x"1ECD79E",
    x"1ECD468",
    x"1ECD134",
    x"1ECCE00",
    x"1ECCACD",
    x"1ECC79A",
    x"1ECC469",
    x"1ECC138",
    x"1ECBE08",
    x"1ECBAD9",
    x"1ECB7AB",
    x"1ECB47D",
    x"1ECB151",
    x"1ECAE25",
    x"1ECAAFA",
    x"1ECA7CF",
    x"1ECA4A6",
    x"1ECA17D",
    x"1EC9E55",
    x"1EC9B2E",
    x"1EC9807",
    x"1EC94E2",
    x"1EC91BD",
    x"1EC8E99",
    x"1EC8B76",
    x"1EC8853",
    x"1EC8531",
    x"1EC8211",
    x"1EC7EF0",
    x"1EC7BD1",
    x"1EC78B3",
    x"1EC7595",
    x"1EC7278",
    x"1EC6F5B",
    x"1EC6C40",
    x"1EC6925",
    x"1EC660B",
    x"1EC62F2",
    x"1EC5FDA",
    x"1EC5CC2",
    x"1EC59AC",
    x"1EC5696",
    x"1EC5380",
    x"1EC506C",
    x"1EC4D58",
    x"1EC4A45",
    x"1EC4733",
    x"1EC4422",
    x"1EC4111",
    x"1EC3E01",
    x"1EC3AF2",
    x"1EC37E4",
    x"1EC34D6",
    x"1EC31C9",
    x"1EC2EBD",
    x"1EC2BB2",
    x"1EC28A7",
    x"1EC259D",
    x"1EC2294",
    x"1EC1F8C",
    x"1EC1C85",
    x"1EC197E",
    x"1EC1678",
    x"1EC1373",
    x"1EC106E",
    x"1EC0D6A",
    x"1EC0A67",
    x"1EC0765",
    x"1EC0464",
    x"1EC0163",
    x"1EBFE63",
    x"1EBFB64",
    x"1EBF865",
    x"1EBF568",
    x"1EBF26B",
    x"1EBEF6E",
    x"1EBEC73",
    x"1EBE978",
    x"1EBE67E",
    x"1EBE385",
    x"1EBE08C",
    x"1EBDD95",
    x"1EBDA9E",
    x"1EBD7A7",
    x"1EBD4B2",
    x"1EBD1BD",
    x"1EBCEC9",
    x"1EBCBD6",
    x"1EBC8E3",
    x"1EBC5F1",
    x"1EBC300",
    x"1EBC010",
    x"1EBBD20",
    x"1EBBA31",
    x"1EBB743",
    x"1EBB455",
    x"1EBB169",
    x"1EBAE7D",
    x"1EBAB92",
    x"1EBA8A7",
    x"1EBA5BD",
    x"1EBA2D4",
    x"1EB9FEC",
    x"1EB9D04",
    x"1EB9A1D",
    x"1EB9737",
    x"1EB9452",
    x"1EB916D",
    x"1EB8E89",
    x"1EB8BA6",
    x"1EB88C3",
    x"1EB85E1",
    x"1EB8300",
    x"1EB8020",
    x"1EB7D40",
    x"1EB7A61",
    x"1EB7783",
    x"1EB74A5",
    x"1EB71C9",
    x"1EB6EED",
    x"1EB6C11",
    x"1EB6936",
    x"1EB665D",
    x"1EB6383",
    x"1EB60AB",
    x"1EB5DD3",
    x"1EB5AFC",
    x"1EB5825",
    x"1EB5550",
    x"1EB527B",
    x"1EB4FA7",
    x"1EB4CD3",
    x"1EB4A00",
    x"1EB472E",
    x"1EB445D",
    x"1EB418C",
    x"1EB3EBC",
    x"1EB3BEC",
    x"1EB391E",
    x"1EB3650",
    x"1EB3383",
    x"1EB30B6",
    x"1EB2DEA",
    x"1EB2B1F",
    x"1EB2855",
    x"1EB258B",
    x"1EB22C2",
    x"1EB1FFA",
    x"1EB1D32",
    x"1EB1A6B",
    x"1EB17A5",
    x"1EB14DF",
    x"1EB121A",
    x"1EB0F56",
    x"1EB0C93",
    x"1EB09D0",
    x"1EB070E",
    x"1EB044C",
    x"1EB018C",
    x"1EAFECC",
    x"1EAFC0C",
    x"1EAF94E",
    x"1EAF690",
    x"1EAF3D2",
    x"1EAF116",
    x"1EAEE5A",
    x"1EAEB9E",
    x"1EAE8E4",
    x"1EAE62A",
    x"1EAE371",
    x"1EAE0B8",
    x"1EADE00",
    x"1EADB49",
    x"1EAD893",
    x"1EAD5DD",
    x"1EAD328",
    x"1EAD073",
    x"1EACDC0",
    x"1EACB0D",
    x"1EAC85A",
    x"1EAC5A8",
    x"1EAC2F7",
    x"1EAC047",
    x"1EABD97",
    x"1EABAE8",
    x"1EAB83A",
    x"1EAB58C",
    x"1EAB2DF",
    x"1EAB033",
    x"1EAAD87",
    x"1EAAADC",
    x"1EAA831",
    x"1EAA588",
    x"1EAA2DF",
    x"1EAA036",
    x"1EA9D8F",
    x"1EA9AE7",
    x"1EA9841",
    x"1EA959B",
    x"1EA92F6",
    x"1EA9052",
    x"1EA8DAE",
    x"1EA8B0B",
    x"1EA8869",
    x"1EA85C7",
    x"1EA8326",
    x"1EA8085",
    x"1EA7DE5",
    x"1EA7B46",
    x"1EA78A8",
    x"1EA760A",
    x"1EA736D",
    x"1EA70D0",
    x"1EA6E34",
    x"1EA6B99",
    x"1EA68FF",
    x"1EA6665",
    x"1EA63CB",
    x"1EA6133",
    x"1EA5E9B",
    x"1EA5C03",
    x"1EA596D",
    x"1EA56D7",
    x"1EA5441",
    x"1EA51AD",
    x"1EA4F18",
    x"1EA4C85",
    x"1EA49F2",
    x"1EA4760",
    x"1EA44CF",
    x"1EA423E",
    x"1EA3FAD",
    x"1EA3D1E",
    x"1EA3A8F",
    x"1EA3801",
    x"1EA3573",
    x"1EA32E6",
    x"1EA3059",
    x"1EA2DCE",
    x"1EA2B43",
    x"1EA28B8",
    x"1EA262E",
    x"1EA23A5",
    x"1EA211C",
    x"1EA1E94",
    x"1EA1C0D",
    x"1EA1986",
    x"1EA1700",
    x"1EA147B",
    x"1EA11F6",
    x"1EA0F72",
    x"1EA0CEE",
    x"1EA0A6B",
    x"1EA07E9",
    x"1EA0567",
    x"1EA02E6",
    x"1EA0066",
    x"1E9FDE6",
    x"1E9FB67",
    x"1E9F8E8",
    x"1E9F66B",
    x"1E9F3ED",
    x"1E9F171",
    x"1E9EEF5",
    x"1E9EC79",
    x"1E9E9FE",
    x"1E9E784",
    x"1E9E50B",
    x"1E9E292",
    x"1E9E019",
    x"1E9DDA2",
    x"1E9DB2A",
    x"1E9D8B4",
    x"1E9D63E",
    x"1E9D3C9",
    x"1E9D154",
    x"1E9CEE0",
    x"1E9CC6D",
    x"1E9C9FA",
    x"1E9C788",
    x"1E9C516",
    x"1E9C2A5",
    x"1E9C035",
    x"1E9BDC5",
    x"1E9BB56",
    x"1E9B8E7",
    x"1E9B67A",
    x"1E9B40C",
    x"1E9B1A0",
    x"1E9AF33",
    x"1E9ACC8",
    x"1E9AA5D",
    x"1E9A7F3",
    x"1E9A589",
    x"1E9A320",
    x"1E9A0B7",
    x"1E99E50",
    x"1E99BE8",
    x"1E99982",
    x"1E9971C",
    x"1E994B6",
    x"1E99251",
    x"1E98FED",
    x"1E98D89",
    x"1E98B26",
    x"1E988C4",
    x"1E98662",
    x"1E98400",
    x"1E981A0",
    x"1E97F40",
    x"1E97CE0",
    x"1E97A81",
    x"1E97823",
    x"1E975C5",
    x"1E97368",
    x"1E9710B",
    x"1E96EAF",
    x"1E96C54",
    x"1E969F9",
    x"1E9679F",
    x"1E96546",
    x"1E962EC",
    x"1E96094",
    x"1E95E3C",
    x"1E95BE5",
    x"1E9598E",
    x"1E95738",
    x"1E954E3",
    x"1E9528E",
    x"1E95039",
    x"1E94DE6",
    x"1E94B92",
    x"1E94940",
    x"1E946EE",
    x"1E9449C",
    x"1E9424B",
    x"1E93FFB",
    x"1E93DAB",
    x"1E93B5C",
    x"1E9390E",
    x"1E936C0",
    x"1E93472",
    x"1E93226",
    x"1E92FD9",
    x"1E92D8E",
    x"1E92B43",
    x"1E928F8",
    x"1E926AE",
    x"1E92465",
    x"1E9221C",
    x"1E91FD4",
    x"1E91D8C",
    x"1E91B45",
    x"1E918FE",
    x"1E916B8",
    x"1E91473",
    x"1E9122E",
    x"1E90FEA",
    x"1E90DA6",
    x"1E90B63",
    x"1E90921",
    x"1E906DF",
    x"1E9049D",
    x"1E9025C",
    x"1E9001C",
    x"1E8FDDC",
    x"1E8FB9D",
    x"1E8F95E",
    x"1E8F720",
    x"1E8F4E3",
    x"1E8F2A6",
    x"1E8F069",
    x"1E8EE2E",
    x"1E8EBF2",
    x"1E8E9B8",
    x"1E8E77D",
    x"1E8E544",
    x"1E8E30B",
    x"1E8E0D2",
    x"1E8DE9A",
    x"1E8DC63",
    x"1E8DA2C",
    x"1E8D7F6",
    x"1E8D5C0",
    x"1E8D38B",
    x"1E8D156",
    x"1E8CF22",
    x"1E8CCEF",
    x"1E8CABC",
    x"1E8C88A",
    x"1E8C658",
    x"1E8C426",
    x"1E8C1F6",
    x"1E8BFC5",
    x"1E8BD96",
    x"1E8BB67",
    x"1E8B938",
    x"1E8B70A",
    x"1E8B4DD",
    x"1E8B2B0",
    x"1E8B083",
    x"1E8AE57",
    x"1E8AC2C",
    x"1E8AA01",
    x"1E8A7D7",
    x"1E8A5AD",
    x"1E8A384",
    x"1E8A15C",
    x"1E89F33",
    x"1E89D0C",
    x"1E89AE5",
    x"1E898BE",
    x"1E89699",
    x"1E89473",
    x"1E8924E",
    x"1E8902A",
    x"1E88E06",
    x"1E88BE3",
    x"1E889C0",
    x"1E8879E",
    x"1E8857D",
    x"1E8835B",
    x"1E8813B",
    x"1E87F1B",
    x"1E87CFB",
    x"1E87ADC",
    x"1E878BE",
    x"1E876A0",
    x"1E87483",
    x"1E87266",
    x"1E87049",
    x"1E86E2E",
    x"1E86C12",
    x"1E869F7",
    x"1E867DD",
    x"1E865C4",
    x"1E863AA",
    x"1E86192",
    x"1E85F7A",
    x"1E85D62",
    x"1E85B4B",
    x"1E85934",
    x"1E8571E",
    x"1E85509",
    x"1E852F4",
    x"1E850DF",
    x"1E84ECB",
    x"1E84CB8",
    x"1E84AA5",
    x"1E84893",
    x"1E84681",
    x"1E8446F",
    x"1E8425E",
    x"1E8404E",
    x"1E83E3E",
    x"1E83C2F",
    x"1E83A20",
    x"1E83812",
    x"1E83604",
    x"1E833F7",
    x"1E831EA",
    x"1E82FDE",
    x"1E82DD2",
    x"1E82BC7",
    x"1E829BC",
    x"1E827B2",
    x"1E825A9",
    x"1E8239F",
    x"1E82197",
    x"1E81F8F",
    x"1E81D87",
    x"1E81B80",
    x"1E81979",
    x"1E81773",
    x"1E8156D",
    x"1E81368",
    x"1E81164",
    x"1E80F60",
    x"1E80D5C",
    x"1E80B59",
    x"1E80956",
    x"1E80754",
    x"1E80553",
    x"1E80352",
    x"1E80151",
    x"1E7FEA2",
    x"1E7FAA3",
    x"1E7F6A5",
    x"1E7F2A8",
    x"1E7EEAC",
    x"1E7EAB1",
    x"1E7E6B6",
    x"1E7E2BD",
    x"1E7DEC5",
    x"1E7DACE",
    x"1E7D6D8",
    x"1E7D2E2",
    x"1E7CEEE",
    x"1E7CAFB",
    x"1E7C709",
    x"1E7C317",
    x"1E7BF27",
    x"1E7BB38",
    x"1E7B74A",
    x"1E7B35C",
    x"1E7AF70",
    x"1E7AB85",
    x"1E7A79A",
    x"1E7A3B1",
    x"1E79FC8",
    x"1E79BE1",
    x"1E797FA",
    x"1E79415",
    x"1E79030",
    x"1E78C4D",
    x"1E7886A",
    x"1E78489",
    x"1E780A8",
    x"1E77CC8",
    x"1E778EA",
    x"1E7750C",
    x"1E7712F",
    x"1E76D53",
    x"1E76978",
    x"1E7659E",
    x"1E761C6",
    x"1E75DEE",
    x"1E75A17",
    x"1E75641",
    x"1E7526B",
    x"1E74E97",
    x"1E74AC4",
    x"1E746F2",
    x"1E74321",
    x"1E73F50",
    x"1E73B81",
    x"1E737B3",
    x"1E733E5",
    x"1E73019",
    x"1E72C4D",
    x"1E72882",
    x"1E724B9",
    x"1E720F0",
    x"1E71D28",
    x"1E71962",
    x"1E7159C",
    x"1E711D7",
    x"1E70E13",
    x"1E70A50",
    x"1E7068E",
    x"1E702CC",
    x"1E6FF0C",
    x"1E6FB4D",
    x"1E6F78F",
    x"1E6F3D1",
    x"1E6F015",
    x"1E6EC59",
    x"1E6E89E",
    x"1E6E4E5",
    x"1E6E12C",
    x"1E6DD74",
    x"1E6D9BD",
    x"1E6D607",
    x"1E6D252",
    x"1E6CE9E",
    x"1E6CAEB",
    x"1E6C739",
    x"1E6C387",
    x"1E6BFD7",
    x"1E6BC27",
    x"1E6B879",
    x"1E6B4CB",
    x"1E6B11E",
    x"1E6AD73",
    x"1E6A9C8",
    x"1E6A61E",
    x"1E6A275",
    x"1E69ECD",
    x"1E69B25",
    x"1E6977F",
    x"1E693DA",
    x"1E69035",
    x"1E68C91",
    x"1E688EF",
    x"1E6854D",
    x"1E681AC",
    x"1E67E0C",
    x"1E67A6D",
    x"1E676CF",
    x"1E67332",
    x"1E66F95",
    x"1E66BFA",
    x"1E6685F",
    x"1E664C6",
    x"1E6612D",
    x"1E65D95",
    x"1E659FE",
    x"1E65668",
    x"1E652D3",
    x"1E64F3F",
    x"1E64BAB",
    x"1E64819",
    x"1E64487",
    x"1E640F7",
    x"1E63D67",
    x"1E639D8",
    x"1E6364A",
    x"1E632BD",
    x"1E62F30",
    x"1E62BA5",
    x"1E6281B",
    x"1E62491",
    x"1E62108",
    x"1E61D81",
    x"1E619FA",
    x"1E61674",
    x"1E612EE",
    x"1E60F6A",
    x"1E60BE7",
    x"1E60864",
    x"1E604E2",
    x"1E60162",
    x"1E5FDE2",
    x"1E5FA63",
    x"1E5F6E5",
    x"1E5F367",
    x"1E5EFEB",
    x"1E5EC6F",
    x"1E5E8F5",
    x"1E5E57B",
    x"1E5E202",
    x"1E5DE8A",
    x"1E5DB13",
    x"1E5D79C",
    x"1E5D427",
    x"1E5D0B2",
    x"1E5CD3F",
    x"1E5C9CC",
    x"1E5C65A",
    x"1E5C2E8",
    x"1E5BF78",
    x"1E5BC09",
    x"1E5B89A",
    x"1E5B52C",
    x"1E5B1C0",
    x"1E5AE54",
    x"1E5AAE8",
    x"1E5A77E",
    x"1E5A415",
    x"1E5A0AC",
    x"1E59D44",
    x"1E599DD",
    x"1E59677",
    x"1E59312",
    x"1E58FAE",
    x"1E58C4A",
    x"1E588E8",
    x"1E58586",
    x"1E58225",
    x"1E57EC5",
    x"1E57B66",
    x"1E57807",
    x"1E574AA",
    x"1E5714D",
    x"1E56DF1",
    x"1E56A96",
    x"1E5673C",
    x"1E563E2",
    x"1E5608A",
    x"1E55D32",
    x"1E559DB",
    x"1E55685",
    x"1E55330",
    x"1E54FDB",
    x"1E54C88",
    x"1E54935",
    x"1E545E3",
    x"1E54292",
    x"1E53F42",
    x"1E53BF3",
    x"1E538A4",
    x"1E53556",
    x"1E53209",
    x"1E52EBD",
    x"1E52B72",
    x"1E52827",
    x"1E524DE",
    x"1E52195",
    x"1E51E4D",
    x"1E51B06",
    x"1E517C0",
    x"1E5147A",
    x"1E51135",
    x"1E50DF1",
    x"1E50AAE",
    x"1E5076C",
    x"1E5042B",
    x"1E500EA",
    x"1E4FDAA",
    x"1E4FA6B",
    x"1E4F72D",
    x"1E4F3F0",
    x"1E4F0B3",
    x"1E4ED77",
    x"1E4EA3C",
    x"1E4E702",
    x"1E4E3C9",
    x"1E4E090",
    x"1E4DD58",
    x"1E4DA22",
    x"1E4D6EB",
    x"1E4D3B6",
    x"1E4D082",
    x"1E4CD4E",
    x"1E4CA1B",
    x"1E4C6E9",
    x"1E4C3B7",
    x"1E4C087",
    x"1E4BD57",
    x"1E4BA28",
    x"1E4B6FA",
    x"1E4B3CD",
    x"1E4B0A0",
    x"1E4AD74",
    x"1E4AA49",
    x"1E4A71F",
    x"1E4A3F6",
    x"1E4A0CD",
    x"1E49DA5",
    x"1E49A7E",
    x"1E49758",
    x"1E49433",
    x"1E4910E",
    x"1E48DEA",
    x"1E48AC7",
    x"1E487A5",
    x"1E48483",
    x"1E48163",
    x"1E47E43",
    x"1E47B23",
    x"1E47805",
    x"1E474E7",
    x"1E471CB",
    x"1E46EAF",
    x"1E46B93",
    x"1E46879",
    x"1E4655F",
    x"1E46246",
    x"1E45F2E",
    x"1E45C17",
    x"1E45900",
    x"1E455EA",
    x"1E452D5",
    x"1E44FC1",
    x"1E44CAD",
    x"1E4499A",
    x"1E44688",
    x"1E44377",
    x"1E44067",
    x"1E43D57",
    x"1E43A48",
    x"1E4373A",
    x"1E4342C",
    x"1E43120",
    x"1E42E14",
    x"1E42B09",
    x"1E427FE",
    x"1E424F5",
    x"1E421EC",
    x"1E41EE4",
    x"1E41BDC",
    x"1E418D6",
    x"1E415D0",
    x"1E412CB",
    x"1E40FC6",
    x"1E40CC3",
    x"1E409C0",
    x"1E406BE",
    x"1E403BD",
    x"1E400BC",
    x"1E3FDBC",
    x"1E3FABD",
    x"1E3F7BF",
    x"1E3F4C1",
    x"1E3F1C5",
    x"1E3EEC8",
    x"1E3EBCD",
    x"1E3E8D3",
    x"1E3E5D9",
    x"1E3E2E0",
    x"1E3DFE7",
    x"1E3DCF0",
    x"1E3D9F9",
    x"1E3D703",
    x"1E3D40D",
    x"1E3D119",
    x"1E3CE25",
    x"1E3CB32",
    x"1E3C83F",
    x"1E3C54D",
    x"1E3C25D",
    x"1E3BF6C",
    x"1E3BC7D",
    x"1E3B98E",
    x"1E3B6A0",
    x"1E3B3B3",
    x"1E3B0C6",
    x"1E3ADDA",
    x"1E3AAEF",
    x"1E3A805",
    x"1E3A51B",
    x"1E3A232",
    x"1E39F4A",
    x"1E39C63",
    x"1E3997C",
    x"1E39696",
    x"1E393B1",
    x"1E390CC",
    x"1E38DE8",
    x"1E38B05",
    x"1E38823",
    x"1E38541",
    x"1E38260",
    x"1E37F80",
    x"1E37CA0",
    x"1E379C2",
    x"1E376E3",
    x"1E37406",
    x"1E37129",
    x"1E36E4E",
    x"1E36B72",
    x"1E36898",
    x"1E365BE",
    x"1E362E5",
    x"1E3600D",
    x"1E35D35",
    x"1E35A5E",
    x"1E35788",
    x"1E354B2",
    x"1E351DD",
    x"1E34F09",
    x"1E34C36",
    x"1E34963",
    x"1E34691",
    x"1E343C0",
    x"1E340EF",
    x"1E33E1F",
    x"1E33B50",
    x"1E33882",
    x"1E335B4",
    x"1E332E7",
    x"1E3301B",
    x"1E32D4F",
    x"1E32A84",
    x"1E327BA",
    x"1E324F0",
    x"1E32227",
    x"1E31F5F",
    x"1E31C97",
    x"1E319D1",
    x"1E3170B",
    x"1E31445",
    x"1E31180",
    x"1E30EBC",
    x"1E30BF9",
    x"1E30936",
    x"1E30674",
    x"1E303B3",
    x"1E300F3",
    x"1E2FE33",
    x"1E2FB73",
    x"1E2F8B5",
    x"1E2F5F7",
    x"1E2F33A",
    x"1E2F07D",
    x"1E2EDC2",
    x"1E2EB07",
    x"1E2E84C",
    x"1E2E592",
    x"1E2E2D9",
    x"1E2E021",
    x"1E2DD69",
    x"1E2DAB2",
    x"1E2D7FC",
    x"1E2D546",
    x"1E2D291",
    x"1E2CFDD",
    x"1E2CD29",
    x"1E2CA76",
    x"1E2C7C4",
    x"1E2C513",
    x"1E2C262",
    x"1E2BFB1",
    x"1E2BD02",
    x"1E2BA53",
    x"1E2B7A5",
    x"1E2B4F7",
    x"1E2B24A",
    x"1E2AF9E",
    x"1E2ACF2",
    x"1E2AA47",
    x"1E2A79D",
    x"1E2A4F4",
    x"1E2A24B",
    x"1E29FA2",
    x"1E29CFB",
    x"1E29A54",
    x"1E297AE",
    x"1E29508",
    x"1E29263",
    x"1E28FBF",
    x"1E28D1B",
    x"1E28A78",
    x"1E287D6",
    x"1E28534",
    x"1E28294",
    x"1E27FF3",
    x"1E27D54",
    x"1E27AB5",
    x"1E27816",
    x"1E27578",
    x"1E272DB",
    x"1E2703F",
    x"1E26DA3",
    x"1E26B08",
    x"1E2686E",
    x"1E265D4",
    x"1E2633B",
    x"1E260A2",
    x"1E25E0B",
    x"1E25B73",
    x"1E258DD",
    x"1E25647",
    x"1E253B2",
    x"1E2511D",
    x"1E24E89",
    x"1E24BF6",
    x"1E24963",
    x"1E246D1",
    x"1E24440",
    x"1E241AF",
    x"1E23F1F",
    x"1E23C8F",
    x"1E23A01",
    x"1E23772",
    x"1E234E5",
    x"1E23258",
    x"1E22FCC",
    x"1E22D40",
    x"1E22AB5",
    x"1E2282B",
    x"1E225A1",
    x"1E22318",
    x"1E2208F",
    x"1E21E08",
    x"1E21B80",
    x"1E218FA",
    x"1E21674",
    x"1E213EF",
    x"1E2116A",
    x"1E20EE6",
    x"1E20C63",
    x"1E209E0",
    x"1E2075E",
    x"1E204DC",
    x"1E2025B",
    x"1E1FFDB",
    x"1E1FD5B",
    x"1E1FADC",
    x"1E1F85E",
    x"1E1F5E0",
    x"1E1F363",
    x"1E1F0E6",
    x"1E1EE6A",
    x"1E1EBEF",
    x"1E1E974",
    x"1E1E6FA",
    x"1E1E481",
    x"1E1E208",
    x"1E1DF90",
    x"1E1DD18",
    x"1E1DAA1",
    x"1E1D82B",
    x"1E1D5B5",
    x"1E1D340",
    x"1E1D0CC",
    x"1E1CE58",
    x"1E1CBE5",
    x"1E1C972",
    x"1E1C700",
    x"1E1C48E",
    x"1E1C21E",
    x"1E1BFAD",
    x"1E1BD3E",
    x"1E1BACF",
    x"1E1B860",
    x"1E1B5F2",
    x"1E1B385",
    x"1E1B119",
    x"1E1AEAD",
    x"1E1AC41",
    x"1E1A9D7",
    x"1E1A76C",
    x"1E1A503",
    x"1E1A29A",
    x"1E1A032",
    x"1E19DCA",
    x"1E19B63",
    x"1E198FC",
    x"1E19696",
    x"1E19431",
    x"1E191CC",
    x"1E18F68",
    x"1E18D04",
    x"1E18AA1",
    x"1E1883F",
    x"1E185DD",
    x"1E1837C",
    x"1E1811C",
    x"1E17EBC",
    x"1E17C5C",
    x"1E179FD",
    x"1E1779F",
    x"1E17542",
    x"1E172E5",
    x"1E17088",
    x"1E16E2C",
    x"1E16BD1",
    x"1E16976",
    x"1E1671C",
    x"1E164C3",
    x"1E1626A",
    x"1E16012",
    x"1E15DBA",
    x"1E15B63",
    x"1E1590C",
    x"1E156B6",
    x"1E15461",
    x"1E1520C",
    x"1E14FB8",
    x"1E14D64",
    x"1E14B11",
    x"1E148BF",
    x"1E1466D",
    x"1E1441B",
    x"1E141CB",
    x"1E13F7B",
    x"1E13D2B",
    x"1E13ADC",
    x"1E1388E",
    x"1E13640",
    x"1E133F2",
    x"1E131A6",
    x"1E12F5A",
    x"1E12D0E",
    x"1E12AC3",
    x"1E12879",
    x"1E1262F",
    x"1E123E6",
    x"1E1219D",
    x"1E11F55",
    x"1E11D0D",
    x"1E11AC6",
    x"1E11880",
    x"1E1163A",
    x"1E113F5",
    x"1E111B0",
    x"1E10F6C",
    x"1E10D28",
    x"1E10AE5",
    x"1E108A3",
    x"1E10661",
    x"1E10420",
    x"1E101DF",
    x"1E0FF9F",
    x"1E0FD5F",
    x"1E0FB20",
    x"1E0F8E2",
    x"1E0F6A4",
    x"1E0F466",
    x"1E0F229",
    x"1E0EFED",
    x"1E0EDB1",
    x"1E0EB76",
    x"1E0E93C",
    x"1E0E702",
    x"1E0E4C8",
    x"1E0E28F",
    x"1E0E057",
    x"1E0DE1F",
    x"1E0DBE8",
    x"1E0D9B1",
    x"1E0D77B",
    x"1E0D545",
    x"1E0D310",
    x"1E0D0DC",
    x"1E0CEA8",
    x"1E0CC75",
    x"1E0CA42",
    x"1E0C80F",
    x"1E0C5DE",
    x"1E0C3AC",
    x"1E0C17C",
    x"1E0BF4C",
    x"1E0BD1C",
    x"1E0BAED",
    x"1E0B8BF",
    x"1E0B691",
    x"1E0B463",
    x"1E0B237",
    x"1E0B00A",
    x"1E0ADDF",
    x"1E0ABB3",
    x"1E0A989",
    x"1E0A75F",
    x"1E0A535",
    x"1E0A30C",
    x"1E0A0E4",
    x"1E09EBC",
    x"1E09C94",
    x"1E09A6D",
    x"1E09847",
    x"1E09621",
    x"1E093FC",
    x"1E091D7",
    x"1E08FB3",
    x"1E08D8F",
    x"1E08B6C",
    x"1E0894A",
    x"1E08728",
    x"1E08506",
    x"1E082E5",
    x"1E080C5",
    x"1E07EA5",
    x"1E07C85",
    x"1E07A66",
    x"1E07848",
    x"1E0762A",
    x"1E0740D",
    x"1E071F0",
    x"1E06FD4",
    x"1E06DB8",
    x"1E06B9D",
    x"1E06982",
    x"1E06768",
    x"1E0654F",
    x"1E06336",
    x"1E0611D",
    x"1E05F05",
    x"1E05CEE",
    x"1E05AD7",
    x"1E058C0",
    x"1E056AA",
    x"1E05495",
    x"1E05280",
    x"1E0506C",
    x"1E04E58",
    x"1E04C44",
    x"1E04A32",
    x"1E0481F",
    x"1E0460E",
    x"1E043FC",
    x"1E041EC",
    x"1E03FDB",
    x"1E03DCC",
    x"1E03BBD",
    x"1E039AE",
    x"1E037A0",
    x"1E03592",
    x"1E03385",
    x"1E03178",
    x"1E02F6C",
    x"1E02D61",
    x"1E02B55",
    x"1E0294B",
    x"1E02741",
    x"1E02537",
    x"1E0232E",
    x"1E02126",
    x"1E01F1E",
    x"1E01D16",
    x"1E01B0F",
    x"1E01909",
    x"1E01703",
    x"1E014FD",
    x"1E012F8",
    x"1E010F4",
    x"1E00EF0",
    x"1E00CEC",
    x"1E00AE9",
    x"1E008E7",
    x"1E006E5",
    x"1E004E3",
    x"1E002E2",
    x"1E000E2",
    x"1DFFDC4",
    x"1DFF9C5",
    x"1DFF5C7",
    x"1DFF1CA",
    x"1DFEDCE",
    x"1DFE9D3",
    x"1DFE5D9",
    x"1DFE1E0",
    x"1DFDDE8",
    x"1DFD9F1",
    x"1DFD5FB",
    x"1DFD206",
    x"1DFCE12",
    x"1DFCA1F",
    x"1DFC62D",
    x"1DFC23C",
    x"1DFBE4C",
    x"1DFBA5D",
    x"1DFB66F",
    x"1DFB282",
    x"1DFAE96",
    x"1DFAAAB",
    x"1DFA6C0",
    x"1DFA2D7",
    x"1DF9EEF",
    x"1DF9B08",
    x"1DF9722",
    x"1DF933C",
    x"1DF8F58",
    x"1DF8B75",
    x"1DF8792",
    x"1DF83B1",
    x"1DF7FD0",
    x"1DF7BF1",
    x"1DF7812",
    x"1DF7435",
    x"1DF7058",
    x"1DF6C7D",
    x"1DF68A2",
    x"1DF64C8",
    x"1DF60F0",
    x"1DF5D18",
    x"1DF5941",
    x"1DF556B",
    x"1DF5196",
    x"1DF4DC2",
    x"1DF49EF",
    x"1DF461D",
    x"1DF424C",
    x"1DF3E7C",
    x"1DF3AAD",
    x"1DF36DF",
    x"1DF3312",
    x"1DF2F45",
    x"1DF2B7A",
    x"1DF27B0",
    x"1DF23E6",
    x"1DF201E",
    x"1DF1C56",
    x"1DF1890",
    x"1DF14CA",
    x"1DF1105",
    x"1DF0D41",
    x"1DF097F",
    x"1DF05BD",
    x"1DF01FC",
    x"1DEFE3C",
    x"1DEFA7D",
    x"1DEF6BE",
    x"1DEF301",
    x"1DEEF45",
    x"1DEEB8A",
    x"1DEE7CF",
    x"1DEE416",
    x"1DEE05D",
    x"1DEDCA5",
    x"1DED8EF",
    x"1DED539",
    x"1DED184",
    x"1DECDD0",
    x"1DECA1D",
    x"1DEC66B",
    x"1DEC2BA",
    x"1DEBF0A",
    x"1DEBB5B",
    x"1DEB7AC",
    x"1DEB3FF",
    x"1DEB052",
    x"1DEACA7",
    x"1DEA8FC",
    x"1DEA552",
    x"1DEA1A9",
    x"1DE9E01",
    x"1DE9A5A",
    x"1DE96B4",
    x"1DE930F",
    x"1DE8F6B",
    x"1DE8BC7",
    x"1DE8825",
    x"1DE8483",
    x"1DE80E2",
    x"1DE7D43",
    x"1DE79A4",
    x"1DE7606",
    x"1DE7269",
    x"1DE6ECD",
    x"1DE6B31",
    x"1DE6797",
    x"1DE63FE",
    x"1DE6065",
    x"1DE5CCD",
    x"1DE5937",
    x"1DE55A1",
    x"1DE520C",
    x"1DE4E78",
    x"1DE4AE5",
    x"1DE4752",
    x"1DE43C1",
    x"1DE4030",
    x"1DE3CA1",
    x"1DE3912",
    x"1DE3584",
    x"1DE31F7",
    x"1DE2E6B",
    x"1DE2AE0",
    x"1DE2756",
    x"1DE23CC",
    x"1DE2044",
    x"1DE1CBC",
    x"1DE1936",
    x"1DE15B0",
    x"1DE122B",
    x"1DE0EA7",
    x"1DE0B23",
    x"1DE07A1",
    x"1DE0420",
    x"1DE009F",
    x"1DDFD1F",
    x"1DDF9A0",
    x"1DDF622",
    x"1DDF2A5",
    x"1DDEF29",
    x"1DDEBAE",
    x"1DDE833",
    x"1DDE4BA",
    x"1DDE141",
    x"1DDDDC9",
    x"1DDDA52",
    x"1DDD6DC",
    x"1DDD367",
    x"1DDCFF2",
    x"1DDCC7F",
    x"1DDC90C",
    x"1DDC59A",
    x"1DDC229",
    x"1DDBEB9",
    x"1DDBB4A",
    x"1DDB7DB",
    x"1DDB46E",
    x"1DDB101",
    x"1DDAD95",
    x"1DDAA2A",
    x"1DDA6C0",
    x"1DDA357",
    x"1DD9FEF",
    x"1DD9C87",
    x"1DD9920",
    x"1DD95BA",
    x"1DD9255",
    x"1DD8EF1",
    x"1DD8B8E",
    x"1DD882B",
    x"1DD84CA",
    x"1DD8169",
    x"1DD7E09",
    x"1DD7AAA",
    x"1DD774C",
    x"1DD73EE",
    x"1DD7092",
    x"1DD6D36",
    x"1DD69DB",
    x"1DD6681",
    x"1DD6328",
    x"1DD5FD0",
    x"1DD5C78",
    x"1DD5921",
    x"1DD55CC",
    x"1DD5276",
    x"1DD4F22",
    x"1DD4BCF",
    x"1DD487C",
    x"1DD452B",
    x"1DD41DA",
    x"1DD3E8A",
    x"1DD3B3B",
    x"1DD37EC",
    x"1DD349F",
    x"1DD3152",
    x"1DD2E06",
    x"1DD2ABB",
    x"1DD2771",
    x"1DD2427",
    x"1DD20DE",
    x"1DD1D97",
    x"1DD1A50",
    x"1DD1709",
    x"1DD13C4",
    x"1DD1080",
    x"1DD0D3C",
    x"1DD09F9",
    x"1DD06B7",
    x"1DD0376",
    x"1DD0035",
    x"1DCFCF6",
    x"1DCF9B7",
    x"1DCF679",
    x"1DCF33B",
    x"1DCEFFF",
    x"1DCECC3",
    x"1DCE989",
    x"1DCE64F",
    x"1DCE316",
    x"1DCDFDD",
    x"1DCDCA6",
    x"1DCD96F",
    x"1DCD639",
    x"1DCD304",
    x"1DCCFCF",
    x"1DCCC9C",
    x"1DCC969",
    x"1DCC637",
    x"1DCC306",
    x"1DCBFD6",
    x"1DCBCA6",
    x"1DCB977",
    x"1DCB649",
    x"1DCB31C",
    x"1DCAFF0",
    x"1DCACC4",
    x"1DCA999",
    x"1DCA66F",
    x"1DCA346",
    x"1DCA01E",
    x"1DC9CF6",
    x"1DC99CF",
    x"1DC96A9",
    x"1DC9384",
    x"1DC905F",
    x"1DC8D3C",
    x"1DC8A19",
    x"1DC86F7",
    x"1DC83D5",
    x"1DC80B5",
    x"1DC7D95",
    x"1DC7A76",
    x"1DC7758",
    x"1DC743A",
    x"1DC711E",
    x"1DC6E02",
    x"1DC6AE7",
    x"1DC67CC",
    x"1DC64B3",
    x"1DC619A",
    x"1DC5E82",
    x"1DC5B6B",
    x"1DC5854",
    x"1DC553E",
    x"1DC522A",
    x"1DC4F15",
    x"1DC4C02",
    x"1DC48EF",
    x"1DC45DE",
    x"1DC42CC",
    x"1DC3FBC",
    x"1DC3CAD",
    x"1DC399E",
    x"1DC3690",
    x"1DC3383",
    x"1DC3076",
    x"1DC2D6A",
    x"1DC2A5F",
    x"1DC2755",
    x"1DC244C",
    x"1DC2143",
    x"1DC1E3B",
    x"1DC1B34",
    x"1DC182D",
    x"1DC1528",
    x"1DC1223",
    x"1DC0F1F",
    x"1DC0C1B",
    x"1DC0919",
    x"1DC0617",
    x"1DC0316",
    x"1DC0015",
    x"1DBFD16",
    x"1DBFA17",
    x"1DBF719",
    x"1DBF41B",
    x"1DBF11E",
    x"1DBEE23",
    x"1DBEB27",
    x"1DBE82D",
    x"1DBE533",
    x"1DBE23A",
    x"1DBDF42",
    x"1DBDC4B",
    x"1DBD954",
    x"1DBD65E",
    x"1DBD369",
    x"1DBD074",
    x"1DBCD81",
    x"1DBCA8E",
    x"1DBC79B",
    x"1DBC4AA",
    x"1DBC1B9",
    x"1DBBEC9",
    x"1DBBBDA",
    x"1DBB8EB",
    x"1DBB5FD",
    x"1DBB310",
    x"1DBB024",
    x"1DBAD38",
    x"1DBAA4D",
    x"1DBA763",
    x"1DBA479",
    x"1DBA191",
    x"1DB9EA9",
    x"1DB9BC1",
    x"1DB98DB",
    x"1DB95F5",
    x"1DB9310",
    x"1DB902B",
    x"1DB8D48",
    x"1DB8A65",
    x"1DB8782",
    x"1DB84A1",
    x"1DB81C0",
    x"1DB7EE0",
    x"1DB7C01",
    x"1DB7922",
    x"1DB7644",
    x"1DB7367",
    x"1DB708A",
    x"1DB6DAF",
    x"1DB6AD4",
    x"1DB67F9",
    x"1DB6520",
    x"1DB6247",
    x"1DB5F6E",
    x"1DB5C97",
    x"1DB59C0",
    x"1DB56EA",
    x"1DB5415",
    x"1DB5140",
    x"1DB4E6C",
    x"1DB4B99",
    x"1DB48C6",
    x"1DB45F4",
    x"1DB4323",
    x"1DB4053",
    x"1DB3D83",
    x"1DB3AB4",
    x"1DB37E6",
    x"1DB3518",
    x"1DB324B",
    x"1DB2F7F",
    x"1DB2CB3",
    x"1DB29E9",
    x"1DB271E",
    x"1DB2455",
    x"1DB218C",
    x"1DB1EC4",
    x"1DB1BFD",
    x"1DB1936",
    x"1DB1670",
    x"1DB13AB",
    x"1DB10E6",
    x"1DB0E23",
    x"1DB0B5F",
    x"1DB089D",
    x"1DB05DB",
    x"1DB031A",
    x"1DB005A",
    x"1DAFD9A",
    x"1DAFADB",
    x"1DAF81C",
    x"1DAF55F",
    x"1DAF2A2",
    x"1DAEFE5",
    x"1DAED2A",
    x"1DAEA6F",
    x"1DAE7B5",
    x"1DAE4FB",
    x"1DAE242",
    x"1DADF8A",
    x"1DADCD2",
    x"1DADA1B",
    x"1DAD765",
    x"1DAD4B0",
    x"1DAD1FB",
    x"1DACF47",
    x"1DACC93",
    x"1DAC9E0",
    x"1DAC72E",
    x"1DAC47D",
    x"1DAC1CC",
    x"1DABF1C",
    x"1DABC6C",
    x"1DAB9BE",
    x"1DAB710",
    x"1DAB462",
    x"1DAB1B5",
    x"1DAAF09",
    x"1DAAC5E",
    x"1DAA9B3",
    x"1DAA709",
    x"1DAA460",
    x"1DAA1B7",
    x"1DA9F0F",
    x"1DA9C67",
    x"1DA99C1",
    x"1DA971A",
    x"1DA9475",
    x"1DA91D0",
    x"1DA8F2C",
    x"1DA8C89",
    x"1DA89E6",
    x"1DA8744",
    x"1DA84A2",
    x"1DA8201",
    x"1DA7F61",
    x"1DA7CC2",
    x"1DA7A23",
    x"1DA7785",
    x"1DA74E7",
    x"1DA724A",
    x"1DA6FAE",
    x"1DA6D12",
    x"1DA6A77",
    x"1DA67DD",
    x"1DA6543",
    x"1DA62AA",
    x"1DA6012",
    x"1DA5D7A",
    x"1DA5AE3",
    x"1DA584D",
    x"1DA55B7",
    x"1DA5322",
    x"1DA508E",
    x"1DA4DFA",
    x"1DA4B67",
    x"1DA48D4",
    x"1DA4642",
    x"1DA43B1",
    x"1DA4120",
    x"1DA3E90",
    x"1DA3C01",
    x"1DA3972",
    x"1DA36E4",
    x"1DA3457",
    x"1DA31CA",
    x"1DA2F3E",
    x"1DA2CB3",
    x"1DA2A28",
    x"1DA279E",
    x"1DA2514",
    x"1DA228B",
    x"1DA2003",
    x"1DA1D7B",
    x"1DA1AF4",
    x"1DA186D",
    x"1DA15E8",
    x"1DA1363",
    x"1DA10DE",
    x"1DA0E5A",
    x"1DA0BD7",
    x"1DA0954",
    x"1DA06D2",
    x"1DA0451",
    x"1DA01D0",
    x"1D9FF50",
    x"1D9FCD0",
    x"1D9FA51",
    x"1D9F7D3",
    x"1D9F556",
    x"1D9F2D9",
    x"1D9F05C",
    x"1D9EDE0",
    x"1D9EB65",
    x"1D9E8EB",
    x"1D9E671",
    x"1D9E3F7",
    x"1D9E17F",
    x"1D9DF07",
    x"1D9DC8F",
    x"1D9DA18",
    x"1D9D7A2",
    x"1D9D52D",
    x"1D9D2B8",
    x"1D9D043",
    x"1D9CDCF",
    x"1D9CB5C",
    x"1D9C8EA",
    x"1D9C678",
    x"1D9C407",
    x"1D9C196",
    x"1D9BF26",
    x"1D9BCB6",
    x"1D9BA47",
    x"1D9B7D9",
    x"1D9B56B",
    x"1D9B2FE",
    x"1D9B092",
    x"1D9AE26",
    x"1D9ABBB",
    x"1D9A950",
    x"1D9A6E6",
    x"1D9A47D",
    x"1D9A214",
    x"1D99FAC",
    x"1D99D44",
    x"1D99ADD",
    x"1D99877",
    x"1D99611",
    x"1D993AC",
    x"1D99147",
    x"1D98EE3",
    x"1D98C80",
    x"1D98A1D",
    x"1D987BB",
    x"1D98559",
    x"1D982F8",
    x"1D98097",
    x"1D97E38",
    x"1D97BD8",
    x"1D9797A",
    x"1D9771C",
    x"1D974BE",
    x"1D97261",
    x"1D97005",
    x"1D96DA9",
    x"1D96B4E",
    x"1D968F4",
    x"1D9669A",
    x"1D96440",
    x"1D961E7",
    x"1D95F8F",
    x"1D95D38",
    x"1D95AE1",
    x"1D9588A",
    x"1D95634",
    x"1D953DF",
    x"1D9518A",
    x"1D94F36",
    x"1D94CE3",
    x"1D94A90",
    x"1D9483E",
    x"1D945EC",
    x"1D9439B",
    x"1D9414A",
    x"1D93EFA",
    x"1D93CAB",
    x"1D93A5C",
    x"1D9380D",
    x"1D935C0",
    x"1D93372",
    x"1D93126",
    x"1D92EDA",
    x"1D92C8E",
    x"1D92A44",
    x"1D927F9",
    x"1D925B0",
    x"1D92366",
    x"1D9211E",
    x"1D91ED6",
    x"1D91C8F",
    x"1D91A48",
    x"1D91801",
    x"1D915BC",
    x"1D91376",
    x"1D91132",
    x"1D90EEE",
    x"1D90CAA",
    x"1D90A68",
    x"1D90825",
    x"1D905E3",
    x"1D903A2",
    x"1D90162",
    x"1D8FF22",
    x"1D8FCE2",
    x"1D8FAA3",
    x"1D8F865",
    x"1D8F627",
    x"1D8F3EA",
    x"1D8F1AD",
    x"1D8EF71",
    x"1D8ED35",
    x"1D8EAFA",
    x"1D8E8C0",
    x"1D8E686",
    x"1D8E44D",
    x"1D8E214",
    x"1D8DFDB",
    x"1D8DDA4",
    x"1D8DB6D",
    x"1D8D936",
    x"1D8D700",
    x"1D8D4CB",
    x"1D8D296",
    x"1D8D061",
    x"1D8CE2D",
    x"1D8CBFA",
    x"1D8C9C7",
    x"1D8C795",
    x"1D8C564",
    x"1D8C333",
    x"1D8C102",
    x"1D8BED2",
    x"1D8BCA3",
    x"1D8BA74",
    x"1D8B845",
    x"1D8B618",
    x"1D8B3EA",
    x"1D8B1BE",
    x"1D8AF92",
    x"1D8AD66",
    x"1D8AB3B",
    x"1D8A910",
    x"1D8A6E6",
    x"1D8A4BD",
    x"1D8A294",
    x"1D8A06C",
    x"1D89E44",
    x"1D89C1C",
    x"1D899F6",
    x"1D897CF",
    x"1D895AA",
    x"1D89385",
    x"1D89160",
    x"1D88F3C",
    x"1D88D18",
    x"1D88AF5",
    x"1D888D3",
    x"1D886B1",
    x"1D88490",
    x"1D8826F",
    x"1D8804E",
    x"1D87E2F",
    x"1D87C0F",
    x"1D879F1",
    x"1D877D2",
    x"1D875B5",
    x"1D87397",
    x"1D8717B",
    x"1D86F5F",
    x"1D86D43",
    x"1D86B28",
    x"1D8690E",
    x"1D866F4",
    x"1D864DA",
    x"1D862C1",
    x"1D860A9",
    x"1D85E91",
    x"1D85C79",
    x"1D85A63",
    x"1D8584C",
    x"1D85636",
    x"1D85421",
    x"1D8520C",
    x"1D84FF8",
    x"1D84DE4",
    x"1D84BD1",
    x"1D849BE",
    x"1D847AC",
    x"1D8459B",
    x"1D84389",
    x"1D84179",
    x"1D83F69",
    x"1D83D59",
    x"1D83B4A",
    x"1D8393B",
    x"1D8372D",
    x"1D83520",
    x"1D83313",
    x"1D83106",
    x"1D82EFA",
    x"1D82CEF",
    x"1D82AE4",
    x"1D828D9",
    x"1D826CF",
    x"1D824C6",
    x"1D822BD",
    x"1D820B5",
    x"1D81EAD",
    x"1D81CA5",
    x"1D81A9E",
    x"1D81898",
    x"1D81692",
    x"1D8148D",
    x"1D81288",
    x"1D81083",
    x"1D80E80",
    x"1D80C7C",
    x"1D80A79",
    x"1D80877",
    x"1D80675",
    x"1D80474",
    x"1D80273",
    x"1D80072",
    x"1D7FCE6",
    x"1D7F8E7",
    x"1D7F4E9",
    x"1D7F0ED",
    x"1D7ECF1",
    x"1D7E8F6",
    x"1D7E4FC",
    x"1D7E104",
    x"1D7DD0C",
    x"1D7D915",
    x"1D7D51F",
    x"1D7D12A",
    x"1D7CD37",
    x"1D7C944",
    x"1D7C552",
    x"1D7C161",
    x"1D7BD71",
    x"1D7B982",
    x"1D7B595",
    x"1D7B1A8",
    x"1D7ADBC",
    x"1D7A9D1",
    x"1D7A5E7",
    x"1D7A1FE",
    x"1D79E16",
    x"1D79A2F",
    x"1D79649",
    x"1D79264",
    x"1D78E80",
    x"1D78A9C",
    x"1D786BA",
    x"1D782D9",
    x"1D77EF9",
    x"1D77B1A",
    x"1D7773B",
    x"1D7735E",
    x"1D76F82",
    x"1D76BA6",
    x"1D767CC",
    x"1D763F2",
    x"1D7601A",
    x"1D75C42",
    x"1D7586C",
    x"1D75496",
    x"1D750C1",
    x"1D74CEE",
    x"1D7491B",
    x"1D74549",
    x"1D74178",
    x"1D73DA8",
    x"1D739D9",
    x"1D7360B",
    x"1D7323E",
    x"1D72E72",
    x"1D72AA7",
    x"1D726DD",
    x"1D72314",
    x"1D71F4B",
    x"1D71B84",
    x"1D717BE",
    x"1D713F8",
    x"1D71034",
    x"1D70C70",
    x"1D708AD",
    x"1D704EC",
    x"1D7012B",
    x"1D6FD6B",
    x"1D6F9AC",
    x"1D6F5EE",
    x"1D6F231",
    x"1D6EE75",
    x"1D6EABA",
    x"1D6E700",
    x"1D6E347",
    x"1D6DF8E",
    x"1D6DBD7",
    x"1D6D820",
    x"1D6D46B",
    x"1D6D0B6",
    x"1D6CD02",
    x"1D6C950",
    x"1D6C59E",
    x"1D6C1ED",
    x"1D6BE3D",
    x"1D6BA8E",
    x"1D6B6E0",
    x"1D6B332",
    x"1D6AF86",
    x"1D6ABDA",
    x"1D6A830",
    x"1D6A486",
    x"1D6A0DE",
    x"1D69D36",
    x"1D6998F",
    x"1D695E9",
    x"1D69244",
    x"1D68EA0",
    x"1D68AFD",
    x"1D6875B",
    x"1D683B9",
    x"1D68019",
    x"1D67C79",
    x"1D678DA",
    x"1D6753D",
    x"1D671A0",
    x"1D66E04",
    x"1D66A69",
    x"1D666CF",
    x"1D66335",
    x"1D65F9D",
    x"1D65C06",
    x"1D6586F",
    x"1D654D9",
    x"1D65145",
    x"1D64DB1",
    x"1D64A1E",
    x"1D6468C",
    x"1D642FB",
    x"1D63F6A",
    x"1D63BDB",
    x"1D6384C",
    x"1D634BF",
    x"1D63132",
    x"1D62DA6",
    x"1D62A1B",
    x"1D62691",
    x"1D62308",
    x"1D61F7F",
    x"1D61BF8",
    x"1D61871",
    x"1D614EC",
    x"1D61167",
    x"1D60DE3",
    x"1D60A60",
    x"1D606DE",
    x"1D6035D",
    x"1D5FFDC",
    x"1D5FC5D",
    x"1D5F8DE",
    x"1D5F560",
    x"1D5F1E3",
    x"1D5EE67",
    x"1D5EAEC",
    x"1D5E772",
    x"1D5E3F8",
    x"1D5E080",
    x"1D5DD08",
    x"1D5D991",
    x"1D5D61B",
    x"1D5D2A6",
    x"1D5CF32",
    x"1D5CBBF",
    x"1D5C84C",
    x"1D5C4DB",
    x"1D5C16A",
    x"1D5BDFA",
    x"1D5BA8B",
    x"1D5B71D",
    x"1D5B3AF",
    x"1D5B043",
    x"1D5ACD7",
    x"1D5A96C",
    x"1D5A602",
    x"1D5A299",
    x"1D59F31",
    x"1D59BCA",
    x"1D59863",
    x"1D594FE",
    x"1D59199",
    x"1D58E35",
    x"1D58AD2",
    x"1D5876F",
    x"1D5840E",
    x"1D580AD",
    x"1D57D4E",
    x"1D579EF",
    x"1D57691",
    x"1D57333",
    x"1D56FD7",
    x"1D56C7B",
    x"1D56921",
    x"1D565C7",
    x"1D5626E",
    x"1D55F16",
    x"1D55BBE",
    x"1D55868",
    x"1D55512",
    x"1D551BD",
    x"1D54E69",
    x"1D54B16",
    x"1D547C4",
    x"1D54472",
    x"1D54121",
    x"1D53DD2",
    x"1D53A83",
    x"1D53734",
    x"1D533E7",
    x"1D5309A",
    x"1D52D4F",
    x"1D52A04",
    x"1D526BA",
    x"1D52370",
    x"1D52028",
    x"1D51CE0",
    x"1D51999",
    x"1D51653",
    x"1D5130E",
    x"1D50FCA",
    x"1D50C86",
    x"1D50944",
    x"1D50602",
    x"1D502C1",
    x"1D4FF80",
    x"1D4FC41",
    x"1D4F902",
    x"1D4F5C4",
    x"1D4F287",
    x"1D4EF4B",
    x"1D4EC10",
    x"1D4E8D5",
    x"1D4E59B",
    x"1D4E262",
    x"1D4DF2A",
    x"1D4DBF3",
    x"1D4D8BC",
    x"1D4D586",
    x"1D4D251",
    x"1D4CF1D",
    x"1D4CBEA",
    x"1D4C8B7",
    x"1D4C585",
    x"1D4C254",
    x"1D4BF24",
    x"1D4BBF5",
    x"1D4B8C6",
    x"1D4B599",
    x"1D4B26C",
    x"1D4AF3F",
    x"1D4AC14",
    x"1D4A8E9",
    x"1D4A5BF",
    x"1D4A296",
    x"1D49F6E",
    x"1D49C47",
    x"1D49920",
    x"1D495FA",
    x"1D492D5",
    x"1D48FB1",
    x"1D48C8D",
    x"1D4896A",
    x"1D48648",
    x"1D48327",
    x"1D48007",
    x"1D47CE7",
    x"1D479C8",
    x"1D476AA",
    x"1D4738D",
    x"1D47071",
    x"1D46D55",
    x"1D46A3A",
    x"1D46720",
    x"1D46406",
    x"1D460EE",
    x"1D45DD6",
    x"1D45ABF",
    x"1D457A9",
    x"1D45493",
    x"1D4517E",
    x"1D44E6A",
    x"1D44B57",
    x"1D44845",
    x"1D44533",
    x"1D44222",
    x"1D43F12",
    x"1D43C02",
    x"1D438F4",
    x"1D435E6",
    x"1D432D9",
    x"1D42FCD",
    x"1D42CC1",
    x"1D429B6",
    x"1D426AC",
    x"1D423A3",
    x"1D4209A",
    x"1D41D93",
    x"1D41A8C",
    x"1D41785",
    x"1D41480",
    x"1D4117B",
    x"1D40E77",
    x"1D40B74",
    x"1D40871",
    x"1D40570",
    x"1D4026F",
    x"1D3FF6E",
    x"1D3FC6F",
    x"1D3F970",
    x"1D3F672",
    x"1D3F375",
    x"1D3F078",
    x"1D3ED7D",
    x"1D3EA82",
    x"1D3E787",
    x"1D3E48E",
    x"1D3E195",
    x"1D3DE9D",
    x"1D3DBA6",
    x"1D3D8AF",
    x"1D3D5B9",
    x"1D3D2C4",
    x"1D3CFD0",
    x"1D3CCDC",
    x"1D3C9EA",
    x"1D3C6F8",
    x"1D3C406",
    x"1D3C116",
    x"1D3BE26",
    x"1D3BB36",
    x"1D3B848",
    x"1D3B55A",
    x"1D3B26D",
    x"1D3AF81",
    x"1D3AC96",
    x"1D3A9AB",
    x"1D3A6C1",
    x"1D3A3D7",
    x"1D3A0EF",
    x"1D39E07",
    x"1D39B20",
    x"1D39839",
    x"1D39554",
    x"1D3926F",
    x"1D38F8A",
    x"1D38CA7",
    x"1D389C4",
    x"1D386E2",
    x"1D38401",
    x"1D38120",
    x"1D37E40",
    x"1D37B61",
    x"1D37882",
    x"1D375A5",
    x"1D372C8",
    x"1D36FEB",
    x"1D36D10",
    x"1D36A35",
    x"1D3675B",
    x"1D36481",
    x"1D361A8",
    x"1D35ED0",
    x"1D35BF9",
    x"1D35922",
    x"1D3564C",
    x"1D35377",
    x"1D350A3",
    x"1D34DCF",
    x"1D34AFC",
    x"1D34829",
    x"1D34558",
    x"1D34287",
    x"1D33FB6",
    x"1D33CE7",
    x"1D33A18",
    x"1D3374A",
    x"1D3347C",
    x"1D331AF",
    x"1D32EE3",
    x"1D32C18",
    x"1D3294D",
    x"1D32683",
    x"1D323BA",
    x"1D320F2",
    x"1D31E2A",
    x"1D31B62",
    x"1D3189C",
    x"1D315D6",
    x"1D31311",
    x"1D3104D",
    x"1D30D89",
    x"1D30AC6",
    x"1D30803",
    x"1D30542",
    x"1D30281",
    x"1D2FFC1",
    x"1D2FD01",
    x"1D2FA42",
    x"1D2F784",
    x"1D2F4C6",
    x"1D2F209",
    x"1D2EF4D",
    x"1D2EC92",
    x"1D2E9D7",
    x"1D2E71D",
    x"1D2E463",
    x"1D2E1AB",
    x"1D2DEF3",
    x"1D2DC3B",
    x"1D2D984",
    x"1D2D6CE",
    x"1D2D419",
    x"1D2D164",
    x"1D2CEB0",
    x"1D2CBFD",
    x"1D2C94A",
    x"1D2C698",
    x"1D2C3E7",
    x"1D2C136",
    x"1D2BE86",
    x"1D2BBD7",
    x"1D2B929",
    x"1D2B67B",
    x"1D2B3CD",
    x"1D2B121",
    x"1D2AE75",
    x"1D2ABC9",
    x"1D2A91F",
    x"1D2A675",
    x"1D2A3CC",
    x"1D2A123",
    x"1D29E7B",
    x"1D29BD4",
    x"1D2992D",
    x"1D29687",
    x"1D293E2",
    x"1D2913D",
    x"1D28E99",
    x"1D28BF6",
    x"1D28953",
    x"1D286B1",
    x"1D28410",
    x"1D2816F",
    x"1D27ECF",
    x"1D27C30",
    x"1D27991",
    x"1D276F3",
    x"1D27456",
    x"1D271B9",
    x"1D26F1D",
    x"1D26C81",
    x"1D269E7",
    x"1D2674C",
    x"1D264B3",
    x"1D2621A",
    x"1D25F82",
    x"1D25CEA",
    x"1D25A53",
    x"1D257BD",
    x"1D25528",
    x"1D25293",
    x"1D24FFE",
    x"1D24D6B",
    x"1D24AD8",
    x"1D24845",
    x"1D245B3",
    x"1D24322",
    x"1D24092",
    x"1D23E02",
    x"1D23B73",
    x"1D238E4",
    x"1D23656",
    x"1D233C9",
    x"1D2313C",
    x"1D22EB0",
    x"1D22C25",
    x"1D2299A",
    x"1D22710",
    x"1D22487",
    x"1D221FE",
    x"1D21F76",
    x"1D21CEE",
    x"1D21A67",
    x"1D217E1",
    x"1D2155B",
    x"1D212D6",
    x"1D21052",
    x"1D20DCE",
    x"1D20B4B",
    x"1D208C9",
    x"1D20647",
    x"1D203C5",
    x"1D20145",
    x"1D1FEC5",
    x"1D1FC45",
    x"1D1F9C7",
    x"1D1F749",
    x"1D1F4CB",
    x"1D1F24E",
    x"1D1EFD2",
    x"1D1ED56",
    x"1D1EADB",
    x"1D1E861",
    x"1D1E5E7",
    x"1D1E36E",
    x"1D1E0F5",
    x"1D1DE7D",
    x"1D1DC06",
    x"1D1D98F",
    x"1D1D719",
    x"1D1D4A4",
    x"1D1D22F",
    x"1D1CFBB",
    x"1D1CD47",
    x"1D1CAD4",
    x"1D1C862",
    x"1D1C5F0",
    x"1D1C37F",
    x"1D1C10E",
    x"1D1BE9E",
    x"1D1BC2F",
    x"1D1B9C0",
    x"1D1B752",
    x"1D1B4E4",
    x"1D1B278",
    x"1D1B00B",
    x"1D1ADA0",
    x"1D1AB34",
    x"1D1A8CA",
    x"1D1A660",
    x"1D1A3F7",
    x"1D1A18E",
    x"1D19F26",
    x"1D19CBE",
    x"1D19A58",
    x"1D197F1",
    x"1D1958C",
    x"1D19327",
    x"1D190C2",
    x"1D18E5E",
    x"1D18BFB",
    x"1D18998",
    x"1D18736",
    x"1D184D5",
    x"1D18274",
    x"1D18013",
    x"1D17DB4",
    x"1D17B54",
    x"1D178F6",
    x"1D17698",
    x"1D1743B",
    x"1D171DE",
    x"1D16F82",
    x"1D16D26",
    x"1D16ACB",
    x"1D16871",
    x"1D16617",
    x"1D163BE",
    x"1D16165",
    x"1D15F0D",
    x"1D15CB5",
    x"1D15A5F",
    x"1D15808",
    x"1D155B3",
    x"1D1535D",
    x"1D15109",
    x"1D14EB5",
    x"1D14C62",
    x"1D14A0F",
    x"1D147BD",
    x"1D1456B",
    x"1D1431A",
    x"1D140C9",
    x"1D13E79",
    x"1D13C2A",
    x"1D139DB",
    x"1D1378D",
    x"1D13540",
    x"1D132F3",
    x"1D130A6",
    x"1D12E5A",
    x"1D12C0F",
    x"1D129C4",
    x"1D1277A",
    x"1D12530",
    x"1D122E7",
    x"1D1209F",
    x"1D11E57",
    x"1D11C10",
    x"1D119C9",
    x"1D11783",
    x"1D1153D",
    x"1D112F8",
    x"1D110B4",
    x"1D10E70",
    x"1D10C2D",
    x"1D109EA",
    x"1D107A8",
    x"1D10566",
    x"1D10325",
    x"1D100E4",
    x"1D0FEA5",
    x"1D0FC65",
    x"1D0FA26",
    x"1D0F7E8",
    x"1D0F5AA",
    x"1D0F36D",
    x"1D0F131",
    x"1D0EEF5",
    x"1D0ECB9",
    x"1D0EA7E",
    x"1D0E844",
    x"1D0E60A",
    x"1D0E3D1",
    x"1D0E198",
    x"1D0DF60",
    x"1D0DD29",
    x"1D0DAF2",
    x"1D0D8BB",
    x"1D0D685",
    x"1D0D450",
    x"1D0D21B",
    x"1D0CFE7",
    x"1D0CDB3",
    x"1D0CB80",
    x"1D0C94D",
    x"1D0C71B",
    x"1D0C4EA",
    x"1D0C2B9",
    x"1D0C088",
    x"1D0BE59",
    x"1D0BC29",
    x"1D0B9FA",
    x"1D0B7CC",
    x"1D0B59F",
    x"1D0B371",
    x"1D0B145",
    x"1D0AF19",
    x"1D0ACED",
    x"1D0AAC2",
    x"1D0A898",
    x"1D0A66E",
    x"1D0A445",
    x"1D0A21C",
    x"1D09FF4",
    x"1D09DCC",
    x"1D09BA5",
    x"1D0997E",
    x"1D09758",
    x"1D09532",
    x"1D0930D",
    x"1D090E9",
    x"1D08EC5",
    x"1D08CA1",
    x"1D08A7F",
    x"1D0885C",
    x"1D0863A",
    x"1D08419",
    x"1D081F8",
    x"1D07FD8",
    x"1D07DB8",
    x"1D07B99",
    x"1D0797B",
    x"1D0775D",
    x"1D0753F",
    x"1D07322",
    x"1D07105",
    x"1D06EE9",
    x"1D06CCE",
    x"1D06AB3",
    x"1D06899",
    x"1D0667F",
    x"1D06465",
    x"1D0624C",
    x"1D06034",
    x"1D05E1C",
    x"1D05C05",
    x"1D059EE",
    x"1D057D8",
    x"1D055C2",
    x"1D053AD",
    x"1D05199",
    x"1D04F84",
    x"1D04D71",
    x"1D04B5E",
    x"1D0494B",
    x"1D04739",
    x"1D04528",
    x"1D04317",
    x"1D04106",
    x"1D03EF6",
    x"1D03CE7",
    x"1D03AD8",
    x"1D038C9",
    x"1D036BB",
    x"1D034AE",
    x"1D032A1",
    x"1D03094",
    x"1D02E89",
    x"1D02C7D",
    x"1D02A72",
    x"1D02868",
    x"1D0265E",
    x"1D02455",
    x"1D0224C",
    x"1D02044",
    x"1D01E3C",
    x"1D01C34",
    x"1D01A2E",
    x"1D01827",
    x"1D01622",
    x"1D0141C",
    x"1D01218",
    x"1D01013",
    x"1D00E10",
    x"1D00C0C",
    x"1D00A09",
    x"1D00807",
    x"1D00605",
    x"1D00404",
    x"1D00203",
    x"1D00003",
    x"1CFFC07",
    x"1CFF809",
    x"1CFF40B",
    x"1CFF00F",
    x"1CFEC13",
    x"1CFE819",
    x"1CFE41F",
    x"1CFE027",
    x"1CFDC2F",
    x"1CFD839",
    x"1CFD443",
    x"1CFD04F",
    x"1CFCC5B",
    x"1CFC868",
    x"1CFC477",
    x"1CFC086",
    x"1CFBC96",
    x"1CFB8A8",
    x"1CFB4BA",
    x"1CFB0CD",
    x"1CFACE2",
    x"1CFA8F7",
    x"1CFA50D",
    x"1CFA124",
    x"1CF9D3D",
    x"1CF9956",
    x"1CF9570",
    x"1CF918B",
    x"1CF8DA7",
    x"1CF89C4",
    x"1CF85E2",
    x"1CF8201",
    x"1CF7E21",
    x"1CF7A42",
    x"1CF7664",
    x"1CF7287",
    x"1CF6EAB",
    x"1CF6AD0",
    x"1CF66F6",
    x"1CF631C",
    x"1CF5F44",
    x"1CF5B6D",
    x"1CF5796",
    x"1CF53C1",
    x"1CF4FEC",
    x"1CF4C19",
    x"1CF4846",
    x"1CF4475",
    x"1CF40A4",
    x"1CF3CD4",
    x"1CF3906",
    x"1CF3538",
    x"1CF316B",
    x"1CF2D9F",
    x"1CF29D4",
    x"1CF260A",
    x"1CF2241",
    x"1CF1E79",
    x"1CF1AB2",
    x"1CF16EC",
    x"1CF1327",
    x"1CF0F62",
    x"1CF0B9F",
    x"1CF07DC",
    x"1CF041B",
    x"1CF005A",
    x"1CEFC9B",
    x"1CEF8DC",
    x"1CEF51E",
    x"1CEF162",
    x"1CEEDA6",
    x"1CEE9EB",
    x"1CEE631",
    x"1CEE278",
    x"1CEDEBF",
    x"1CEDB08",
    x"1CED752",
    x"1CED39D",
    x"1CECFE8",
    x"1CECC35",
    x"1CEC882",
    x"1CEC4D0",
    x"1CEC120",
    x"1CEBD70",
    x"1CEB9C1",
    x"1CEB613",
    x"1CEB266",
    x"1CEAEBA",
    x"1CEAB0E",
    x"1CEA764",
    x"1CEA3BB",
    x"1CEA012",
    x"1CE9C6B",
    x"1CE98C4",
    x"1CE951E",
    x"1CE917A",
    x"1CE8DD6",
    x"1CE8A33",
    x"1CE8691",
    x"1CE82EF",
    x"1CE7F4F",
    x"1CE7BB0",
    x"1CE7811",
    x"1CE7474",
    x"1CE70D7",
    x"1CE6D3B",
    x"1CE69A0",
    x"1CE6606",
    x"1CE626D",
    x"1CE5ED5",
    x"1CE5B3E",
    x"1CE57A8",
    x"1CE5412",
    x"1CE507E",
    x"1CE4CEA",
    x"1CE4957",
    x"1CE45C5",
    x"1CE4234",
    x"1CE3EA4",
    x"1CE3B15",
    x"1CE3787",
    x"1CE33F9",
    x"1CE306D",
    x"1CE2CE1",
    x"1CE2956",
    x"1CE25CC",
    x"1CE2243",
    x"1CE1EBB",
    x"1CE1B34",
    x"1CE17AD",
    x"1CE1428",
    x"1CE10A3",
    x"1CE0D20",
    x"1CE099D",
    x"1CE061B",
    x"1CE029A",
    x"1CDFF1A",
    x"1CDFB9A",
    x"1CDF81C",
    x"1CDF49E",
    x"1CDF121",
    x"1CDEDA6",
    x"1CDEA2B",
    x"1CDE6B1",
    x"1CDE337",
    x"1CDDFBF",
    x"1CDDC47",
    x"1CDD8D1",
    x"1CDD55B",
    x"1CDD1E6",
    x"1CDCE72",
    x"1CDCAFF",
    x"1CDC78D",
    x"1CDC41B",
    x"1CDC0AB",
    x"1CDBD3B",
    x"1CDB9CC",
    x"1CDB65E",
    x"1CDB2F1",
    x"1CDAF84",
    x"1CDAC19",
    x"1CDA8AE",
    x"1CDA545",
    x"1CDA1DC",
    x"1CD9E74",
    x"1CD9B0C",
    x"1CD97A6",
    x"1CD9441",
    x"1CD90DC",
    x"1CD8D78",
    x"1CD8A15",
    x"1CD86B3",
    x"1CD8352",
    x"1CD7FF2",
    x"1CD7C92",
    x"1CD7933",
    x"1CD75D5",
    x"1CD7278",
    x"1CD6F1C",
    x"1CD6BC1",
    x"1CD6866",
    x"1CD650D",
    x"1CD61B4",
    x"1CD5E5C",
    x"1CD5B05",
    x"1CD57AE",
    x"1CD5459",
    x"1CD5104",
    x"1CD4DB0",
    x"1CD4A5D",
    x"1CD470B",
    x"1CD43BA",
    x"1CD4069",
    x"1CD3D19",
    x"1CD39CB",
    x"1CD367D",
    x"1CD332F",
    x"1CD2FE3",
    x"1CD2C97",
    x"1CD294D",
    x"1CD2603",
    x"1CD22BA",
    x"1CD1F71",
    x"1CD1C2A",
    x"1CD18E3",
    x"1CD159E",
    x"1CD1259",
    x"1CD0F14",
    x"1CD0BD1",
    x"1CD088E",
    x"1CD054D",
    x"1CD020C",
    x"1CCFECC",
    x"1CCFB8C",
    x"1CCF84E",
    x"1CCF510",
    x"1CCF1D3",
    x"1CCEE97",
    x"1CCEB5C",
    x"1CCE822",
    x"1CCE4E8",
    x"1CCE1AF",
    x"1CCDE77",
    x"1CCDB40",
    x"1CCD80A",
    x"1CCD4D4",
    x"1CCD19F",
    x"1CCCE6B",
    x"1CCCB38",
    x"1CCC805",
    x"1CCC4D4",
    x"1CCC1A3",
    x"1CCBE73",
    x"1CCBB44",
    x"1CCB815",
    x"1CCB4E8",
    x"1CCB1BB",
    x"1CCAE8F",
    x"1CCAB64",
    x"1CCA839",
    x"1CCA510",
    x"1CCA1E7",
    x"1CC9EBF",
    x"1CC9B97",
    x"1CC9871",
    x"1CC954B",
    x"1CC9226",
    x"1CC8F02",
    x"1CC8BDF",
    x"1CC88BC",
    x"1CC859A",
    x"1CC8279",
    x"1CC7F59",
    x"1CC7C3A",
    x"1CC791B",
    x"1CC75FD",
    x"1CC72E0",
    x"1CC6FC4",
    x"1CC6CA8",
    x"1CC698D",
    x"1CC6673",
    x"1CC635A",
    x"1CC6042",
    x"1CC5D2A",
    x"1CC5A13",
    x"1CC56FD",
    x"1CC53E8",
    x"1CC50D3",
    x"1CC4DBF",
    x"1CC4AAC",
    x"1CC479A",
    x"1CC4488",
    x"1CC4178",
    x"1CC3E68",
    x"1CC3B58",
    x"1CC384A",
    x"1CC353C",
    x"1CC322F",
    x"1CC2F23",
    x"1CC2C18",
    x"1CC290D",
    x"1CC2603",
    x"1CC22FA",
    x"1CC1FF2",
    x"1CC1CEA",
    x"1CC19E3",
    x"1CC16DD",
    x"1CC13D8",
    x"1CC10D3",
    x"1CC0DCF",
    x"1CC0ACC",
    x"1CC07CA",
    x"1CC04C8",
    x"1CC01C8",
    x"1CBFEC8",
    x"1CBFBC8",
    x"1CBF8CA",
    x"1CBF5CC",
    x"1CBF2CF",
    x"1CBEFD2",
    x"1CBECD7",
    x"1CBE9DC",
    x"1CBE6E2",
    x"1CBE3E9",
    x"1CBE0F0",
    x"1CBDDF8",
    x"1CBDB01",
    x"1CBD80B",
    x"1CBD515",
    x"1CBD220",
    x"1CBCF2C",
    x"1CBCC38",
    x"1CBC946",
    x"1CBC654",
    x"1CBC363",
    x"1CBC072",
    x"1CBBD82",
    x"1CBBA93",
    x"1CBB7A5",
    x"1CBB4B8",
    x"1CBB1CB",
    x"1CBAEDF",
    x"1CBABF3",
    x"1CBA909",
    x"1CBA61F",
    x"1CBA336",
    x"1CBA04D",
    x"1CB9D65",
    x"1CB9A7E",
    x"1CB9798",
    x"1CB94B3",
    x"1CB91CE",
    x"1CB8EEA",
    x"1CB8C06",
    x"1CB8924",
    x"1CB8642",
    x"1CB8361",
    x"1CB8080",
    x"1CB7DA0",
    x"1CB7AC1",
    x"1CB77E3",
    x"1CB7505",
    x"1CB7228",
    x"1CB6F4C",
    x"1CB6C71",
    x"1CB6996",
    x"1CB66BC",
    x"1CB63E3",
    x"1CB610A",
    x"1CB5E32",
    x"1CB5B5B",
    x"1CB5884",
    x"1CB55AF",
    x"1CB52DA",
    x"1CB5005",
    x"1CB4D32",
    x"1CB4A5F",
    x"1CB478C",
    x"1CB44BB",
    x"1CB41EA",
    x"1CB3F1A",
    x"1CB3C4B",
    x"1CB397C",
    x"1CB36AE",
    x"1CB33E0",
    x"1CB3114",
    x"1CB2E48",
    x"1CB2B7D",
    x"1CB28B2",
    x"1CB25E8",
    x"1CB231F",
    x"1CB2057",
    x"1CB1D8F",
    x"1CB1AC8",
    x"1CB1802",
    x"1CB153C",
    x"1CB1277",
    x"1CB0FB3",
    x"1CB0CEF",
    x"1CB0A2C",
    x"1CB076A",
    x"1CB04A9",
    x"1CB01E8",
    x"1CAFF28",
    x"1CAFC68",
    x"1CAF9A9",
    x"1CAF6EB",
    x"1CAF42E",
    x"1CAF171",
    x"1CAEEB5",
    x"1CAEBFA",
    x"1CAE93F",
    x"1CAE685",
    x"1CAE3CC",
    x"1CAE113",
    x"1CADE5B",
    x"1CADBA4",
    x"1CAD8EE",
    x"1CAD638",
    x"1CAD383",
    x"1CAD0CE",
    x"1CACE1A",
    x"1CACB67",
    x"1CAC8B4",
    x"1CAC603",
    x"1CAC351",
    x"1CAC0A1",
    x"1CABDF1",
    x"1CABB42",
    x"1CAB893",
    x"1CAB5E6",
    x"1CAB339",
    x"1CAB08C",
    x"1CAADE0",
    x"1CAAB35",
    x"1CAA88B",
    x"1CAA5E1",
    x"1CAA338",
    x"1CAA08F",
    x"1CA9DE7",
    x"1CA9B40",
    x"1CA989A",
    x"1CA95F4",
    x"1CA934F",
    x"1CA90AA",
    x"1CA8E06",
    x"1CA8B63",
    x"1CA88C1",
    x"1CA861F",
    x"1CA837E",
    x"1CA80DD",
    x"1CA7E3D",
    x"1CA7B9E",
    x"1CA78FF",
    x"1CA7662",
    x"1CA73C4",
    x"1CA7128",
    x"1CA6E8C",
    x"1CA6BF0",
    x"1CA6956",
    x"1CA66BC",
    x"1CA6422",
    x"1CA618A",
    x"1CA5EF2",
    x"1CA5C5A",
    x"1CA59C3",
    x"1CA572D",
    x"1CA5498",
    x"1CA5203",
    x"1CA4F6F",
    x"1CA4CDB",
    x"1CA4A48",
    x"1CA47B6",
    x"1CA4525",
    x"1CA4294",
    x"1CA4003",
    x"1CA3D74",
    x"1CA3AE5",
    x"1CA3856",
    x"1CA35C8",
    x"1CA333B",
    x"1CA30AF",
    x"1CA2E23",
    x"1CA2B98",
    x"1CA290D",
    x"1CA2683",
    x"1CA23FA",
    x"1CA2171",
    x"1CA1EE9",
    x"1CA1C62",
    x"1CA19DB",
    x"1CA1755",
    x"1CA14CF",
    x"1CA124A",
    x"1CA0FC6",
    x"1CA0D42",
    x"1CA0ABF",
    x"1CA083D",
    x"1CA05BB",
    x"1CA033A",
    x"1CA00BA",
    x"1C9FE3A",
    x"1C9FBBB",
    x"1C9F93C",
    x"1C9F6BE",
    x"1C9F441",
    x"1C9F1C4",
    x"1C9EF48",
    x"1C9ECCC",
    x"1C9EA51",
    x"1C9E7D7",
    x"1C9E55D",
    x"1C9E2E4",
    x"1C9E06C",
    x"1C9DDF4",
    x"1C9DB7D",
    x"1C9D906",
    x"1C9D690",
    x"1C9D41B",
    x"1C9D1A6",
    x"1C9CF32",
    x"1C9CCBF",
    x"1C9CA4C",
    x"1C9C7DA",
    x"1C9C568",
    x"1C9C2F7",
    x"1C9C087",
    x"1C9BE17",
    x"1C9BBA7",
    x"1C9B939",
    x"1C9B6CB",
    x"1C9B45D",
    x"1C9B1F1",
    x"1C9AF85",
    x"1C9AD19",
    x"1C9AAAE",
    x"1C9A844",
    x"1C9A5DA",
    x"1C9A371",
    x"1C9A108",
    x"1C99EA0",
    x"1C99C39",
    x"1C999D2",
    x"1C9976C",
    x"1C99506",
    x"1C992A1",
    x"1C9903D",
    x"1C98DD9",
    x"1C98B76",
    x"1C98914",
    x"1C986B2",
    x"1C98450",
    x"1C981EF",
    x"1C97F8F",
    x"1C97D30",
    x"1C97AD1",
    x"1C97872",
    x"1C97614",
    x"1C973B7",
    x"1C9715B",
    x"1C96EFE",
    x"1C96CA3",
    x"1C96A48",
    x"1C967EE",
    x"1C96594",
    x"1C9633B",
    x"1C960E3",
    x"1C95E8B",
    x"1C95C33",
    x"1C959DD",
    x"1C95786",
    x"1C95531",
    x"1C952DC",
    x"1C95087",
    x"1C94E34",
    x"1C94BE0",
    x"1C9498E",
    x"1C9473B",
    x"1C944EA",
    x"1C94299",
    x"1C94049",
    x"1C93DF9",
    x"1C93BAA",
    x"1C9395B",
    x"1C9370D",
    x"1C934C0",
    x"1C93273",
    x"1C93026",
    x"1C92DDB",
    x"1C92B8F",
    x"1C92945",
    x"1C926FB",
    x"1C924B1",
    x"1C92268",
    x"1C92020",
    x"1C91DD8",
    x"1C91B91",
    x"1C9194B",
    x"1C91704",
    x"1C914BF",
    x"1C9127A",
    x"1C91036",
    x"1C90DF2",
    x"1C90BAF",
    x"1C9096C",
    x"1C9072A",
    x"1C904E9",
    x"1C902A8",
    x"1C90067",
    x"1C8FE27",
    x"1C8FBE8",
    x"1C8F9A9",
    x"1C8F76B",
    x"1C8F52E",
    x"1C8F2F1",
    x"1C8F0B4",
    x"1C8EE78",
    x"1C8EC3D",
    x"1C8EA02",
    x"1C8E7C8",
    x"1C8E58E",
    x"1C8E355",
    x"1C8E11D",
    x"1C8DEE5",
    x"1C8DCAD",
    x"1C8DA76",
    x"1C8D840",
    x"1C8D60A",
    x"1C8D3D5",
    x"1C8D1A0",
    x"1C8CF6C",
    x"1C8CD39",
    x"1C8CB06",
    x"1C8C8D3",
    x"1C8C6A1",
    x"1C8C470",
    x"1C8C23F",
    x"1C8C00F",
    x"1C8BDDF",
    x"1C8BBB0",
    x"1C8B981",
    x"1C8B753",
    x"1C8B525",
    x"1C8B2F8",
    x"1C8B0CC",
    x"1C8AEA0",
    x"1C8AC75",
    x"1C8AA4A",
    x"1C8A81F",
    x"1C8A5F6",
    x"1C8A3CD",
    x"1C8A1A4",
    x"1C89F7C",
    x"1C89D54",
    x"1C89B2D",
    x"1C89906",
    x"1C896E1",
    x"1C894BB",
    x"1C89296",
    x"1C89072",
    x"1C88E4E",
    x"1C88C2B",
    x"1C88A08",
    x"1C887E6",
    x"1C885C4",
    x"1C883A3",
    x"1C88182",
    x"1C87F62",
    x"1C87D42",
    x"1C87B23",
    x"1C87905",
    x"1C876E7",
    x"1C874C9",
    x"1C872AC",
    x"1C87090",
    x"1C86E74",
    x"1C86C59",
    x"1C86A3E",
    x"1C86824",
    x"1C8660A",
    x"1C863F1",
    x"1C861D8",
    x"1C85FC0",
    x"1C85DA8",
    x"1C85B91",
    x"1C8597A",
    x"1C85764",
    x"1C8554F",
    x"1C85339",
    x"1C85125",
    x"1C84F11",
    x"1C84CFD",
    x"1C84AEA",
    x"1C848D8",
    x"1C846C6",
    x"1C844B5",
    x"1C842A4",
    x"1C84093",
    x"1C83E83",
    x"1C83C74",
    x"1C83A65",
    x"1C83857",
    x"1C83649",
    x"1C8343C",
    x"1C8322F",
    x"1C83023",
    x"1C82E17",
    x"1C82C0C",
    x"1C82A01",
    x"1C827F7",
    x"1C825ED",
    x"1C823E4",
    x"1C821DB",
    x"1C81FD3",
    x"1C81DCB",
    x"1C81BC4",
    x"1C819BD",
    x"1C817B7",
    x"1C815B1",
    x"1C813AC",
    x"1C811A7",
    x"1C80FA3",
    x"1C80DA0",
    x"1C80B9C",
    x"1C8099A",
    x"1C80798",
    x"1C80596",
    x"1C80395",
    x"1C80194",
    x"1C7FF28",
    x"1C7FB29",
    x"1C7F72B",
    x"1C7F32E",
    x"1C7EF31",
    x"1C7EB36",
    x"1C7E73C",
    x"1C7E342",
    x"1C7DF4A",
    x"1C7DB53",
    x"1C7D75C",
    x"1C7D367",
    x"1C7CF73",
    x"1C7CB7F",
    x"1C7C78D",
    x"1C7C39B",
    x"1C7BFAB",
    x"1C7BBBC",
    x"1C7B7CD",
    x"1C7B3E0",
    x"1C7AFF3",
    x"1C7AC08",
    x"1C7A81D",
    x"1C7A434",
    x"1C7A04B",
    x"1C79C64",
    x"1C7987D",
    x"1C79497",
    x"1C790B3",
    x"1C78CCF",
    x"1C788EC",
    x"1C7850B",
    x"1C7812A",
    x"1C77D4A",
    x"1C7796B",
    x"1C7758D",
    x"1C771B0",
    x"1C76DD4",
    x"1C769F9",
    x"1C7661F",
    x"1C76246",
    x"1C75E6E",
    x"1C75A97",
    x"1C756C1",
    x"1C752EC",
    x"1C74F17",
    x"1C74B44",
    x"1C74772",
    x"1C743A0",
    x"1C73FD0",
    x"1C73C01",
    x"1C73832",
    x"1C73464",
    x"1C73098",
    x"1C72CCC",
    x"1C72901",
    x"1C72538",
    x"1C7216F",
    x"1C71DA7",
    x"1C719E0",
    x"1C7161A",
    x"1C71255",
    x"1C70E91",
    x"1C70ACE",
    x"1C7070B",
    x"1C7034A",
    x"1C6FF8A",
    x"1C6FBCA",
    x"1C6F80C",
    x"1C6F44E",
    x"1C6F092",
    x"1C6ECD6",
    x"1C6E91B",
    x"1C6E562",
    x"1C6E1A9",
    x"1C6DDF1",
    x"1C6DA3A",
    x"1C6D684",
    x"1C6D2CE",
    x"1C6CF1A",
    x"1C6CB67",
    x"1C6C7B4",
    x"1C6C403",
    x"1C6C052",
    x"1C6BCA3",
    x"1C6B8F4",
    x"1C6B546",
    x"1C6B199",
    x"1C6ADEE",
    x"1C6AA43",
    x"1C6A698",
    x"1C6A2EF",
    x"1C69F47",
    x"1C69BA0",
    x"1C697F9",
    x"1C69454",
    x"1C690AF",
    x"1C68D0B",
    x"1C68968",
    x"1C685C7",
    x"1C68226",
    x"1C67E85",
    x"1C67AE6",
    x"1C67748",
    x"1C673AB",
    x"1C6700E",
    x"1C66C73",
    x"1C668D8",
    x"1C6653E",
    x"1C661A5",
    x"1C65E0D",
    x"1C65A76",
    x"1C656E0",
    x"1C6534B",
    x"1C64FB7",
    x"1C64C23",
    x"1C64890",
    x"1C644FF",
    x"1C6416E",
    x"1C63DDE",
    x"1C63A4F",
    x"1C636C1",
    x"1C63334",
    x"1C62FA7",
    x"1C62C1C",
    x"1C62891",
    x"1C62508",
    x"1C6217F",
    x"1C61DF7",
    x"1C61A70",
    x"1C616EA",
    x"1C61364",
    x"1C60FE0",
    x"1C60C5C",
    x"1C608DA",
    x"1C60558",
    x"1C601D7",
    x"1C5FE57",
    x"1C5FAD8",
    x"1C5F75A",
    x"1C5F3DC",
    x"1C5F060",
    x"1C5ECE4",
    x"1C5E969",
    x"1C5E5EF",
    x"1C5E276",
    x"1C5DEFE",
    x"1C5DB87",
    x"1C5D810",
    x"1C5D49B",
    x"1C5D126",
    x"1C5CDB2",
    x"1C5CA3F",
    x"1C5C6CD",
    x"1C5C35C",
    x"1C5BFEB",
    x"1C5BC7C",
    x"1C5B90D",
    x"1C5B59F",
    x"1C5B232",
    x"1C5AEC6",
    x"1C5AB5B",
    x"1C5A7F0",
    x"1C5A487",
    x"1C5A11E",
    x"1C59DB6",
    x"1C59A4F",
    x"1C596E9",
    x"1C59384",
    x"1C5901F",
    x"1C58CBC",
    x"1C58959",
    x"1C585F7",
    x"1C58296",
    x"1C57F36",
    x"1C57BD6",
    x"1C57878",
    x"1C5751A",
    x"1C571BD",
    x"1C56E61",
    x"1C56B06",
    x"1C567AC",
    x"1C56452",
    x"1C560FA",
    x"1C55DA2",
    x"1C55A4B",
    x"1C556F5",
    x"1C5539F",
    x"1C5504B",
    x"1C54CF7",
    x"1C549A4",
    x"1C54652",
    x"1C54301",
    x"1C53FB1",
    x"1C53C61",
    x"1C53913",
    x"1C535C5",
    x"1C53278",
    x"1C52F2C",
    x"1C52BE0",
    x"1C52896",
    x"1C5254C",
    x"1C52203",
    x"1C51EBB",
    x"1C51B74",
    x"1C5182D",
    x"1C514E8",
    x"1C511A3",
    x"1C50E5F",
    x"1C50B1C",
    x"1C507D9",
    x"1C50498",
    x"1C50157",
    x"1C4FE17",
    x"1C4FAD8",
    x"1C4F79A",
    x"1C4F45C",
    x"1C4F11F",
    x"1C4EDE3",
    x"1C4EAA8",
    x"1C4E76E",
    x"1C4E435",
    x"1C4E0FC",
    x"1C4DDC4",
    x"1C4DA8D",
    x"1C4D757",
    x"1C4D421",
    x"1C4D0ED",
    x"1C4CDB9",
    x"1C4CA86",
    x"1C4C754",
    x"1C4C422",
    x"1C4C0F2",
    x"1C4BDC2",
    x"1C4BA93",
    x"1C4B765",
    x"1C4B437",
    x"1C4B10A",
    x"1C4ADDF",
    x"1C4AAB4",
    x"1C4A789",
    x"1C4A460",
    x"1C4A137",
    x"1C49E0F",
    x"1C49AE8",
    x"1C497C2",
    x"1C4949C",
    x"1C49177",
    x"1C48E53",
    x"1C48B30",
    x"1C4880E",
    x"1C484EC",
    x"1C481CB",
    x"1C47EAB",
    x"1C47B8C",
    x"1C4786E",
    x"1C47550",
    x"1C47233",
    x"1C46F17",
    x"1C46BFB",
    x"1C468E1",
    x"1C465C7",
    x"1C462AE",
    x"1C45F96",
    x"1C45C7E",
    x"1C45967",
    x"1C45651",
    x"1C4533C",
    x"1C45028",
    x"1C44D14",
    x"1C44A01",
    x"1C446EF",
    x"1C443DE",
    x"1C440CD",
    x"1C43DBD",
    x"1C43AAE",
    x"1C437A0",
    x"1C43492",
    x"1C43186",
    x"1C42E7A",
    x"1C42B6E",
    x"1C42864",
    x"1C4255A",
    x"1C42251",
    x"1C41F49",
    x"1C41C42",
    x"1C4193B",
    x"1C41635",
    x"1C41330",
    x"1C4102B",
    x"1C40D28",
    x"1C40A25",
    x"1C40723",
    x"1C40421",
    x"1C40121",
    x"1C3FE21",
    x"1C3FB22",
    x"1C3F823",
    x"1C3F525",
    x"1C3F229",
    x"1C3EF2C",
    x"1C3EC31",
    x"1C3E936",
    x"1C3E63C",
    x"1C3E343",
    x"1C3E04B",
    x"1C3DD53",
    x"1C3DA5C",
    x"1C3D766",
    x"1C3D470",
    x"1C3D17C",
    x"1C3CE88",
    x"1C3CB94",
    x"1C3C8A2",
    x"1C3C5B0",
    x"1C3C2BF",
    x"1C3BFCF",
    x"1C3BCDF",
    x"1C3B9F0",
    x"1C3B702",
    x"1C3B415",
    x"1C3B128",
    x"1C3AE3C",
    x"1C3AB51",
    x"1C3A866",
    x"1C3A57D",
    x"1C3A294",
    x"1C39FAB",
    x"1C39CC4",
    x"1C399DD",
    x"1C396F7",
    x"1C39412",
    x"1C3912D",
    x"1C38E49",
    x"1C38B66",
    x"1C38883",
    x"1C385A2",
    x"1C382C0",
    x"1C37FE0",
    x"1C37D01",
    x"1C37A22",
    x"1C37743",
    x"1C37466",
    x"1C37189",
    x"1C36EAD",
    x"1C36BD2",
    x"1C368F7",
    x"1C3661D",
    x"1C36344",
    x"1C3606C",
    x"1C35D94",
    x"1C35ABD",
    x"1C357E7",
    x"1C35511",
    x"1C3523C",
    x"1C34F68",
    x"1C34C94",
    x"1C349C2",
    x"1C346F0",
    x"1C3441E",
    x"1C3414E",
    x"1C33E7E",
    x"1C33BAE",
    x"1C338E0",
    x"1C33612",
    x"1C33345",
    x"1C33078",
    x"1C32DAC",
    x"1C32AE1",
    x"1C32817",
    x"1C3254D",
    x"1C32284",
    x"1C31FBC",
    x"1C31CF4",
    x"1C31A2E",
    x"1C31767",
    x"1C314A2",
    x"1C311DD",
    x"1C30F19",
    x"1C30C56",
    x"1C30993",
    x"1C306D1",
    x"1C3040F",
    x"1C3014F",
    x"1C2FE8F",
    x"1C2FBCF",
    x"1C2F911",
    x"1C2F653",
    x"1C2F396",
    x"1C2F0D9",
    x"1C2EE1D",
    x"1C2EB62",
    x"1C2E8A8",
    x"1C2E5EE",
    x"1C2E335",
    x"1C2E07C",
    x"1C2DDC4",
    x"1C2DB0D",
    x"1C2D857",
    x"1C2D5A1",
    x"1C2D2EC",
    x"1C2D038",
    x"1C2CD84",
    x"1C2CAD1",
    x"1C2C81E",
    x"1C2C56D",
    x"1C2C2BC",
    x"1C2C00B",
    x"1C2BD5C",
    x"1C2BAAD",
    x"1C2B7FE",
    x"1C2B551",
    x"1C2B2A4",
    x"1C2AFF7",
    x"1C2AD4C",
    x"1C2AAA1",
    x"1C2A7F6",
    x"1C2A54D",
    x"1C2A2A4",
    x"1C29FFB",
    x"1C29D54",
    x"1C29AAD",
    x"1C29806",
    x"1C29561",
    x"1C292BC",
    x"1C29017",
    x"1C28D74",
    x"1C28AD1",
    x"1C2882E",
    x"1C2858D",
    x"1C282EC",
    x"1C2804B",
    x"1C27DAB",
    x"1C27B0C",
    x"1C2786E",
    x"1C275D0",
    x"1C27333",
    x"1C27096",
    x"1C26DFB",
    x"1C26B5F",
    x"1C268C5",
    x"1C2662B",
    x"1C26392",
    x"1C260F9",
    x"1C25E61",
    x"1C25BCA",
    x"1C25933",
    x"1C2569E",
    x"1C25408",
    x"1C25174",
    x"1C24EDF",
    x"1C24C4C",
    x"1C249B9",
    x"1C24727",
    x"1C24496",
    x"1C24205",
    x"1C23F75",
    x"1C23CE5",
    x"1C23A56",
    x"1C237C8",
    x"1C2353A",
    x"1C232AD",
    x"1C23021",
    x"1C22D95",
    x"1C22B0A",
    x"1C22880",
    x"1C225F6",
    x"1C2236D",
    x"1C220E4",
    x"1C21E5C",
    x"1C21BD5",
    x"1C2194E",
    x"1C216C8",
    x"1C21443",
    x"1C211BE",
    x"1C20F3A",
    x"1C20CB7",
    x"1C20A34",
    x"1C207B2",
    x"1C20530",
    x"1C202AF",
    x"1C2002F",
    x"1C1FDAF",
    x"1C1FB30",
    x"1C1F8B1",
    x"1C1F633",
    x"1C1F3B6",
    x"1C1F13A",
    x"1C1EEBE",
    x"1C1EC42",
    x"1C1E9C7",
    x"1C1E74D",
    x"1C1E4D4",
    x"1C1E25B",
    x"1C1DFE3",
    x"1C1DD6B",
    x"1C1DAF4",
    x"1C1D87E",
    x"1C1D608",
    x"1C1D392",
    x"1C1D11E",
    x"1C1CEAA",
    x"1C1CC37",
    x"1C1C9C4",
    x"1C1C752",
    x"1C1C4E0",
    x"1C1C26F",
    x"1C1BFFF",
    x"1C1BD8F",
    x"1C1BB20",
    x"1C1B8B2",
    x"1C1B644",
    x"1C1B3D7",
    x"1C1B16A",
    x"1C1AEFE",
    x"1C1AC92",
    x"1C1AA28",
    x"1C1A7BD",
    x"1C1A554",
    x"1C1A2EB",
    x"1C1A082",
    x"1C19E1A",
    x"1C19BB3",
    x"1C1994D",
    x"1C196E7",
    x"1C19481",
    x"1C1921C",
    x"1C18FB8",
    x"1C18D54",
    x"1C18AF1",
    x"1C1888F",
    x"1C1862D",
    x"1C183CC",
    x"1C1816B",
    x"1C17F0B",
    x"1C17CAC",
    x"1C17A4D",
    x"1C177EF",
    x"1C17591",
    x"1C17334",
    x"1C170D7",
    x"1C16E7B",
    x"1C16C20",
    x"1C169C5",
    x"1C1676B",
    x"1C16512",
    x"1C162B9",
    x"1C16060",
    x"1C15E08",
    x"1C15BB1",
    x"1C1595B",
    x"1C15704",
    x"1C154AF",
    x"1C1525A",
    x"1C15006",
    x"1C14DB2",
    x"1C14B5F",
    x"1C1490C",
    x"1C146BA",
    x"1C14469",
    x"1C14218",
    x"1C13FC8",
    x"1C13D78",
    x"1C13B29",
    x"1C138DB",
    x"1C1368D",
    x"1C13440",
    x"1C131F3",
    x"1C12FA7",
    x"1C12D5B",
    x"1C12B10",
    x"1C128C5",
    x"1C1267B",
    x"1C12432",
    x"1C121E9",
    x"1C11FA1",
    x"1C11D5A",
    x"1C11B13",
    x"1C118CC",
    x"1C11686",
    x"1C11441",
    x"1C111FC",
    x"1C10FB8",
    x"1C10D74",
    x"1C10B31",
    x"1C108EF",
    x"1C106AD",
    x"1C1046B",
    x"1C1022A",
    x"1C0FFEA",
    x"1C0FDAA",
    x"1C0FB6B",
    x"1C0F92D",
    x"1C0F6EF",
    x"1C0F4B1",
    x"1C0F274",
    x"1C0F038",
    x"1C0EDFC",
    x"1C0EBC1",
    x"1C0E986",
    x"1C0E74C",
    x"1C0E513",
    x"1C0E2DA",
    x"1C0E0A1",
    x"1C0DE69",
    x"1C0DC32",
    x"1C0D9FB",
    x"1C0D7C5",
    x"1C0D58F",
    x"1C0D35A",
    x"1C0D126",
    x"1C0CEF2",
    x"1C0CCBE",
    x"1C0CA8B",
    x"1C0C859",
    x"1C0C627",
    x"1C0C3F6",
    x"1C0C1C5",
    x"1C0BF95",
    x"1C0BD65",
    x"1C0BB36",
    x"1C0B908",
    x"1C0B6DA",
    x"1C0B4AC",
    x"1C0B27F",
    x"1C0B053",
    x"1C0AE27",
    x"1C0ABFC",
    x"1C0A9D1",
    x"1C0A7A7",
    x"1C0A57D",
    x"1C0A354",
    x"1C0A12C",
    x"1C09F04",
    x"1C09CDC",
    x"1C09AB5",
    x"1C0988F",
    x"1C09669",
    x"1C09444",
    x"1C0921F",
    x"1C08FFB",
    x"1C08DD7",
    x"1C08BB4",
    x"1C08991",
    x"1C0876F",
    x"1C0854D",
    x"1C0832C",
    x"1C0810C",
    x"1C07EEC",
    x"1C07CCC",
    x"1C07AAD",
    x"1C0788F",
    x"1C07671",
    x"1C07454",
    x"1C07237",
    x"1C0701B",
    x"1C06DFF",
    x"1C06BE4",
    x"1C069C9",
    x"1C067AF",
    x"1C06595",
    x"1C0637C",
    x"1C06163",
    x"1C05F4B",
    x"1C05D34",
    x"1C05B1D",
    x"1C05906",
    x"1C056F0",
    x"1C054DB",
    x"1C052C6",
    x"1C050B1",
    x"1C04E9D",
    x"1C04C8A",
    x"1C04A77",
    x"1C04865",
    x"1C04653",
    x"1C04442",
    x"1C04231",
    x"1C04020",
    x"1C03E11",
    x"1C03C01",
    x"1C039F3",
    x"1C037E4",
    x"1C035D7",
    x"1C033CA",
    x"1C031BD",
    x"1C02FB1",
    x"1C02DA5",
    x"1C02B9A",
    x"1C0298F",
    x"1C02785",
    x"1C0257B",
    x"1C02372",
    x"1C0216A",
    x"1C01F62",
    x"1C01D5A",
    x"1C01B53",
    x"1C0194C",
    x"1C01746",
    x"1C01541",
    x"1C0133C",
    x"1C01137",
    x"1C00F33",
    x"1C00D30",
    x"1C00B2C",
    x"1C0092A",
    x"1C00728",
    x"1C00526",
    x"1C00325",
    x"1C00125",
    x"1BFFE4A",
    x"1BFFA4B",
    x"1BFF64D",
    x"1BFF250",
    x"1BFEE54",
    x"1BFEA59",
    x"1BFE65F",
    x"1BFE265",
    x"1BFDE6D",
    x"1BFDA76",
    x"1BFD680",
    x"1BFD28B",
    x"1BFCE97",
    x"1BFCAA4",
    x"1BFC6B1",
    x"1BFC2C0",
    x"1BFBED0",
    x"1BFBAE1",
    x"1BFB6F3",
    x"1BFB305",
    x"1BFAF19",
    x"1BFAB2E",
    x"1BFA744",
    x"1BFA35A",
    x"1BF9F72",
    x"1BF9B8B",
    x"1BF97A4",
    x"1BF93BF",
    x"1BF8FDA",
    x"1BF8BF7",
    x"1BF8814",
    x"1BF8433",
    x"1BF8052",
    x"1BF7C73",
    x"1BF7894",
    x"1BF74B6",
    x"1BF70DA",
    x"1BF6CFE",
    x"1BF6923",
    x"1BF6549",
    x"1BF6170",
    x"1BF5D99",
    x"1BF59C2",
    x"1BF55EC",
    x"1BF5217",
    x"1BF4E43",
    x"1BF4A70",
    x"1BF469D",
    x"1BF42CC",
    x"1BF3EFC",
    x"1BF3B2D",
    x"1BF375E",
    x"1BF3391",
    x"1BF2FC5",
    x"1BF2BF9",
    x"1BF282F",
    x"1BF2465",
    x"1BF209C",
    x"1BF1CD5",
    x"1BF190E",
    x"1BF1548",
    x"1BF1183",
    x"1BF0DBF",
    x"1BF09FD",
    x"1BF063A",
    x"1BF0279",
    x"1BEFEB9",
    x"1BEFAFA",
    x"1BEF73C",
    x"1BEF37E",
    x"1BEEFC2",
    x"1BEEC07",
    x"1BEE84C",
    x"1BEE492",
    x"1BEE0DA",
    x"1BEDD22",
    x"1BED96B",
    x"1BED5B5",
    x"1BED200",
    x"1BECE4C",
    x"1BECA99",
    x"1BEC6E7",
    x"1BEC336",
    x"1BEBF85",
    x"1BEBBD6",
    x"1BEB827",
    x"1BEB47A",
    x"1BEB0CD",
    x"1BEAD21",
    x"1BEA977",
    x"1BEA5CD",
    x"1BEA224",
    x"1BE9E7C",
    x"1BE9AD4",
    x"1BE972E",
    x"1BE9389",
    x"1BE8FE4",
    x"1BE8C41",
    x"1BE889E",
    x"1BE84FD",
    x"1BE815C",
    x"1BE7DBC",
    x"1BE7A1D",
    x"1BE767F",
    x"1BE72E2",
    x"1BE6F45",
    x"1BE6BAA",
    x"1BE6810",
    x"1BE6476",
    x"1BE60DD",
    x"1BE5D46",
    x"1BE59AF",
    x"1BE5619",
    x"1BE5284",
    x"1BE4EF0",
    x"1BE4B5C",
    x"1BE47CA",
    x"1BE4438",
    x"1BE40A8",
    x"1BE3D18",
    x"1BE3989",
    x"1BE35FB",
    x"1BE326E",
    x"1BE2EE2",
    x"1BE2B57",
    x"1BE27CC",
    x"1BE2443",
    x"1BE20BA",
    x"1BE1D32",
    x"1BE19AC",
    x"1BE1626",
    x"1BE12A1",
    x"1BE0F1C",
    x"1BE0B99",
    x"1BE0817",
    x"1BE0495",
    x"1BE0114",
    x"1BDFD94",
    x"1BDFA15",
    x"1BDF697",
    x"1BDF31A",
    x"1BDEF9E",
    x"1BDEC22",
    x"1BDE8A8",
    x"1BDE52E",
    x"1BDE1B5",
    x"1BDDE3D",
    x"1BDDAC6",
    x"1BDD750",
    x"1BDD3DA",
    x"1BDD066",
    x"1BDCCF2",
    x"1BDC97F",
    x"1BDC60D",
    x"1BDC29C",
    x"1BDBF2C",
    x"1BDBBBD",
    x"1BDB84E",
    x"1BDB4E1",
    x"1BDB174",
    x"1BDAE08",
    x"1BDAA9D",
    x"1BDA733",
    x"1BDA3C9",
    x"1BDA061",
    x"1BD9CF9",
    x"1BD9992",
    x"1BD962C",
    x"1BD92C7",
    x"1BD8F63",
    x"1BD8BFF",
    x"1BD889D",
    x"1BD853B",
    x"1BD81DA",
    x"1BD7E7A",
    x"1BD7B1B",
    x"1BD77BD",
    x"1BD745F",
    x"1BD7102",
    x"1BD6DA7",
    x"1BD6A4C",
    x"1BD66F1",
    x"1BD6398",
    x"1BD6040",
    x"1BD5CE8",
    x"1BD5991",
    x"1BD563B",
    x"1BD52E6",
    x"1BD4F92",
    x"1BD4C3E",
    x"1BD48EC",
    x"1BD459A",
    x"1BD4249",
    x"1BD3EF9",
    x"1BD3BA9",
    x"1BD385B",
    x"1BD350D",
    x"1BD31C0",
    x"1BD2E74",
    x"1BD2B29",
    x"1BD27DF",
    x"1BD2495",
    x"1BD214C",
    x"1BD1E04",
    x"1BD1ABD",
    x"1BD1777",
    x"1BD1432",
    x"1BD10ED",
    x"1BD0DA9",
    x"1BD0A66",
    x"1BD0724",
    x"1BD03E3",
    x"1BD00A2",
    x"1BCFD62",
    x"1BCFA23",
    x"1BCF6E5",
    x"1BCF3A8",
    x"1BCF06B",
    x"1BCED30",
    x"1BCE9F5",
    x"1BCE6BB",
    x"1BCE381",
    x"1BCE049",
    x"1BCDD11",
    x"1BCD9DA",
    x"1BCD6A4",
    x"1BCD36F",
    x"1BCD03B",
    x"1BCCD07",
    x"1BCC9D4",
    x"1BCC6A2",
    x"1BCC371",
    x"1BCC040",
    x"1BCBD11",
    x"1BCB9E2",
    x"1BCB6B4",
    x"1BCB386",
    x"1BCB05A",
    x"1BCAD2E",
    x"1BCAA03",
    x"1BCA6D9",
    x"1BCA3B0",
    x"1BCA087",
    x"1BC9D60",
    x"1BC9A39",
    x"1BC9713",
    x"1BC93ED",
    x"1BC90C9",
    x"1BC8DA5",
    x"1BC8A82",
    x"1BC8760",
    x"1BC843E",
    x"1BC811D",
    x"1BC7DFE",
    x"1BC7ADE",
    x"1BC77C0",
    x"1BC74A3",
    x"1BC7186",
    x"1BC6E6A",
    x"1BC6B4F",
    x"1BC6834",
    x"1BC651A",
    x"1BC6202",
    x"1BC5EE9",
    x"1BC5BD2",
    x"1BC58BC",
    x"1BC55A6",
    x"1BC5291",
    x"1BC4F7C",
    x"1BC4C69",
    x"1BC4956",
    x"1BC4644",
    x"1BC4333",
    x"1BC4023",
    x"1BC3D13",
    x"1BC3A04",
    x"1BC36F6",
    x"1BC33E9",
    x"1BC30DC",
    x"1BC2DD0",
    x"1BC2AC5",
    x"1BC27BB",
    x"1BC24B1",
    x"1BC21A9",
    x"1BC1EA1",
    x"1BC1B99",
    x"1BC1893",
    x"1BC158D",
    x"1BC1288",
    x"1BC0F84",
    x"1BC0C80",
    x"1BC097D",
    x"1BC067B",
    x"1BC037A",
    x"1BC007A",
    x"1BBFD7A",
    x"1BBFA7B",
    x"1BBF77D",
    x"1BBF47F",
    x"1BBF182",
    x"1BBEE86",
    x"1BBEB8B",
    x"1BBE891",
    x"1BBE597",
    x"1BBE29E",
    x"1BBDFA6",
    x"1BBDCAE",
    x"1BBD9B7",
    x"1BBD6C1",
    x"1BBD3CC",
    x"1BBD0D7",
    x"1BBCDE3",
    x"1BBCAF0",
    x"1BBC7FE",
    x"1BBC50C",
    x"1BBC21B",
    x"1BBBF2B",
    x"1BBBC3C",
    x"1BBB94D",
    x"1BBB65F",
    x"1BBB372",
    x"1BBB086",
    x"1BBAD9A",
    x"1BBAAAF",
    x"1BBA7C4",
    x"1BBA4DB",
    x"1BBA1F2",
    x"1BB9F0A",
    x"1BB9C22",
    x"1BB993C",
    x"1BB9656",
    x"1BB9371",
    x"1BB908C",
    x"1BB8DA8",
    x"1BB8AC5",
    x"1BB87E3",
    x"1BB8501",
    x"1BB8220",
    x"1BB7F40",
    x"1BB7C61",
    x"1BB7982",
    x"1BB76A4",
    x"1BB73C7",
    x"1BB70EA",
    x"1BB6E0E",
    x"1BB6B33",
    x"1BB6859",
    x"1BB657F",
    x"1BB62A6",
    x"1BB5FCE",
    x"1BB5CF6",
    x"1BB5A1F",
    x"1BB5749",
    x"1BB5474",
    x"1BB519F",
    x"1BB4ECB",
    x"1BB4BF7",
    x"1BB4925",
    x"1BB4653",
    x"1BB4382",
    x"1BB40B1",
    x"1BB3DE1",
    x"1BB3B12",
    x"1BB3844",
    x"1BB3576",
    x"1BB32A9",
    x"1BB2FDD",
    x"1BB2D11",
    x"1BB2A46",
    x"1BB277C",
    x"1BB24B2",
    x"1BB21EA",
    x"1BB1F21",
    x"1BB1C5A",
    x"1BB1993",
    x"1BB16CD",
    x"1BB1408",
    x"1BB1143",
    x"1BB0E7F",
    x"1BB0BBC",
    x"1BB08F9",
    x"1BB0637",
    x"1BB0376",
    x"1BB00B6",
    x"1BAFDF6",
    x"1BAFB37",
    x"1BAF878",
    x"1BAF5BA",
    x"1BAF2FD",
    x"1BAF041",
    x"1BAED85",
    x"1BAEACA",
    x"1BAE810",
    x"1BAE556",
    x"1BAE29D",
    x"1BADFE5",
    x"1BADD2D",
    x"1BADA76",
    x"1BAD7C0",
    x"1BAD50A",
    x"1BAD255",
    x"1BACFA1",
    x"1BACCEE",
    x"1BACA3B",
    x"1BAC789",
    x"1BAC4D7",
    x"1BAC226",
    x"1BABF76",
    x"1BABCC6",
    x"1BABA18",
    x"1BAB769",
    x"1BAB4BC",
    x"1BAB20F",
    x"1BAAF63",
    x"1BAACB7",
    x"1BAAA0C",
    x"1BAA762",
    x"1BAA4B9",
    x"1BAA210",
    x"1BA9F68",
    x"1BA9CC0",
    x"1BA9A19",
    x"1BA9773",
    x"1BA94CE",
    x"1BA9229",
    x"1BA8F85",
    x"1BA8CE1",
    x"1BA8A3E",
    x"1BA879C",
    x"1BA84FA",
    x"1BA8259",
    x"1BA7FB9",
    x"1BA7D1A",
    x"1BA7A7B",
    x"1BA77DC",
    x"1BA753F",
    x"1BA72A2",
    x"1BA7005",
    x"1BA6D6A",
    x"1BA6ACF",
    x"1BA6834",
    x"1BA659B",
    x"1BA6301",
    x"1BA6069",
    x"1BA5DD1",
    x"1BA5B3A",
    x"1BA58A4",
    x"1BA560E",
    x"1BA5379",
    x"1BA50E4",
    x"1BA4E50",
    x"1BA4BBD",
    x"1BA492A",
    x"1BA4698",
    x"1BA4407",
    x"1BA4176",
    x"1BA3EE6",
    x"1BA3C57",
    x"1BA39C8",
    x"1BA373A",
    x"1BA34AC",
    x"1BA3220",
    x"1BA2F93",
    x"1BA2D08",
    x"1BA2A7D",
    x"1BA27F3",
    x"1BA2569",
    x"1BA22E0",
    x"1BA2057",
    x"1BA1DD0",
    x"1BA1B49",
    x"1BA18C2",
    x"1BA163C",
    x"1BA13B7",
    x"1BA1132",
    x"1BA0EAE",
    x"1BA0C2B",
    x"1BA09A8",
    x"1BA0726",
    x"1BA04A5",
    x"1BA0224",
    x"1B9FFA4",
    x"1B9FD24",
    x"1B9FAA5",
    x"1B9F827",
    x"1B9F5A9",
    x"1B9F32C",
    x"1B9F0AF",
    x"1B9EE33",
    x"1B9EBB8",
    x"1B9E93E",
    x"1B9E6C4",
    x"1B9E44A",
    x"1B9E1D1",
    x"1B9DF59",
    x"1B9DCE2",
    x"1B9DA6B",
    x"1B9D7F5",
    x"1B9D57F",
    x"1B9D30A",
    x"1B9D095",
    x"1B9CE22",
    x"1B9CBAE",
    x"1B9C93C",
    x"1B9C6CA",
    x"1B9C458",
    x"1B9C1E8",
    x"1B9BF77",
    x"1B9BD08",
    x"1B9BA99",
    x"1B9B82B",
    x"1B9B5BD",
    x"1B9B350",
    x"1B9B0E3",
    x"1B9AE77",
    x"1B9AC0C",
    x"1B9A9A1",
    x"1B9A737",
    x"1B9A4CE",
    x"1B9A265",
    x"1B99FFC",
    x"1B99D95",
    x"1B99B2E",
    x"1B998C7",
    x"1B99661",
    x"1B993FC",
    x"1B99197",
    x"1B98F33",
    x"1B98CD0",
    x"1B98A6D",
    x"1B9880A",
    x"1B985A9",
    x"1B98348",
    x"1B980E7",
    x"1B97E87",
    x"1B97C28",
    x"1B979C9",
    x"1B9776B",
    x"1B9750D",
    x"1B972B0",
    x"1B97054",
    x"1B96DF8",
    x"1B96B9D",
    x"1B96942",
    x"1B966E8",
    x"1B9648F",
    x"1B96236",
    x"1B95FDE",
    x"1B95D86",
    x"1B95B2F",
    x"1B958D9",
    x"1B95683",
    x"1B9542D",
    x"1B951D9",
    x"1B94F84",
    x"1B94D31",
    x"1B94ADE",
    x"1B9488B",
    x"1B94639",
    x"1B943E8",
    x"1B94198",
    x"1B93F47",
    x"1B93CF8",
    x"1B93AA9",
    x"1B9385B",
    x"1B9360D",
    x"1B933C0",
    x"1B93173",
    x"1B92F27",
    x"1B92CDB",
    x"1B92A90",
    x"1B92846",
    x"1B925FC",
    x"1B923B3",
    x"1B9216A",
    x"1B91F22",
    x"1B91CDB",
    x"1B91A94",
    x"1B9184E",
    x"1B91608",
    x"1B913C3",
    x"1B9117E",
    x"1B90F3A",
    x"1B90CF6",
    x"1B90AB3",
    x"1B90871",
    x"1B9062F",
    x"1B903EE",
    x"1B901AD",
    x"1B8FF6D",
    x"1B8FD2D",
    x"1B8FAEE",
    x"1B8F8B0",
    x"1B8F672",
    x"1B8F435",
    x"1B8F1F8",
    x"1B8EFBC",
    x"1B8ED80",
    x"1B8EB45",
    x"1B8E90A",
    x"1B8E6D0",
    x"1B8E497",
    x"1B8E25E",
    x"1B8E026",
    x"1B8DDEE",
    x"1B8DBB7",
    x"1B8D980",
    x"1B8D74A",
    x"1B8D515",
    x"1B8D2E0",
    x"1B8D0AB",
    x"1B8CE77",
    x"1B8CC44",
    x"1B8CA11",
    x"1B8C7DF",
    x"1B8C5AD",
    x"1B8C37C",
    x"1B8C14B",
    x"1B8BF1B",
    x"1B8BCEC",
    x"1B8BABD",
    x"1B8B88E",
    x"1B8B661",
    x"1B8B433",
    x"1B8B207",
    x"1B8AFDA",
    x"1B8ADAF",
    x"1B8AB83",
    x"1B8A959",
    x"1B8A72F",
    x"1B8A505",
    x"1B8A2DC",
    x"1B8A0B4",
    x"1B89E8C",
    x"1B89C65",
    x"1B89A3E",
    x"1B89817",
    x"1B895F2",
    x"1B893CC",
    x"1B891A8",
    x"1B88F84",
    x"1B88D60",
    x"1B88B3D",
    x"1B8891A",
    x"1B886F8",
    x"1B884D7",
    x"1B882B6",
    x"1B88096",
    x"1B87E76",
    x"1B87C56",
    x"1B87A37",
    x"1B87819",
    x"1B875FB",
    x"1B873DE",
    x"1B871C2",
    x"1B86FA5",
    x"1B86D8A",
    x"1B86B6F",
    x"1B86954",
    x"1B8673A",
    x"1B86520",
    x"1B86307",
    x"1B860EF",
    x"1B85ED7",
    x"1B85CBF",
    x"1B85AA8",
    x"1B85892",
    x"1B8567C",
    x"1B85467",
    x"1B85252",
    x"1B8503E",
    x"1B84E2A",
    x"1B84C17",
    x"1B84A04",
    x"1B847F2",
    x"1B845E0",
    x"1B843CF",
    x"1B841BE",
    x"1B83FAE",
    x"1B83D9E",
    x"1B83B8F",
    x"1B83980",
    x"1B83772",
    x"1B83565",
    x"1B83358",
    x"1B8314B",
    x"1B82F3F",
    x"1B82D33",
    x"1B82B28",
    x"1B8291E",
    x"1B82714",
    x"1B8250A",
    x"1B82301",
    x"1B820F9",
    x"1B81EF1",
    x"1B81CE9",
    x"1B81AE2",
    x"1B818DC",
    x"1B816D6",
    x"1B814D0",
    x"1B812CB",
    x"1B810C7",
    x"1B80EC3",
    x"1B80CC0",
    x"1B80ABD",
    x"1B808BA",
    x"1B806B8",
    x"1B804B7",
    x"1B802B6",
    x"1B800B5",
    x"1B7FD6C",
    x"1B7F96D",
    x"1B7F56F",
    x"1B7F172",
    x"1B7ED76",
    x"1B7E97B",
    x"1B7E581",
    x"1B7E189",
    x"1B7DD91",
    x"1B7D99A",
    x"1B7D5A4",
    x"1B7D1AF",
    x"1B7CDBB",
    x"1B7C9C8",
    x"1B7C5D6",
    x"1B7C1E5",
    x"1B7BDF5",
    x"1B7BA06",
    x"1B7B618",
    x"1B7B22B",
    x"1B7AE3F",
    x"1B7AA54",
    x"1B7A66A",
    x"1B7A281",
    x"1B79E99",
    x"1B79AB1",
    x"1B796CB",
    x"1B792E6",
    x"1B78F02",
    x"1B78B1F",
    x"1B7873C",
    x"1B7835B",
    x"1B77F7B",
    x"1B77B9B",
    x"1B777BD",
    x"1B773DF",
    x"1B77003",
    x"1B76C27",
    x"1B7684D",
    x"1B76473",
    x"1B7609B",
    x"1B75CC3",
    x"1B758EC",
    x"1B75516",
    x"1B75142",
    x"1B74D6E",
    x"1B7499B",
    x"1B745C9",
    x"1B741F8",
    x"1B73E28",
    x"1B73A59",
    x"1B7368B",
    x"1B732BE",
    x"1B72EF1",
    x"1B72B26",
    x"1B7275C",
    x"1B72393",
    x"1B71FCA",
    x"1B71C03",
    x"1B7183C",
    x"1B71477",
    x"1B710B2",
    x"1B70CEE",
    x"1B7092B",
    x"1B7056A",
    x"1B701A9",
    x"1B6FDE9",
    x"1B6FA2A",
    x"1B6F66C",
    x"1B6F2AF",
    x"1B6EEF2",
    x"1B6EB37",
    x"1B6E77D",
    x"1B6E3C3",
    x"1B6E00B",
    x"1B6DC53",
    x"1B6D89D",
    x"1B6D4E7",
    x"1B6D132",
    x"1B6CD7E",
    x"1B6C9CB",
    x"1B6C619",
    x"1B6C268",
    x"1B6BEB8",
    x"1B6BB09",
    x"1B6B75B",
    x"1B6B3AD",
    x"1B6B001",
    x"1B6AC55",
    x"1B6A8AB",
    x"1B6A501",
    x"1B6A158",
    x"1B69DB0",
    x"1B69A09",
    x"1B69663",
    x"1B692BE",
    x"1B68F1A",
    x"1B68B77",
    x"1B687D4",
    x"1B68433",
    x"1B68092",
    x"1B67CF2",
    x"1B67954",
    x"1B675B6",
    x"1B67219",
    x"1B66E7D",
    x"1B66AE2",
    x"1B66747",
    x"1B663AE",
    x"1B66015",
    x"1B65C7E",
    x"1B658E7",
    x"1B65551",
    x"1B651BD",
    x"1B64E29",
    x"1B64A95",
    x"1B64703",
    x"1B64372",
    x"1B63FE2",
    x"1B63C52",
    x"1B638C3",
    x"1B63536",
    x"1B631A9",
    x"1B62E1D",
    x"1B62A92",
    x"1B62708",
    x"1B6237E",
    x"1B61FF6",
    x"1B61C6E",
    x"1B618E8",
    x"1B61562",
    x"1B611DD",
    x"1B60E59",
    x"1B60AD6",
    x"1B60753",
    x"1B603D2",
    x"1B60051",
    x"1B5FCD2",
    x"1B5F953",
    x"1B5F5D5",
    x"1B5F258",
    x"1B5EEDC",
    x"1B5EB61",
    x"1B5E7E6",
    x"1B5E46D",
    x"1B5E0F4",
    x"1B5DD7C",
    x"1B5DA05",
    x"1B5D68F",
    x"1B5D31A",
    x"1B5CFA6",
    x"1B5CC32",
    x"1B5C8C0",
    x"1B5C54E",
    x"1B5C1DD",
    x"1B5BE6D",
    x"1B5BAFE",
    x"1B5B78F",
    x"1B5B422",
    x"1B5B0B5",
    x"1B5AD4A",
    x"1B5A9DF",
    x"1B5A675",
    x"1B5A30C",
    x"1B59FA3",
    x"1B59C3C",
    x"1B598D5",
    x"1B5956F",
    x"1B5920A",
    x"1B58EA6",
    x"1B58B43",
    x"1B587E1",
    x"1B5847F",
    x"1B5811E",
    x"1B57DBF",
    x"1B57A60",
    x"1B57701",
    x"1B573A4",
    x"1B57048",
    x"1B56CEC",
    x"1B56991",
    x"1B56637",
    x"1B562DE",
    x"1B55F86",
    x"1B55C2E",
    x"1B558D8",
    x"1B55582",
    x"1B5522D",
    x"1B54ED9",
    x"1B54B85",
    x"1B54833",
    x"1B544E1",
    x"1B54190",
    x"1B53E40",
    x"1B53AF1",
    x"1B537A3",
    x"1B53456",
    x"1B53109",
    x"1B52DBD",
    x"1B52A72",
    x"1B52728",
    x"1B523DE",
    x"1B52096",
    x"1B51D4E",
    x"1B51A07",
    x"1B516C1",
    x"1B5137C",
    x"1B51037",
    x"1B50CF4",
    x"1B509B1",
    x"1B5066F",
    x"1B5032E",
    x"1B4FFED",
    x"1B4FCAE",
    x"1B4F96F",
    x"1B4F631",
    x"1B4F2F4",
    x"1B4EFB7",
    x"1B4EC7C",
    x"1B4E941",
    x"1B4E607",
    x"1B4E2CE",
    x"1B4DF96",
    x"1B4DC5E",
    x"1B4D928",
    x"1B4D5F2",
    x"1B4D2BD",
    x"1B4CF88",
    x"1B4CC55",
    x"1B4C922",
    x"1B4C5F0",
    x"1B4C2BF",
    x"1B4BF8F",
    x"1B4BC60",
    x"1B4B931",
    x"1B4B603",
    x"1B4B2D6",
    x"1B4AFAA",
    x"1B4AC7E",
    x"1B4A953",
    x"1B4A629",
    x"1B4A300",
    x"1B49FD8",
    x"1B49CB0",
    x"1B4998A",
    x"1B49664",
    x"1B4933E",
    x"1B4901A",
    x"1B48CF6",
    x"1B489D3",
    x"1B486B1",
    x"1B48390",
    x"1B48070",
    x"1B47D50",
    x"1B47A31",
    x"1B47713",
    x"1B473F5",
    x"1B470D9",
    x"1B46DBD",
    x"1B46AA2",
    x"1B46788",
    x"1B4646E",
    x"1B46155",
    x"1B45E3D",
    x"1B45B26",
    x"1B45810",
    x"1B454FA",
    x"1B451E5",
    x"1B44ED1",
    x"1B44BBE",
    x"1B448AB",
    x"1B4459A",
    x"1B44289",
    x"1B43F78",
    x"1B43C69",
    x"1B4395A",
    x"1B4364C",
    x"1B4333F",
    x"1B43033",
    x"1B42D27",
    x"1B42A1C",
    x"1B42712",
    x"1B42408",
    x"1B42100",
    x"1B41DF8",
    x"1B41AF1",
    x"1B417EB",
    x"1B414E5",
    x"1B411E0",
    x"1B40EDC",
    x"1B40BD9",
    x"1B408D6",
    x"1B405D4",
    x"1B402D3",
    x"1B3FFD3",
    x"1B3FCD3",
    x"1B3F9D4",
    x"1B3F6D6",
    x"1B3F3D9",
    x"1B3F0DC",
    x"1B3EDE1",
    x"1B3EAE5",
    x"1B3E7EB",
    x"1B3E4F1",
    x"1B3E1F9",
    x"1B3DF01",
    x"1B3DC09",
    x"1B3D912",
    x"1B3D61D",
    x"1B3D327",
    x"1B3D033",
    x"1B3CD3F",
    x"1B3CA4C",
    x"1B3C75A",
    x"1B3C469",
    x"1B3C178",
    x"1B3BE88",
    x"1B3BB99",
    x"1B3B8AA",
    x"1B3B5BC",
    x"1B3B2CF",
    x"1B3AFE3",
    x"1B3ACF7",
    x"1B3AA0C",
    x"1B3A722",
    x"1B3A439",
    x"1B3A150",
    x"1B39E68",
    x"1B39B81",
    x"1B3989B",
    x"1B395B5",
    x"1B392D0",
    x"1B38FEB",
    x"1B38D08",
    x"1B38A25",
    x"1B38743",
    x"1B38461",
    x"1B38180",
    x"1B37EA0",
    x"1B37BC1",
    x"1B378E3",
    x"1B37605",
    x"1B37328",
    x"1B3704B",
    x"1B36D6F",
    x"1B36A94",
    x"1B367BA",
    x"1B364E1",
    x"1B36208",
    x"1B35F2F",
    x"1B35C58",
    x"1B35981",
    x"1B356AB",
    x"1B353D6",
    x"1B35101",
    x"1B34E2D",
    x"1B34B5A",
    x"1B34888",
    x"1B345B6",
    x"1B342E5",
    x"1B34015",
    x"1B33D45",
    x"1B33A76",
    x"1B337A8",
    x"1B334DA",
    x"1B3320D",
    x"1B32F41",
    x"1B32C76",
    x"1B329AB",
    x"1B326E1",
    x"1B32417",
    x"1B3214F",
    x"1B31E87",
    x"1B31BBF",
    x"1B318F9",
    x"1B31633",
    x"1B3136E",
    x"1B310A9",
    x"1B30DE5",
    x"1B30B22",
    x"1B30860",
    x"1B3059E",
    x"1B302DD",
    x"1B3001D",
    x"1B2FD5D",
    x"1B2FA9E",
    x"1B2F7E0",
    x"1B2F522",
    x"1B2F265",
    x"1B2EFA9",
    x"1B2ECED",
    x"1B2EA32",
    x"1B2E778",
    x"1B2E4BF",
    x"1B2E206",
    x"1B2DF4E",
    x"1B2DC96",
    x"1B2D9DF",
    x"1B2D729",
    x"1B2D474",
    x"1B2D1BF",
    x"1B2CF0B",
    x"1B2CC57",
    x"1B2C9A5",
    x"1B2C6F3",
    x"1B2C441",
    x"1B2C191",
    x"1B2BEE0",
    x"1B2BC31",
    x"1B2B982",
    x"1B2B6D4",
    x"1B2B427",
    x"1B2B17A",
    x"1B2AECE",
    x"1B2AC23",
    x"1B2A978",
    x"1B2A6CE",
    x"1B2A425",
    x"1B2A17C",
    x"1B29ED4",
    x"1B29C2D",
    x"1B29986",
    x"1B296E0",
    x"1B2943A",
    x"1B29196",
    x"1B28EF2",
    x"1B28C4E",
    x"1B289AC",
    x"1B28709",
    x"1B28468",
    x"1B281C7",
    x"1B27F27",
    x"1B27C88",
    x"1B279E9",
    x"1B2774B",
    x"1B274AD",
    x"1B27210",
    x"1B26F74",
    x"1B26CD9",
    x"1B26A3E",
    x"1B267A4",
    x"1B2650A",
    x"1B26271",
    x"1B25FD9",
    x"1B25D41",
    x"1B25AAA",
    x"1B25814",
    x"1B2557E",
    x"1B252E9",
    x"1B25055",
    x"1B24DC1",
    x"1B24B2E",
    x"1B2489B",
    x"1B24609",
    x"1B24378",
    x"1B240E8",
    x"1B23E58",
    x"1B23BC8",
    x"1B2393A",
    x"1B236AC",
    x"1B2341F",
    x"1B23192",
    x"1B22F06",
    x"1B22C7A",
    x"1B229F0",
    x"1B22765",
    x"1B224DC",
    x"1B22253",
    x"1B21FCB",
    x"1B21D43",
    x"1B21ABC",
    x"1B21836",
    x"1B215B0",
    x"1B2132B",
    x"1B210A6",
    x"1B20E22",
    x"1B20B9F",
    x"1B2091D",
    x"1B2069B",
    x"1B20419",
    x"1B20199",
    x"1B1FF19",
    x"1B1FC99",
    x"1B1FA1A",
    x"1B1F79C",
    x"1B1F51E",
    x"1B1F2A1",
    x"1B1F025",
    x"1B1EDA9",
    x"1B1EB2E",
    x"1B1E8B4",
    x"1B1E63A",
    x"1B1E3C1",
    x"1B1E148",
    x"1B1DED0",
    x"1B1DC59",
    x"1B1D9E2",
    x"1B1D76C",
    x"1B1D4F6",
    x"1B1D281",
    x"1B1D00D",
    x"1B1CD99",
    x"1B1CB26",
    x"1B1C8B4",
    x"1B1C642",
    x"1B1C3D1",
    x"1B1C160",
    x"1B1BEF0",
    x"1B1BC80",
    x"1B1BA12",
    x"1B1B7A3",
    x"1B1B536",
    x"1B1B2C9",
    x"1B1B05C",
    x"1B1ADF1",
    x"1B1AB85",
    x"1B1A91B",
    x"1B1A6B1",
    x"1B1A447",
    x"1B1A1DF",
    x"1B19F77",
    x"1B19D0F",
    x"1B19AA8",
    x"1B19842",
    x"1B195DC",
    x"1B19377",
    x"1B19112",
    x"1B18EAE",
    x"1B18C4B",
    x"1B189E8",
    x"1B18786",
    x"1B18524",
    x"1B182C3",
    x"1B18063",
    x"1B17E03",
    x"1B17BA4",
    x"1B17945",
    x"1B176E7",
    x"1B1748A",
    x"1B1722D",
    x"1B16FD1",
    x"1B16D75",
    x"1B16B1A",
    x"1B168BF",
    x"1B16666",
    x"1B1640C",
    x"1B161B4",
    x"1B15F5B",
    x"1B15D04",
    x"1B15AAD",
    x"1B15857",
    x"1B15601",
    x"1B153AC",
    x"1B15157",
    x"1B14F03",
    x"1B14CAF",
    x"1B14A5D",
    x"1B1480A",
    x"1B145B9",
    x"1B14367",
    x"1B14117",
    x"1B13EC7",
    x"1B13C77",
    x"1B13A29",
    x"1B137DA",
    x"1B1358D",
    x"1B13340",
    x"1B130F3",
    x"1B12EA7",
    x"1B12C5C",
    x"1B12A11",
    x"1B127C7",
    x"1B1257D",
    x"1B12334",
    x"1B120EB",
    x"1B11EA3",
    x"1B11C5C",
    x"1B11A15",
    x"1B117CF",
    x"1B11589",
    x"1B11344",
    x"1B11100",
    x"1B10EBC",
    x"1B10C78",
    x"1B10A36",
    x"1B107F3",
    x"1B105B2",
    x"1B10370",
    x"1B10130",
    x"1B0FEF0",
    x"1B0FCB0",
    x"1B0FA71",
    x"1B0F833",
    x"1B0F5F5",
    x"1B0F3B8",
    x"1B0F17C",
    x"1B0EF3F",
    x"1B0ED04",
    x"1B0EAC9",
    x"1B0E88F",
    x"1B0E655",
    x"1B0E41B",
    x"1B0E1E3",
    x"1B0DFAA",
    x"1B0DD73",
    x"1B0DB3C",
    x"1B0D905",
    x"1B0D6CF",
    x"1B0D49A",
    x"1B0D265",
    x"1B0D031",
    x"1B0CDFD",
    x"1B0CBCA",
    x"1B0C997",
    x"1B0C765",
    x"1B0C533",
    x"1B0C302",
    x"1B0C0D2",
    x"1B0BEA2",
    x"1B0BC72",
    x"1B0BA44",
    x"1B0B815",
    x"1B0B5E7",
    x"1B0B3BA",
    x"1B0B18E",
    x"1B0AF61",
    x"1B0AD36",
    x"1B0AB0B",
    x"1B0A8E0",
    x"1B0A6B6",
    x"1B0A48D",
    x"1B0A264",
    x"1B0A03C",
    x"1B09E14",
    x"1B09BED",
    x"1B099C6",
    x"1B097A0",
    x"1B0957A",
    x"1B09355",
    x"1B09131",
    x"1B08F0D",
    x"1B08CE9",
    x"1B08AC6",
    x"1B088A4",
    x"1B08682",
    x"1B08460",
    x"1B08240",
    x"1B0801F",
    x"1B07E00",
    x"1B07BE0",
    x"1B079C2",
    x"1B077A3",
    x"1B07586",
    x"1B07369",
    x"1B0714C",
    x"1B06F30",
    x"1B06D14",
    x"1B06AF9",
    x"1B068DF",
    x"1B066C5",
    x"1B064AC",
    x"1B06293",
    x"1B0607A",
    x"1B05E62",
    x"1B05C4B",
    x"1B05A34",
    x"1B0581E",
    x"1B05608",
    x"1B053F3",
    x"1B051DE",
    x"1B04FCA",
    x"1B04DB6",
    x"1B04BA3",
    x"1B04991",
    x"1B0477E",
    x"1B0456D",
    x"1B0435C",
    x"1B0414B",
    x"1B03F3B",
    x"1B03D2C",
    x"1B03B1C",
    x"1B0390E",
    x"1B03700",
    x"1B034F2",
    x"1B032E5",
    x"1B030D9",
    x"1B02ECD",
    x"1B02CC2",
    x"1B02AB7",
    x"1B028AC",
    x"1B026A2",
    x"1B02499",
    x"1B02290",
    x"1B02088",
    x"1B01E80",
    x"1B01C78",
    x"1B01A72",
    x"1B0186B",
    x"1B01665",
    x"1B01460",
    x"1B0125B",
    x"1B01057",
    x"1B00E53",
    x"1B00C50",
    x"1B00A4D",
    x"1B0084A",
    x"1B00649",
    x"1B00447",
    x"1B00247",
    x"1B00046",
    x"1AFFC8D",
    x"1AFF88F",
    x"1AFF491",
    x"1AFF094",
    x"1AFEC99",
    x"1AFE89E",
    x"1AFE4A4",
    x"1AFE0AC",
    x"1AFDCB4",
    x"1AFD8BD",
    x"1AFD4C8",
    x"1AFD0D3",
    x"1AFCCDF",
    x"1AFC8ED",
    x"1AFC4FB",
    x"1AFC10A",
    x"1AFBD1A",
    x"1AFB92B",
    x"1AFB53E",
    x"1AFB151",
    x"1AFAD65",
    x"1AFA97A",
    x"1AFA590",
    x"1AFA1A7",
    x"1AF9DBF",
    x"1AF99D9",
    x"1AF95F3",
    x"1AF920E",
    x"1AF8E2A",
    x"1AF8A46",
    x"1AF8664",
    x"1AF8283",
    x"1AF7EA3",
    x"1AF7AC4",
    x"1AF76E6",
    x"1AF7308",
    x"1AF6F2C",
    x"1AF6B51",
    x"1AF6777",
    x"1AF639D",
    x"1AF5FC5",
    x"1AF5BED",
    x"1AF5817",
    x"1AF5441",
    x"1AF506D",
    x"1AF4C99",
    x"1AF48C6",
    x"1AF44F5",
    x"1AF4124",
    x"1AF3D54",
    x"1AF3985",
    x"1AF35B7",
    x"1AF31EA",
    x"1AF2E1E",
    x"1AF2A53",
    x"1AF2689",
    x"1AF22C0",
    x"1AF1EF8",
    x"1AF1B31",
    x"1AF176A",
    x"1AF13A5",
    x"1AF0FE0",
    x"1AF0C1D",
    x"1AF085A",
    x"1AF0499",
    x"1AF00D8",
    x"1AEFD18",
    x"1AEF959",
    x"1AEF59C",
    x"1AEF1DF",
    x"1AEEE23",
    x"1AEEA68",
    x"1AEE6AD",
    x"1AEE2F4",
    x"1AEDF3C",
    x"1AEDB85",
    x"1AED7CE",
    x"1AED419",
    x"1AED064",
    x"1AECCB1",
    x"1AEC8FE",
    x"1AEC54C",
    x"1AEC19B",
    x"1AEBDEB",
    x"1AEBA3C",
    x"1AEB68E",
    x"1AEB2E1",
    x"1AEAF35",
    x"1AEAB89",
    x"1AEA7DF",
    x"1AEA435",
    x"1AEA08D",
    x"1AE9CE5",
    x"1AE993E",
    x"1AE9599",
    x"1AE91F4",
    x"1AE8E50",
    x"1AE8AAC",
    x"1AE870A",
    x"1AE8369",
    x"1AE7FC8",
    x"1AE7C29",
    x"1AE788A",
    x"1AE74ED",
    x"1AE7150",
    x"1AE6DB4",
    x"1AE6A19",
    x"1AE667F",
    x"1AE62E6",
    x"1AE5F4E",
    x"1AE5BB6",
    x"1AE5820",
    x"1AE548A",
    x"1AE50F5",
    x"1AE4D62",
    x"1AE49CF",
    x"1AE463D",
    x"1AE42AC",
    x"1AE3F1B",
    x"1AE3B8C",
    x"1AE37FE",
    x"1AE3470",
    x"1AE30E3",
    x"1AE2D58",
    x"1AE29CD",
    x"1AE2643",
    x"1AE22BA",
    x"1AE1F31",
    x"1AE1BAA",
    x"1AE1824",
    x"1AE149E",
    x"1AE1119",
    x"1AE0D95",
    x"1AE0A12",
    x"1AE0690",
    x"1AE030F",
    x"1ADFF8F",
    x"1ADFC0F",
    x"1ADF891",
    x"1ADF513",
    x"1ADF196",
    x"1ADEE1A",
    x"1ADEA9F",
    x"1ADE725",
    x"1ADE3AC",
    x"1ADE033",
    x"1ADDCBC",
    x"1ADD945",
    x"1ADD5CF",
    x"1ADD25A",
    x"1ADCEE6",
    x"1ADCB72",
    x"1ADC800",
    x"1ADC48E",
    x"1ADC11E",
    x"1ADBDAE",
    x"1ADBA3F",
    x"1ADB6D1",
    x"1ADB363",
    x"1ADAFF7",
    x"1ADAC8B",
    x"1ADA921",
    x"1ADA5B7",
    x"1ADA24E",
    x"1AD9EE6",
    x"1AD9B7E",
    x"1AD9818",
    x"1AD94B2",
    x"1AD914E",
    x"1AD8DEA",
    x"1AD8A87",
    x"1AD8724",
    x"1AD83C3",
    x"1AD8063",
    x"1AD7D03",
    x"1AD79A4",
    x"1AD7646",
    x"1AD72E9",
    x"1AD6F8D",
    x"1AD6C31",
    x"1AD68D7",
    x"1AD657D",
    x"1AD6224",
    x"1AD5ECC",
    x"1AD5B74",
    x"1AD581E",
    x"1AD54C8",
    x"1AD5174",
    x"1AD4E20",
    x"1AD4ACD",
    x"1AD477A",
    x"1AD4429",
    x"1AD40D8",
    x"1AD3D88",
    x"1AD3A39",
    x"1AD36EB",
    x"1AD339E",
    x"1AD3051",
    x"1AD2D06",
    x"1AD29BB",
    x"1AD2671",
    x"1AD2328",
    x"1AD1FDF",
    x"1AD1C98",
    x"1AD1951",
    x"1AD160B",
    x"1AD12C6",
    x"1AD0F82",
    x"1AD0C3E",
    x"1AD08FC",
    x"1AD05BA",
    x"1AD0279",
    x"1ACFF38",
    x"1ACFBF9",
    x"1ACF8BB",
    x"1ACF57D",
    x"1ACF240",
    x"1ACEF04",
    x"1ACEBC8",
    x"1ACE88E",
    x"1ACE554",
    x"1ACE21B",
    x"1ACDEE3",
    x"1ACDBAC",
    x"1ACD875",
    x"1ACD53F",
    x"1ACD20A",
    x"1ACCED6",
    x"1ACCBA3",
    x"1ACC871",
    x"1ACC53F",
    x"1ACC20E",
    x"1ACBEDE",
    x"1ACBBAE",
    x"1ACB880",
    x"1ACB552",
    x"1ACB225",
    x"1ACAEF9",
    x"1ACABCE",
    x"1ACA8A3",
    x"1ACA579",
    x"1ACA251",
    x"1AC9F28",
    x"1AC9C01",
    x"1AC98DA",
    x"1AC95B5",
    x"1AC928F",
    x"1AC8F6B",
    x"1AC8C48",
    x"1AC8925",
    x"1AC8603",
    x"1AC82E2",
    x"1AC7FC2",
    x"1AC7CA2",
    x"1AC7983",
    x"1AC7665",
    x"1AC7348",
    x"1AC702C",
    x"1AC6D10",
    x"1AC69F5",
    x"1AC66DB",
    x"1AC63C2",
    x"1AC60A9",
    x"1AC5D91",
    x"1AC5A7A",
    x"1AC5764",
    x"1AC544F",
    x"1AC513A",
    x"1AC4E26",
    x"1AC4B13",
    x"1AC4801",
    x"1AC44EF",
    x"1AC41DE",
    x"1AC3ECE",
    x"1AC3BBF",
    x"1AC38B0",
    x"1AC35A2",
    x"1AC3295",
    x"1AC2F89",
    x"1AC2C7E",
    x"1AC2973",
    x"1AC2669",
    x"1AC2360",
    x"1AC2057",
    x"1AC1D50",
    x"1AC1A49",
    x"1AC1742",
    x"1AC143D",
    x"1AC1138",
    x"1AC0E34",
    x"1AC0B31",
    x"1AC082F",
    x"1AC052D",
    x"1AC022C",
    x"1ABFF2C",
    x"1ABFC2D",
    x"1ABF92E",
    x"1ABF630",
    x"1ABF333",
    x"1ABF036",
    x"1ABED3B",
    x"1ABEA40",
    x"1ABE746",
    x"1ABE44C",
    x"1ABE153",
    x"1ABDE5B",
    x"1ABDB64",
    x"1ABD86E",
    x"1ABD578",
    x"1ABD283",
    x"1ABCF8F",
    x"1ABCC9B",
    x"1ABC9A8",
    x"1ABC6B6",
    x"1ABC3C5",
    x"1ABC0D5",
    x"1ABBDE5",
    x"1ABBAF6",
    x"1ABB807",
    x"1ABB51A",
    x"1ABB22D",
    x"1ABAF40",
    x"1ABAC55",
    x"1ABA96A",
    x"1ABA680",
    x"1ABA397",
    x"1ABA0AF",
    x"1AB9DC7",
    x"1AB9AE0",
    x"1AB97F9",
    x"1AB9514",
    x"1AB922F",
    x"1AB8F4B",
    x"1AB8C67",
    x"1AB8984",
    x"1AB86A2",
    x"1AB83C1",
    x"1AB80E0",
    x"1AB7E01",
    x"1AB7B21",
    x"1AB7843",
    x"1AB7565",
    x"1AB7288",
    x"1AB6FAC",
    x"1AB6CD0",
    x"1AB69F6",
    x"1AB671B",
    x"1AB6442",
    x"1AB6169",
    x"1AB5E91",
    x"1AB5BBA",
    x"1AB58E3",
    x"1AB560E",
    x"1AB5338",
    x"1AB5064",
    x"1AB4D90",
    x"1AB4ABD",
    x"1AB47EB",
    x"1AB4519",
    x"1AB4248",
    x"1AB3F78",
    x"1AB3CA9",
    x"1AB39DA",
    x"1AB370C",
    x"1AB343E",
    x"1AB3172",
    x"1AB2EA6",
    x"1AB2BDA",
    x"1AB2910",
    x"1AB2646",
    x"1AB237C",
    x"1AB20B4",
    x"1AB1DEC",
    x"1AB1B25",
    x"1AB185F",
    x"1AB1599",
    x"1AB12D4",
    x"1AB100F",
    x"1AB0D4C",
    x"1AB0A89",
    x"1AB07C6",
    x"1AB0505",
    x"1AB0244",
    x"1AAFF84",
    x"1AAFCC4",
    x"1AAFA05",
    x"1AAF747",
    x"1AAF48A",
    x"1AAF1CD",
    x"1AAEF11",
    x"1AAEC55",
    x"1AAE99B",
    x"1AAE6E1",
    x"1AAE427",
    x"1AAE16E",
    x"1AADEB6",
    x"1AADBFF",
    x"1AAD948",
    x"1AAD692",
    x"1AAD3DD",
    x"1AAD129",
    x"1AACE75",
    x"1AACBC1",
    x"1AAC90F",
    x"1AAC65D",
    x"1AAC3AC",
    x"1AAC0FB",
    x"1AABE4B",
    x"1AABB9C",
    x"1AAB8ED",
    x"1AAB63F",
    x"1AAB392",
    x"1AAB0E6",
    x"1AAAE3A",
    x"1AAAB8E",
    x"1AAA8E4",
    x"1AAA63A",
    x"1AAA391",
    x"1AAA0E8",
    x"1AA9E40",
    x"1AA9B99",
    x"1AA98F3",
    x"1AA964D",
    x"1AA93A7",
    x"1AA9103",
    x"1AA8E5F",
    x"1AA8BBC",
    x"1AA8919",
    x"1AA8677",
    x"1AA83D6",
    x"1AA8135",
    x"1AA7E95",
    x"1AA7BF6",
    x"1AA7957",
    x"1AA76B9",
    x"1AA741C",
    x"1AA717F",
    x"1AA6EE3",
    x"1AA6C48",
    x"1AA69AD",
    x"1AA6713",
    x"1AA6479",
    x"1AA61E1",
    x"1AA5F48",
    x"1AA5CB1",
    x"1AA5A1A",
    x"1AA5784",
    x"1AA54EE",
    x"1AA5259",
    x"1AA4FC5",
    x"1AA4D32",
    x"1AA4A9F",
    x"1AA480C",
    x"1AA457B",
    x"1AA42EA",
    x"1AA4059",
    x"1AA3DC9",
    x"1AA3B3A",
    x"1AA38AC",
    x"1AA361E",
    x"1AA3391",
    x"1AA3104",
    x"1AA2E78",
    x"1AA2BED",
    x"1AA2962",
    x"1AA26D8",
    x"1AA244F",
    x"1AA21C6",
    x"1AA1F3E",
    x"1AA1CB6",
    x"1AA1A30",
    x"1AA17A9",
    x"1AA1524",
    x"1AA129F",
    x"1AA101A",
    x"1AA0D97",
    x"1AA0B14",
    x"1AA0891",
    x"1AA060F",
    x"1AA038E",
    x"1AA010E",
    x"1A9FE8E",
    x"1A9FC0E",
    x"1A9F990",
    x"1A9F711",
    x"1A9F494",
    x"1A9F217",
    x"1A9EF9B",
    x"1A9ED1F",
    x"1A9EAA4",
    x"1A9E82A",
    x"1A9E5B0",
    x"1A9E337",
    x"1A9E0BF",
    x"1A9DE47",
    x"1A9DBD0",
    x"1A9D959",
    x"1A9D6E3",
    x"1A9D46D",
    x"1A9D1F9",
    x"1A9CF84",
    x"1A9CD11",
    x"1A9CA9E",
    x"1A9C82C",
    x"1A9C5BA",
    x"1A9C349",
    x"1A9C0D8",
    x"1A9BE68",
    x"1A9BBF9",
    x"1A9B98A",
    x"1A9B71C",
    x"1A9B4AF",
    x"1A9B242",
    x"1A9AFD6",
    x"1A9AD6A",
    x"1A9AAFF",
    x"1A9A894",
    x"1A9A62B",
    x"1A9A3C1",
    x"1A9A159",
    x"1A99EF1",
    x"1A99C89",
    x"1A99A22",
    x"1A997BC",
    x"1A99557",
    x"1A992F2",
    x"1A9908D",
    x"1A98E29",
    x"1A98BC6",
    x"1A98963",
    x"1A98701",
    x"1A984A0",
    x"1A9823F",
    x"1A97FDF",
    x"1A97D7F",
    x"1A97B20",
    x"1A978C2",
    x"1A97664",
    x"1A97406",
    x"1A971AA",
    x"1A96F4D",
    x"1A96CF2",
    x"1A96A97",
    x"1A9683D",
    x"1A965E3",
    x"1A9638A",
    x"1A96131",
    x"1A95ED9",
    x"1A95C82",
    x"1A95A2B",
    x"1A957D5",
    x"1A9557F",
    x"1A9532A",
    x"1A950D5",
    x"1A94E81",
    x"1A94C2E",
    x"1A949DB",
    x"1A94789",
    x"1A94538",
    x"1A942E7",
    x"1A94096",
    x"1A93E46",
    x"1A93BF7",
    x"1A939A8",
    x"1A9375A",
    x"1A9350D",
    x"1A932C0",
    x"1A93073",
    x"1A92E27",
    x"1A92BDC",
    x"1A92991",
    x"1A92747",
    x"1A924FE",
    x"1A922B5",
    x"1A9206C",
    x"1A91E25",
    x"1A91BDD",
    x"1A91997",
    x"1A91751",
    x"1A9150B",
    x"1A912C6",
    x"1A91082",
    x"1A90E3E",
    x"1A90BFB",
    x"1A909B8",
    x"1A90776",
    x"1A90534",
    x"1A902F3",
    x"1A900B3",
    x"1A8FE73",
    x"1A8FC33",
    x"1A8F9F5",
    x"1A8F7B6",
    x"1A8F579",
    x"1A8F33C",
    x"1A8F0FF",
    x"1A8EEC3",
    x"1A8EC88",
    x"1A8EA4D",
    x"1A8E813",
    x"1A8E5D9",
    x"1A8E3A0",
    x"1A8E167",
    x"1A8DF2F",
    x"1A8DCF8",
    x"1A8DAC1",
    x"1A8D88A",
    x"1A8D654",
    x"1A8D41F",
    x"1A8D1EA",
    x"1A8CFB6",
    x"1A8CD82",
    x"1A8CB4F",
    x"1A8C91D",
    x"1A8C6EB",
    x"1A8C4B9",
    x"1A8C288",
    x"1A8C058",
    x"1A8BE28",
    x"1A8BBF9",
    x"1A8B9CA",
    x"1A8B79C",
    x"1A8B56E",
    x"1A8B341",
    x"1A8B115",
    x"1A8AEE9",
    x"1A8ACBD",
    x"1A8AA92",
    x"1A8A868",
    x"1A8A63E",
    x"1A8A415",
    x"1A8A1EC",
    x"1A89FC4",
    x"1A89D9C",
    x"1A89B75",
    x"1A8994F",
    x"1A89728",
    x"1A89503",
    x"1A892DE",
    x"1A890B9",
    x"1A88E96",
    x"1A88C72",
    x"1A88A4F",
    x"1A8882D",
    x"1A8860B",
    x"1A883EA",
    x"1A881C9",
    x"1A87FA9",
    x"1A87D89",
    x"1A87B6A",
    x"1A8794C",
    x"1A8772E",
    x"1A87510",
    x"1A872F3",
    x"1A870D7",
    x"1A86EBB",
    x"1A86C9F",
    x"1A86A84",
    x"1A8686A",
    x"1A86650",
    x"1A86437",
    x"1A8621E",
    x"1A86006",
    x"1A85DEE",
    x"1A85BD7",
    x"1A859C0",
    x"1A857AA",
    x"1A85594",
    x"1A8537F",
    x"1A8516B",
    x"1A84F57",
    x"1A84D43",
    x"1A84B30",
    x"1A8491D",
    x"1A8470B",
    x"1A844FA",
    x"1A842E9",
    x"1A840D8",
    x"1A83EC8",
    x"1A83CB9",
    x"1A83AAA",
    x"1A8389C",
    x"1A8368E",
    x"1A83480",
    x"1A83273",
    x"1A83067",
    x"1A82E5B",
    x"1A82C50",
    x"1A82A45",
    x"1A8283B",
    x"1A82631",
    x"1A82428",
    x"1A8221F",
    x"1A82017",
    x"1A81E0F",
    x"1A81C08",
    x"1A81A01",
    x"1A817FB",
    x"1A815F5",
    x"1A813F0",
    x"1A811EB",
    x"1A80FE7",
    x"1A80DE3",
    x"1A80BE0",
    x"1A809DD",
    x"1A807DB",
    x"1A805D9",
    x"1A803D8",
    x"1A801D7",
    x"1A7FFAE",
    x"1A7FBAF",
    x"1A7F7B1",
    x"1A7F3B3",
    x"1A7EFB7",
    x"1A7EBBB",
    x"1A7E7C1",
    x"1A7E3C7",
    x"1A7DFCF",
    x"1A7DBD7",
    x"1A7D7E1",
    x"1A7D3EC",
    x"1A7CFF7",
    x"1A7CC04",
    x"1A7C811",
    x"1A7C420",
    x"1A7C02F",
    x"1A7BC3F",
    x"1A7B851",
    x"1A7B463",
    x"1A7B077",
    x"1A7AC8B",
    x"1A7A8A0",
    x"1A7A4B7",
    x"1A7A0CE",
    x"1A79CE6",
    x"1A79900",
    x"1A7951A",
    x"1A79135",
    x"1A78D51",
    x"1A7896E",
    x"1A7858C",
    x"1A781AC",
    x"1A77DCC",
    x"1A779ED",
    x"1A7760F",
    x"1A77232",
    x"1A76E56",
    x"1A76A7A",
    x"1A766A0",
    x"1A762C7",
    x"1A75EEF",
    x"1A75B18",
    x"1A75741",
    x"1A7536C",
    x"1A74F98",
    x"1A74BC4",
    x"1A747F2",
    x"1A74420",
    x"1A74050",
    x"1A73C80",
    x"1A738B2",
    x"1A734E4",
    x"1A73117",
    x"1A72D4B",
    x"1A72980",
    x"1A725B7",
    x"1A721EE",
    x"1A71E26",
    x"1A71A5E",
    x"1A71698",
    x"1A712D3",
    x"1A70F0F",
    x"1A70B4C",
    x"1A70789",
    x"1A703C8",
    x"1A70007",
    x"1A6FC48",
    x"1A6F889",
    x"1A6F4CC",
    x"1A6F10F",
    x"1A6ED53",
    x"1A6E998",
    x"1A6E5DE",
    x"1A6E225",
    x"1A6DE6D",
    x"1A6DAB6",
    x"1A6D700",
    x"1A6D34B",
    x"1A6CF96",
    x"1A6CBE3",
    x"1A6C830",
    x"1A6C47F",
    x"1A6C0CE",
    x"1A6BD1E",
    x"1A6B96F",
    x"1A6B5C2",
    x"1A6B215",
    x"1A6AE68",
    x"1A6AABD",
    x"1A6A713",
    x"1A6A36A",
    x"1A69FC1",
    x"1A69C1A",
    x"1A69873",
    x"1A694CE",
    x"1A69129",
    x"1A68D85",
    x"1A689E2",
    x"1A68640",
    x"1A6829F",
    x"1A67EFF",
    x"1A67B60",
    x"1A677C1",
    x"1A67424",
    x"1A67087",
    x"1A66CEB",
    x"1A66951",
    x"1A665B7",
    x"1A6621E",
    x"1A65E86",
    x"1A65AEF",
    x"1A65758",
    x"1A653C3",
    x"1A6502E",
    x"1A64C9B",
    x"1A64908",
    x"1A64576",
    x"1A641E5",
    x"1A63E55",
    x"1A63AC6",
    x"1A63738",
    x"1A633AB",
    x"1A6301E",
    x"1A62C92",
    x"1A62908",
    x"1A6257E",
    x"1A621F5",
    x"1A61E6D",
    x"1A61AE6",
    x"1A61760",
    x"1A613DA",
    x"1A61056",
    x"1A60CD2",
    x"1A6094F",
    x"1A605CD",
    x"1A6024C",
    x"1A5FECC",
    x"1A5FB4D",
    x"1A5F7CF",
    x"1A5F451",
    x"1A5F0D4",
    x"1A5ED59",
    x"1A5E9DE",
    x"1A5E664",
    x"1A5E2EA",
    x"1A5DF72",
    x"1A5DBFB",
    x"1A5D884",
    x"1A5D50F",
    x"1A5D19A",
    x"1A5CE26",
    x"1A5CAB3",
    x"1A5C740",
    x"1A5C3CF",
    x"1A5C05E",
    x"1A5BCEF",
    x"1A5B980",
    x"1A5B612",
    x"1A5B2A5",
    x"1A5AF39",
    x"1A5ABCD",
    x"1A5A863",
    x"1A5A4F9",
    x"1A5A190",
    x"1A59E28",
    x"1A59AC1",
    x"1A5975B",
    x"1A593F6",
    x"1A59091",
    x"1A58D2D",
    x"1A589CA",
    x"1A58668",
    x"1A58307",
    x"1A57FA7",
    x"1A57C47",
    x"1A578E9",
    x"1A5758B",
    x"1A5722E",
    x"1A56ED2",
    x"1A56B77",
    x"1A5681C",
    x"1A564C2",
    x"1A5616A",
    x"1A55E12",
    x"1A55ABB",
    x"1A55764",
    x"1A5540F",
    x"1A550BA",
    x"1A54D67",
    x"1A54A14",
    x"1A546C2",
    x"1A54370",
    x"1A54020",
    x"1A53CD0",
    x"1A53981",
    x"1A53633",
    x"1A532E6",
    x"1A52F9A",
    x"1A52C4F",
    x"1A52904",
    x"1A525BA",
    x"1A52271",
    x"1A51F29",
    x"1A51BE1",
    x"1A5189B",
    x"1A51555",
    x"1A51210",
    x"1A50ECC",
    x"1A50B89",
    x"1A50846",
    x"1A50505",
    x"1A501C4",
    x"1A4FE84",
    x"1A4FB45",
    x"1A4F806",
    x"1A4F4C9",
    x"1A4F18C",
    x"1A4EE50",
    x"1A4EB15",
    x"1A4E7DA",
    x"1A4E4A1",
    x"1A4E168",
    x"1A4DE30",
    x"1A4DAF9",
    x"1A4D7C2",
    x"1A4D48D",
    x"1A4D158",
    x"1A4CE24",
    x"1A4CAF1",
    x"1A4C7BF",
    x"1A4C48D",
    x"1A4C15D",
    x"1A4BE2D",
    x"1A4BAFD",
    x"1A4B7CF",
    x"1A4B4A2",
    x"1A4B175",
    x"1A4AE49",
    x"1A4AB1E",
    x"1A4A7F3",
    x"1A4A4CA",
    x"1A4A1A1",
    x"1A49E79",
    x"1A49B52",
    x"1A4982B",
    x"1A49506",
    x"1A491E1",
    x"1A48EBD",
    x"1A48B99",
    x"1A48877",
    x"1A48555",
    x"1A48234",
    x"1A47F14",
    x"1A47BF5",
    x"1A478D6",
    x"1A475B8",
    x"1A4729B",
    x"1A46F7F",
    x"1A46C63",
    x"1A46949",
    x"1A4662F",
    x"1A46316",
    x"1A45FFD",
    x"1A45CE6",
    x"1A459CF",
    x"1A456B9",
    x"1A453A3",
    x"1A4508F",
    x"1A44D7B",
    x"1A44A68",
    x"1A44756",
    x"1A44444",
    x"1A44134",
    x"1A43E24",
    x"1A43B15",
    x"1A43806",
    x"1A434F9",
    x"1A431EC",
    x"1A42EE0",
    x"1A42BD4",
    x"1A428CA",
    x"1A425C0",
    x"1A422B7",
    x"1A41FAF",
    x"1A41CA7",
    x"1A419A0",
    x"1A4169A",
    x"1A41395",
    x"1A41090",
    x"1A40D8D",
    x"1A40A8A",
    x"1A40787",
    x"1A40486",
    x"1A40185",
    x"1A3FE85",
    x"1A3FB86",
    x"1A3F887",
    x"1A3F58A",
    x"1A3F28D",
    x"1A3EF90",
    x"1A3EC95",
    x"1A3E99A",
    x"1A3E6A0",
    x"1A3E3A7",
    x"1A3E0AE",
    x"1A3DDB6",
    x"1A3DABF",
    x"1A3D7C9",
    x"1A3D4D3",
    x"1A3D1DF",
    x"1A3CEEB",
    x"1A3CBF7",
    x"1A3C905",
    x"1A3C613",
    x"1A3C321",
    x"1A3C031",
    x"1A3BD41",
    x"1A3BA52",
    x"1A3B764",
    x"1A3B477",
    x"1A3B18A",
    x"1A3AE9E",
    x"1A3ABB3",
    x"1A3A8C8",
    x"1A3A5DE",
    x"1A3A2F5",
    x"1A3A00D",
    x"1A39D25",
    x"1A39A3E",
    x"1A39758",
    x"1A39473",
    x"1A3918E",
    x"1A38EAA",
    x"1A38BC6",
    x"1A388E4",
    x"1A38602",
    x"1A38321",
    x"1A38040",
    x"1A37D61",
    x"1A37A82",
    x"1A377A4",
    x"1A374C6",
    x"1A371E9",
    x"1A36F0D",
    x"1A36C32",
    x"1A36957",
    x"1A3667D",
    x"1A363A4",
    x"1A360CB",
    x"1A35DF3",
    x"1A35B1C",
    x"1A35846",
    x"1A35570",
    x"1A3529B",
    x"1A34FC7",
    x"1A34CF3",
    x"1A34A20",
    x"1A3474E",
    x"1A3447D",
    x"1A341AC",
    x"1A33EDC",
    x"1A33C0C",
    x"1A3393E",
    x"1A33670",
    x"1A333A2",
    x"1A330D6",
    x"1A32E0A",
    x"1A32B3F",
    x"1A32874",
    x"1A325AB",
    x"1A322E2",
    x"1A32019",
    x"1A31D52",
    x"1A31A8B",
    x"1A317C4",
    x"1A314FF",
    x"1A3123A",
    x"1A30F76",
    x"1A30CB2",
    x"1A309EF",
    x"1A3072D",
    x"1A3046C",
    x"1A301AB",
    x"1A2FEEB",
    x"1A2FC2B",
    x"1A2F96D",
    x"1A2F6AF",
    x"1A2F3F1",
    x"1A2F135",
    x"1A2EE79",
    x"1A2EBBD",
    x"1A2E903",
    x"1A2E649",
    x"1A2E390",
    x"1A2E0D7",
    x"1A2DE1F",
    x"1A2DB68",
    x"1A2D8B2",
    x"1A2D5FC",
    x"1A2D347",
    x"1A2D092",
    x"1A2CDDE",
    x"1A2CB2B",
    x"1A2C879",
    x"1A2C5C7",
    x"1A2C316",
    x"1A2C065",
    x"1A2BDB6",
    x"1A2BB07",
    x"1A2B858",
    x"1A2B5AA",
    x"1A2B2FD",
    x"1A2B051",
    x"1A2ADA5",
    x"1A2AAFA",
    x"1A2A850",
    x"1A2A5A6",
    x"1A2A2FD",
    x"1A2A054",
    x"1A29DAD",
    x"1A29B06",
    x"1A2985F",
    x"1A295B9",
    x"1A29314",
    x"1A29070",
    x"1A28DCC",
    x"1A28B29",
    x"1A28887",
    x"1A285E5",
    x"1A28344",
    x"1A280A3",
    x"1A27E03",
    x"1A27B64",
    x"1A278C6",
    x"1A27628",
    x"1A2738A",
    x"1A270EE",
    x"1A26E52",
    x"1A26BB7",
    x"1A2691C",
    x"1A26682",
    x"1A263E9",
    x"1A26150",
    x"1A25EB8",
    x"1A25C21",
    x"1A2598A",
    x"1A256F4",
    x"1A2545F",
    x"1A251CA",
    x"1A24F36",
    x"1A24CA2",
    x"1A24A0F",
    x"1A2477D",
    x"1A244EC",
    x"1A2425B",
    x"1A23FCB",
    x"1A23D3B",
    x"1A23AAC",
    x"1A2381E",
    x"1A23590",
    x"1A23303",
    x"1A23076",
    x"1A22DEB",
    x"1A22B5F",
    x"1A228D5",
    x"1A2264B",
    x"1A223C2",
    x"1A22139",
    x"1A21EB1",
    x"1A21C2A",
    x"1A219A3",
    x"1A2171D",
    x"1A21497",
    x"1A21213",
    x"1A20F8E",
    x"1A20D0B",
    x"1A20A88",
    x"1A20806",
    x"1A20584",
    x"1A20303",
    x"1A20082",
    x"1A1FE03",
    x"1A1FB83",
    x"1A1F905",
    x"1A1F687",
    x"1A1F40A",
    x"1A1F18D",
    x"1A1EF11",
    x"1A1EC95",
    x"1A1EA1A",
    x"1A1E7A0",
    x"1A1E527",
    x"1A1E2AE",
    x"1A1E035",
    x"1A1DDBE",
    x"1A1DB46",
    x"1A1D8D0",
    x"1A1D65A",
    x"1A1D3E5",
    x"1A1D170",
    x"1A1CEFC",
    x"1A1CC89",
    x"1A1CA16",
    x"1A1C7A4",
    x"1A1C532",
    x"1A1C2C1",
    x"1A1C051",
    x"1A1BDE1",
    x"1A1BB72",
    x"1A1B903",
    x"1A1B695",
    x"1A1B428",
    x"1A1B1BB",
    x"1A1AF4F",
    x"1A1ACE3",
    x"1A1AA78",
    x"1A1A80E",
    x"1A1A5A4",
    x"1A1A33B",
    x"1A1A0D3",
    x"1A19E6B",
    x"1A19C04",
    x"1A1999D",
    x"1A19737",
    x"1A194D1",
    x"1A1926C",
    x"1A19008",
    x"1A18DA4",
    x"1A18B41",
    x"1A188DF",
    x"1A1867D",
    x"1A1841C",
    x"1A181BB",
    x"1A17F5B",
    x"1A17CFB",
    x"1A17A9C",
    x"1A1783E",
    x"1A175E0",
    x"1A17383",
    x"1A17126",
    x"1A16ECA",
    x"1A16C6F",
    x"1A16A14",
    x"1A167BA",
    x"1A16560",
    x"1A16307",
    x"1A160AF",
    x"1A15E57",
    x"1A15C00",
    x"1A159A9",
    x"1A15753",
    x"1A154FD",
    x"1A152A8",
    x"1A15054",
    x"1A14E00",
    x"1A14BAD",
    x"1A1495A",
    x"1A14708",
    x"1A144B7",
    x"1A14266",
    x"1A14015",
    x"1A13DC6",
    x"1A13B77",
    x"1A13928",
    x"1A136DA",
    x"1A1348D",
    x"1A13240",
    x"1A12FF3",
    x"1A12DA8",
    x"1A12B5D",
    x"1A12912",
    x"1A126C8",
    x"1A1247F",
    x"1A12236",
    x"1A11FEE",
    x"1A11DA6",
    x"1A11B5F",
    x"1A11918",
    x"1A116D2",
    x"1A1148D",
    x"1A11248",
    x"1A11004",
    x"1A10DC0",
    x"1A10B7D",
    x"1A1093A",
    x"1A106F8",
    x"1A104B7",
    x"1A10276",
    x"1A10035",
    x"1A0FDF6",
    x"1A0FBB6",
    x"1A0F978",
    x"1A0F73A",
    x"1A0F4FC",
    x"1A0F2BF",
    x"1A0F083",
    x"1A0EE47",
    x"1A0EC0C",
    x"1A0E9D1",
    x"1A0E797",
    x"1A0E55D",
    x"1A0E324",
    x"1A0E0EC",
    x"1A0DEB4",
    x"1A0DC7C",
    x"1A0DA45",
    x"1A0D80F",
    x"1A0D5D9",
    x"1A0D3A4",
    x"1A0D170",
    x"1A0CF3B",
    x"1A0CD08",
    x"1A0CAD5",
    x"1A0C8A3",
    x"1A0C671",
    x"1A0C43F",
    x"1A0C20F",
    x"1A0BFDE",
    x"1A0BDAF",
    x"1A0BB7F",
    x"1A0B951",
    x"1A0B723",
    x"1A0B4F5",
    x"1A0B2C8",
    x"1A0B09C",
    x"1A0AE70",
    x"1A0AC45",
    x"1A0AA1A",
    x"1A0A7F0",
    x"1A0A5C6",
    x"1A0A39D",
    x"1A0A174",
    x"1A09F4C",
    x"1A09D24",
    x"1A09AFD",
    x"1A098D7",
    x"1A096B1",
    x"1A0948C",
    x"1A09267",
    x"1A09042",
    x"1A08E1F",
    x"1A08BFB",
    x"1A089D9",
    x"1A087B6",
    x"1A08595",
    x"1A08374",
    x"1A08153",
    x"1A07F33",
    x"1A07D13",
    x"1A07AF4",
    x"1A078D6",
    x"1A076B8",
    x"1A0749B",
    x"1A0727E",
    x"1A07061",
    x"1A06E45",
    x"1A06C2A",
    x"1A06A0F",
    x"1A067F5",
    x"1A065DB",
    x"1A063C2",
    x"1A061AA",
    x"1A05F91",
    x"1A05D7A",
    x"1A05B63",
    x"1A0594C",
    x"1A05736",
    x"1A05520",
    x"1A0530B",
    x"1A050F7",
    x"1A04EE3",
    x"1A04CCF",
    x"1A04ABD",
    x"1A048AA",
    x"1A04698",
    x"1A04487",
    x"1A04276",
    x"1A04066",
    x"1A03E56",
    x"1A03C46",
    x"1A03A38",
    x"1A03829",
    x"1A0361C",
    x"1A0340E",
    x"1A03202",
    x"1A02FF5",
    x"1A02DEA",
    x"1A02BDE",
    x"1A029D4",
    x"1A027C9",
    x"1A025C0",
    x"1A023B7",
    x"1A021AE",
    x"1A01FA6",
    x"1A01D9E",
    x"1A01B97",
    x"1A01990",
    x"1A0178A",
    x"1A01584",
    x"1A0137F",
    x"1A0117B",
    x"1A00F77",
    x"1A00D73",
    x"1A00B70",
    x"1A0096D",
    x"1A0076B",
    x"1A0056A",
    x"1A00368",
    x"1A00168",
    x"19FFED0",
    x"19FFAD1",
    x"19FF6D3",
    x"19FF2D5",
    x"19FEED9",
    x"19FEADE",
    x"19FE6E4",
    x"19FE2EA",
    x"19FDEF2",
    x"19FDAFB",
    x"19FD705",
    x"19FD30F",
    x"19FCF1B",
    x"19FCB28",
    x"19FC736",
    x"19FC344",
    x"19FBF54",
    x"19FBB65",
    x"19FB776",
    x"19FB389",
    x"19FAF9D",
    x"19FABB1",
    x"19FA7C7",
    x"19FA3DD",
    x"19F9FF5",
    x"19F9C0D",
    x"19F9827",
    x"19F9441",
    x"19F905D",
    x"19F8C79",
    x"19F8896",
    x"19F84B5",
    x"19F80D4",
    x"19F7CF4",
    x"19F7915",
    x"19F7538",
    x"19F715B",
    x"19F6D7F",
    x"19F69A4",
    x"19F65CA",
    x"19F61F1",
    x"19F5E19",
    x"19F5A42",
    x"19F566C",
    x"19F5297",
    x"19F4EC3",
    x"19F4AF0",
    x"19F471D",
    x"19F434C",
    x"19F3F7C",
    x"19F3BAC",
    x"19F37DE",
    x"19F3410",
    x"19F3044",
    x"19F2C78",
    x"19F28AE",
    x"19F24E4",
    x"19F211B",
    x"19F1D53",
    x"19F198C",
    x"19F15C7",
    x"19F1202",
    x"19F0E3E",
    x"19F0A7A",
    x"19F06B8",
    x"19F02F7",
    x"19EFF37",
    x"19EFB77",
    x"19EF7B9",
    x"19EF3FC",
    x"19EF03F",
    x"19EEC84",
    x"19EE8C9",
    x"19EE50F",
    x"19EE156",
    x"19EDD9E",
    x"19ED9E8",
    x"19ED631",
    x"19ED27C",
    x"19ECEC8",
    x"19ECB15",
    x"19EC763",
    x"19EC3B1",
    x"19EC001",
    x"19EBC51",
    x"19EB8A3",
    x"19EB4F5",
    x"19EB148",
    x"19EAD9C",
    x"19EA9F1",
    x"19EA647",
    x"19EA29E",
    x"19E9EF6",
    x"19E9B4F",
    x"19E97A8",
    x"19E9403",
    x"19E905E",
    x"19E8CBB",
    x"19E8918",
    x"19E8576",
    x"19E81D5",
    x"19E7E35",
    x"19E7A96",
    x"19E76F8",
    x"19E735B",
    x"19E6FBE",
    x"19E6C23",
    x"19E6888",
    x"19E64EF",
    x"19E6156",
    x"19E5DBE",
    x"19E5A27",
    x"19E5691",
    x"19E52FC",
    x"19E4F67",
    x"19E4BD4",
    x"19E4841",
    x"19E44B0",
    x"19E411F",
    x"19E3D8F",
    x"19E3A00",
    x"19E3672",
    x"19E32E5",
    x"19E2F59",
    x"19E2BCD",
    x"19E2843",
    x"19E24B9",
    x"19E2131",
    x"19E1DA9",
    x"19E1A22",
    x"19E169C",
    x"19E1316",
    x"19E0F92",
    x"19E0C0F",
    x"19E088C",
    x"19E050A",
    x"19E018A",
    x"19DFE0A",
    x"19DFA8A",
    x"19DF70C",
    x"19DF38F",
    x"19DF013",
    x"19DEC97",
    x"19DE91C",
    x"19DE5A2",
    x"19DE229",
    x"19DDEB1",
    x"19DDB3A",
    x"19DD7C4",
    x"19DD44E",
    x"19DD0DA",
    x"19DCD66",
    x"19DC9F3",
    x"19DC681",
    x"19DC310",
    x"19DBF9F",
    x"19DBC30",
    x"19DB8C1",
    x"19DB553",
    x"19DB1E6",
    x"19DAE7A",
    x"19DAB0F",
    x"19DA7A5",
    x"19DA43B",
    x"19DA0D3",
    x"19D9D6B",
    x"19D9A04",
    x"19D969E",
    x"19D9339",
    x"19D8FD4",
    x"19D8C71",
    x"19D890E",
    x"19D85AC",
    x"19D824B",
    x"19D7EEB",
    x"19D7B8C",
    x"19D782D",
    x"19D74D0",
    x"19D7173",
    x"19D6E17",
    x"19D6ABC",
    x"19D6762",
    x"19D6408",
    x"19D60B0",
    x"19D5D58",
    x"19D5A01",
    x"19D56AB",
    x"19D5356",
    x"19D5001",
    x"19D4CAE",
    x"19D495B",
    x"19D4609",
    x"19D42B8",
    x"19D3F68",
    x"19D3C18",
    x"19D38CA",
    x"19D357C",
    x"19D322F",
    x"19D2EE3",
    x"19D2B97",
    x"19D284D",
    x"19D2503",
    x"19D21BA",
    x"19D1E72",
    x"19D1B2B",
    x"19D17E5",
    x"19D149F",
    x"19D115A",
    x"19D0E17",
    x"19D0AD3",
    x"19D0791",
    x"19D0450",
    x"19D010F",
    x"19CFDCF",
    x"19CFA90",
    x"19CF752",
    x"19CF414",
    x"19CF0D8",
    x"19CED9C",
    x"19CEA61",
    x"19CE727",
    x"19CE3ED",
    x"19CE0B5",
    x"19CDD7D",
    x"19CDA46",
    x"19CD710",
    x"19CD3DB",
    x"19CD0A6",
    x"19CCD72",
    x"19CCA3F",
    x"19CC70D",
    x"19CC3DC",
    x"19CC0AB",
    x"19CBD7B",
    x"19CBA4C",
    x"19CB71E",
    x"19CB3F1",
    x"19CB0C4",
    x"19CAD98",
    x"19CAA6D",
    x"19CA743",
    x"19CA41A",
    x"19CA0F1",
    x"19C9DC9",
    x"19C9AA2",
    x"19C977C",
    x"19C9457",
    x"19C9132",
    x"19C8E0E",
    x"19C8AEB",
    x"19C87C9",
    x"19C84A7",
    x"19C8186",
    x"19C7E66",
    x"19C7B47",
    x"19C7829",
    x"19C750B",
    x"19C71EE",
    x"19C6ED2",
    x"19C6BB7",
    x"19C689C",
    x"19C6582",
    x"19C6269",
    x"19C5F51",
    x"19C5C3A",
    x"19C5923",
    x"19C560D",
    x"19C52F8",
    x"19C4FE4",
    x"19C4CD0",
    x"19C49BD",
    x"19C46AB",
    x"19C439A",
    x"19C4089",
    x"19C3D7A",
    x"19C3A6B",
    x"19C375C",
    x"19C344F",
    x"19C3142",
    x"19C2E36",
    x"19C2B2B",
    x"19C2821",
    x"19C2517",
    x"19C220E",
    x"19C1F06",
    x"19C1BFF",
    x"19C18F8",
    x"19C15F2",
    x"19C12ED",
    x"19C0FE9",
    x"19C0CE5",
    x"19C09E2",
    x"19C06E0",
    x"19C03DF",
    x"19C00DE",
    x"19BFDDE",
    x"19BFADF",
    x"19BF7E1",
    x"19BF4E3",
    x"19BF1E6",
    x"19BEEEA",
    x"19BEBEF",
    x"19BE8F4",
    x"19BE5FB",
    x"19BE301",
    x"19BE009",
    x"19BDD11",
    x"19BDA1B",
    x"19BD724",
    x"19BD42F",
    x"19BD13A",
    x"19BCE46",
    x"19BCB53",
    x"19BC861",
    x"19BC56F",
    x"19BC27E",
    x"19BBF8E",
    x"19BBC9E",
    x"19BB9AF",
    x"19BB6C1",
    x"19BB3D4",
    x"19BB0E7",
    x"19BADFC",
    x"19BAB10",
    x"19BA826",
    x"19BA53C",
    x"19BA253",
    x"19B9F6B",
    x"19B9C84",
    x"19B999D",
    x"19B96B7",
    x"19B93D2",
    x"19B90ED",
    x"19B8E09",
    x"19B8B26",
    x"19B8844",
    x"19B8562",
    x"19B8281",
    x"19B7FA1",
    x"19B7CC1",
    x"19B79E2",
    x"19B7704",
    x"19B7427",
    x"19B714A",
    x"19B6E6E",
    x"19B6B93",
    x"19B68B8",
    x"19B65DE",
    x"19B6305",
    x"19B602D",
    x"19B5D55",
    x"19B5A7E",
    x"19B57A8",
    x"19B54D2",
    x"19B51FE",
    x"19B4F29",
    x"19B4C56",
    x"19B4983",
    x"19B46B1",
    x"19B43E0",
    x"19B410F",
    x"19B3E3F",
    x"19B3B70",
    x"19B38A2",
    x"19B35D4",
    x"19B3307",
    x"19B303A",
    x"19B2D6F",
    x"19B2AA4",
    x"19B27D9",
    x"19B2510",
    x"19B2247",
    x"19B1F7F",
    x"19B1CB7",
    x"19B19F0",
    x"19B172A",
    x"19B1465",
    x"19B11A0",
    x"19B0EDC",
    x"19B0C18",
    x"19B0956",
    x"19B0694",
    x"19B03D2",
    x"19B0112",
    x"19AFE52",
    x"19AFB93",
    x"19AF8D4",
    x"19AF616",
    x"19AF359",
    x"19AF09D",
    x"19AEDE1",
    x"19AEB26",
    x"19AE86B",
    x"19AE5B1",
    x"19AE2F8",
    x"19AE040",
    x"19ADD88",
    x"19ADAD1",
    x"19AD81B",
    x"19AD565",
    x"19AD2B0",
    x"19ACFFC",
    x"19ACD48",
    x"19ACA95",
    x"19AC7E3",
    x"19AC531",
    x"19AC280",
    x"19ABFD0",
    x"19ABD20",
    x"19ABA71",
    x"19AB7C3",
    x"19AB515",
    x"19AB269",
    x"19AAFBC",
    x"19AAD11",
    x"19AAA66",
    x"19AA7BB",
    x"19AA512",
    x"19AA269",
    x"19A9FC1",
    x"19A9D19",
    x"19A9A72",
    x"19A97CC",
    x"19A9526",
    x"19A9281",
    x"19A8FDD",
    x"19A8D39",
    x"19A8A96",
    x"19A87F4",
    x"19A8552",
    x"19A82B1",
    x"19A8011",
    x"19A7D71",
    x"19A7AD2",
    x"19A7834",
    x"19A7596",
    x"19A72F9",
    x"19A705D",
    x"19A6DC1",
    x"19A6B26",
    x"19A688B",
    x"19A65F2",
    x"19A6358",
    x"19A60C0",
    x"19A5E28",
    x"19A5B91",
    x"19A58FA",
    x"19A5664",
    x"19A53CF",
    x"19A513A",
    x"19A4EA6",
    x"19A4C13",
    x"19A4980",
    x"19A46EE",
    x"19A445D",
    x"19A41CC",
    x"19A3F3C",
    x"19A3CAD",
    x"19A3A1E",
    x"19A378F",
    x"19A3502",
    x"19A3275",
    x"19A2FE9",
    x"19A2D5D",
    x"19A2AD2",
    x"19A2848",
    x"19A25BE",
    x"19A2335",
    x"19A20AC",
    x"19A1E24",
    x"19A1B9D",
    x"19A1917",
    x"19A1691",
    x"19A140B",
    x"19A1187",
    x"19A0F03",
    x"19A0C7F",
    x"19A09FC",
    x"19A077A",
    x"19A04F9",
    x"19A0278",
    x"199FFF7",
    x"199FD78",
    x"199FAF9",
    x"199F87A",
    x"199F5FC",
    x"199F37F",
    x"199F103",
    x"199EE87",
    x"199EC0B",
    x"199E991",
    x"199E717",
    x"199E49D",
    x"199E224",
    x"199DFAC",
    x"199DD34",
    x"199DABD",
    x"199D847",
    x"199D5D1",
    x"199D35C",
    x"199D0E8",
    x"199CE74",
    x"199CC00",
    x"199C98E",
    x"199C71C",
    x"199C4AA",
    x"199C239",
    x"199BFC9",
    x"199BD59",
    x"199BAEA",
    x"199B87C",
    x"199B60E",
    x"199B3A1",
    x"199B134",
    x"199AEC8",
    x"199AC5D",
    x"199A9F2",
    x"199A788",
    x"199A51E",
    x"199A2B5",
    x"199A04D",
    x"1999DE5",
    x"1999B7E",
    x"1999917",
    x"19996B1",
    x"199944C",
    x"19991E7",
    x"1998F83",
    x"1998D20",
    x"1998ABD",
    x"199885A",
    x"19985F8",
    x"1998397",
    x"1998137",
    x"1997ED7",
    x"1997C77",
    x"1997A18",
    x"19977BA",
    x"199755D",
    x"19972FF",
    x"19970A3",
    x"1996E47",
    x"1996BEC",
    x"1996991",
    x"1996737",
    x"19964DE",
    x"1996285",
    x"199602C",
    x"1995DD5",
    x"1995B7D",
    x"1995927",
    x"19956D1",
    x"199547B",
    x"1995227",
    x"1994FD2",
    x"1994D7F",
    x"1994B2C",
    x"19948D9",
    x"1994687",
    x"1994436",
    x"19941E5",
    x"1993F95",
    x"1993D45",
    x"1993AF6",
    x"19938A8",
    x"199365A",
    x"199340D",
    x"19931C0",
    x"1992F74",
    x"1992D28",
    x"1992ADD",
    x"1992893",
    x"1992649",
    x"1992400",
    x"19921B7",
    x"1991F6F",
    x"1991D27",
    x"1991AE0",
    x"199189A",
    x"1991654",
    x"199140F",
    x"19911CA",
    x"1990F86",
    x"1990D42",
    x"1990AFF",
    x"19908BD",
    x"199067B",
    x"1990439",
    x"19901F9",
    x"198FFB8",
    x"198FD79",
    x"198FB3A",
    x"198F8FB",
    x"198F6BD",
    x"198F480",
    x"198F243",
    x"198F007",
    x"198EDCB",
    x"198EB90",
    x"198E955",
    x"198E71B",
    x"198E4E1",
    x"198E2A9",
    x"198E070",
    x"198DE38",
    x"198DC01",
    x"198D9CA",
    x"198D794",
    x"198D55F",
    x"198D329",
    x"198D0F5",
    x"198CEC1",
    x"198CC8E",
    x"198CA5B",
    x"198C828",
    x"198C5F7",
    x"198C3C5",
    x"198C195",
    x"198BF65",
    x"198BD35",
    x"198BB06",
    x"198B8D8",
    x"198B6AA",
    x"198B47C",
    x"198B24F",
    x"198B023",
    x"198ADF7",
    x"198ABCC",
    x"198A9A1",
    x"198A777",
    x"198A54E",
    x"198A325",
    x"198A0FC",
    x"1989ED4",
    x"1989CAD",
    x"1989A86",
    x"198985F",
    x"198963A",
    x"1989414",
    x"19891F0",
    x"1988FCB",
    x"1988DA8",
    x"1988B84",
    x"1988962",
    x"1988740",
    x"198851E",
    x"19882FD",
    x"19880DD",
    x"1987EBD",
    x"1987C9D",
    x"1987A7E",
    x"1987860",
    x"1987642",
    x"1987425",
    x"1987208",
    x"1986FEC",
    x"1986DD0",
    x"1986BB5",
    x"198699A",
    x"1986780",
    x"1986567",
    x"198634E",
    x"1986135",
    x"1985F1D",
    x"1985D05",
    x"1985AEE",
    x"19858D8",
    x"19856C2",
    x"19854AD",
    x"1985298",
    x"1985083",
    x"1984E6F",
    x"1984C5C",
    x"1984A49",
    x"1984837",
    x"1984625",
    x"1984414",
    x"1984203",
    x"1983FF3",
    x"1983DE3",
    x"1983BD4",
    x"19839C5",
    x"19837B7",
    x"19835A9",
    x"198339C",
    x"1983190",
    x"1982F83",
    x"1982D78",
    x"1982B6D",
    x"1982962",
    x"1982758",
    x"198254E",
    x"1982345",
    x"198213D",
    x"1981F35",
    x"1981D2D",
    x"1981B26",
    x"1981920",
    x"198171A",
    x"1981514",
    x"198130F",
    x"198110B",
    x"1980F07",
    x"1980D03",
    x"1980B00",
    x"19808FD",
    x"19806FB",
    x"19804FA",
    x"19802F9",
    x"19800F9",
    x"197FDF2",
    x"197F9F3",
    x"197F5F5",
    x"197F1F8",
    x"197EDFC",
    x"197EA01",
    x"197E607",
    x"197E20E",
    x"197DE16",
    x"197DA1E",
    x"197D628",
    x"197D233",
    x"197CE3F",
    x"197CA4C",
    x"197C65A",
    x"197C269",
    x"197BE79",
    x"197BA8A",
    x"197B69C",
    x"197B2AF",
    x"197AEC2",
    x"197AAD7",
    x"197A6ED",
    x"197A304",
    x"1979F1B",
    x"1979B34",
    x"197974E",
    x"1979369",
    x"1978F84",
    x"1978BA1",
    x"19787BE",
    x"19783DD",
    x"1977FFC",
    x"1977C1D",
    x"197783E",
    x"1977461",
    x"1977084",
    x"1976CA9",
    x"19768CE",
    x"19764F4",
    x"197611B",
    x"1975D44",
    x"197596D",
    x"1975597",
    x"19751C2",
    x"1974DEE",
    x"1974A1B",
    x"1974649",
    x"1974278",
    x"1973EA8",
    x"1973AD8",
    x"197370A",
    x"197333D",
    x"1972F71",
    x"1972BA5",
    x"19727DB",
    x"1972411",
    x"1972049",
    x"1971C81",
    x"19718BB",
    x"19714F5",
    x"1971130",
    x"1970D6C",
    x"19709A9",
    x"19705E7",
    x"1970226",
    x"196FE66",
    x"196FAA7",
    x"196F6E9",
    x"196F32C",
    x"196EF6F",
    x"196EBB4",
    x"196E7FA",
    x"196E440",
    x"196E087",
    x"196DCD0",
    x"196D919",
    x"196D563",
    x"196D1AE",
    x"196CDFA",
    x"196CA47",
    x"196C695",
    x"196C2E4",
    x"196BF34",
    x"196BB84",
    x"196B7D6",
    x"196B428",
    x"196B07C",
    x"196ACD0",
    x"196A926",
    x"196A57C",
    x"196A1D3",
    x"1969E2B",
    x"1969A84",
    x"19696DE",
    x"1969338",
    x"1968F94",
    x"1968BF0",
    x"196884E",
    x"19684AC",
    x"196810C",
    x"1967D6C",
    x"19679CD",
    x"196762F",
    x"1967292",
    x"1966EF6",
    x"1966B5A",
    x"19667C0",
    x"1966426",
    x"196608E",
    x"1965CF6",
    x"196595F",
    x"19655C9",
    x"1965234",
    x"1964EA0",
    x"1964B0D",
    x"196477B",
    x"19643E9",
    x"1964059",
    x"1963CC9",
    x"196393A",
    x"19635AD",
    x"1963220",
    x"1962E94",
    x"1962B08",
    x"196277E",
    x"19623F5",
    x"196206C",
    x"1961CE4",
    x"196195E",
    x"19615D8",
    x"1961253",
    x"1960ECF",
    x"1960B4B",
    x"19607C9",
    x"1960447",
    x"19600C7",
    x"195FD47",
    x"195F9C8",
    x"195F64A",
    x"195F2CD",
    x"195EF51",
    x"195EBD5",
    x"195E85B",
    x"195E4E1",
    x"195E168",
    x"195DDF0",
    x"195DA79",
    x"195D703",
    x"195D38E",
    x"195D019",
    x"195CCA6",
    x"195C933",
    x"195C5C1",
    x"195C250",
    x"195BEE0",
    x"195BB71",
    x"195B802",
    x"195B495",
    x"195B128",
    x"195ADBC",
    x"195AA51",
    x"195A6E7",
    x"195A37E",
    x"195A015",
    x"1959CAE",
    x"1959947",
    x"19595E1",
    x"195927C",
    x"1958F18",
    x"1958BB4",
    x"1958852",
    x"19584F0",
    x"195818F",
    x"1957E30",
    x"1957AD0",
    x"1957772",
    x"1957415",
    x"19570B8",
    x"1956D5C",
    x"1956A01",
    x"19566A7",
    x"195634E",
    x"1955FF6",
    x"1955C9E",
    x"1955947",
    x"19555F1",
    x"195529C",
    x"1954F48",
    x"1954BF5",
    x"19548A2",
    x"1954550",
    x"19541FF",
    x"1953EAF",
    x"1953B60",
    x"1953812",
    x"19534C4",
    x"1953177",
    x"1952E2B",
    x"1952AE0",
    x"1952796",
    x"195244C",
    x"1952104",
    x"1951DBC",
    x"1951A75",
    x"195172F",
    x"19513E9",
    x"19510A5",
    x"1950D61",
    x"1950A1E",
    x"19506DC",
    x"195039B",
    x"195005A",
    x"194FD1A",
    x"194F9DC",
    x"194F69E",
    x"194F360",
    x"194F024",
    x"194ECE8",
    x"194E9AD",
    x"194E673",
    x"194E33A",
    x"194E002",
    x"194DCCA",
    x"194D993",
    x"194D65D",
    x"194D328",
    x"194CFF4",
    x"194CCC0",
    x"194C98D",
    x"194C65B",
    x"194C32A",
    x"194BFFA",
    x"194BCCA",
    x"194B99B",
    x"194B66D",
    x"194B340",
    x"194B014",
    x"194ACE8",
    x"194A9BD",
    x"194A693",
    x"194A36A",
    x"194A042",
    x"1949D1A",
    x"19499F3",
    x"19496CD",
    x"19493A8",
    x"1949083",
    x"1948D5F",
    x"1948A3C",
    x"194871A",
    x"19483F9",
    x"19480D8",
    x"1947DB8",
    x"1947A99",
    x"194777B",
    x"194745E",
    x"1947141",
    x"1946E25",
    x"1946B0A",
    x"19467F0",
    x"19464D6",
    x"19461BD",
    x"1945EA5",
    x"1945B8E",
    x"1945877",
    x"1945562",
    x"194524D",
    x"1944F38",
    x"1944C25",
    x"1944912",
    x"1944600",
    x"19442EF",
    x"1943FDF",
    x"1943CCF",
    x"19439C1",
    x"19436B3",
    x"19433A5",
    x"1943099",
    x"1942D8D",
    x"1942A82",
    x"1942778",
    x"194246E",
    x"1942165",
    x"1941E5D",
    x"1941B56",
    x"1941850",
    x"194154A",
    x"1941245",
    x"1940F41",
    x"1940C3E",
    x"194093B",
    x"1940639",
    x"1940338",
    x"1940037",
    x"193FD38",
    x"193FA39",
    x"193F73B",
    x"193F43D",
    x"193F140",
    x"193EE44",
    x"193EB49",
    x"193E84F",
    x"193E555",
    x"193E25C",
    x"193DF64",
    x"193DC6C",
    x"193D976",
    x"193D680",
    x"193D38A",
    x"193D096",
    x"193CDA2",
    x"193CAAF",
    x"193C7BD",
    x"193C4CB",
    x"193C1DA",
    x"193BEEA",
    x"193BBFB",
    x"193B90C",
    x"193B61E",
    x"193B331",
    x"193B045",
    x"193AD59",
    x"193AA6E",
    x"193A784",
    x"193A49A",
    x"193A1B2",
    x"1939ECA",
    x"1939BE2",
    x"19398FC",
    x"1939616",
    x"1939331",
    x"193904C",
    x"1938D68",
    x"1938A85",
    x"19387A3",
    x"19384C2",
    x"19381E1",
    x"1937F01",
    x"1937C21",
    x"1937943",
    x"1937665",
    x"1937387",
    x"19370AB",
    x"1936DCF",
    x"1936AF4",
    x"193681A",
    x"1936540",
    x"1936267",
    x"1935F8F",
    x"1935CB7",
    x"19359E0",
    x"193570A",
    x"1935435",
    x"1935160",
    x"1934E8C",
    x"1934BB9",
    x"19348E6",
    x"1934614",
    x"1934343",
    x"1934073",
    x"1933DA3",
    x"1933AD4",
    x"1933806",
    x"1933538",
    x"193326B",
    x"1932F9F",
    x"1932CD3",
    x"1932A08",
    x"193273E",
    x"1932475",
    x"19321AC",
    x"1931EE4",
    x"1931C1C",
    x"1931956",
    x"1931690",
    x"19313CB",
    x"1931106",
    x"1930E42",
    x"1930B7F",
    x"19308BC",
    x"19305FA",
    x"1930339",
    x"1930079",
    x"192FDB9",
    x"192FAFA",
    x"192F83C",
    x"192F57E",
    x"192F2C1",
    x"192F004",
    x"192ED49",
    x"192EA8E",
    x"192E7D4",
    x"192E51A",
    x"192E261",
    x"192DFA9",
    x"192DCF1",
    x"192DA3A",
    x"192D784",
    x"192D4CE",
    x"192D21A",
    x"192CF65",
    x"192CCB2",
    x"192C9FF",
    x"192C74D",
    x"192C49B",
    x"192C1EB",
    x"192BF3A",
    x"192BC8B",
    x"192B9DC",
    x"192B72E",
    x"192B481",
    x"192B1D4",
    x"192AF28",
    x"192AC7C",
    x"192A9D1",
    x"192A727",
    x"192A47E",
    x"192A1D5",
    x"1929F2D",
    x"1929C85",
    x"19299DF",
    x"1929739",
    x"1929493",
    x"19291EE",
    x"1928F4A",
    x"1928CA7",
    x"1928A04",
    x"1928762",
    x"19284C0",
    x"192821F",
    x"1927F7F",
    x"1927CDF",
    x"1927A41",
    x"19277A2",
    x"1927505",
    x"1927268",
    x"1926FCC",
    x"1926D30",
    x"1926A95",
    x"19267FB",
    x"1926561",
    x"19262C8",
    x"1926030",
    x"1925D98",
    x"1925B01",
    x"192586A",
    x"19255D5",
    x"192533F",
    x"19250AB",
    x"1924E17",
    x"1924B84",
    x"19248F1",
    x"192465F",
    x"19243CE",
    x"192413E",
    x"1923EAE",
    x"1923C1E",
    x"192398F",
    x"1923701",
    x"1923474",
    x"19231E7",
    x"1922F5B",
    x"1922CD0",
    x"1922A45",
    x"19227BA",
    x"1922531",
    x"19222A8",
    x"192201F",
    x"1921D98",
    x"1921B11",
    x"192188A",
    x"1921604",
    x"192137F",
    x"19210FB",
    x"1920E77",
    x"1920BF3",
    x"1920971",
    x"19206EF",
    x"192046D",
    x"19201EC",
    x"191FF6C",
    x"191FCED",
    x"191FA6E",
    x"191F7F0",
    x"191F572",
    x"191F2F5",
    x"191F078",
    x"191EDFD",
    x"191EB81",
    x"191E907",
    x"191E68D",
    x"191E414",
    x"191E19B",
    x"191DF23",
    x"191DCAB",
    x"191DA34",
    x"191D7BE",
    x"191D549",
    x"191D2D4",
    x"191D05F",
    x"191CDEB",
    x"191CB78",
    x"191C906",
    x"191C694",
    x"191C422",
    x"191C1B2",
    x"191BF41",
    x"191BCD2",
    x"191BA63",
    x"191B7F5",
    x"191B587",
    x"191B31A",
    x"191B0AE",
    x"191AE42",
    x"191ABD6",
    x"191A96C",
    x"191A702",
    x"191A498",
    x"191A22F",
    x"1919FC7",
    x"1919D5F",
    x"1919AF8",
    x"1919892",
    x"191962C",
    x"19193C7",
    x"1919162",
    x"1918EFE",
    x"1918C9B",
    x"1918A38",
    x"19187D6",
    x"1918574",
    x"1918313",
    x"19180B2",
    x"1917E53",
    x"1917BF3",
    x"1917995",
    x"1917736",
    x"19174D9",
    x"191727C",
    x"1917020",
    x"1916DC4",
    x"1916B69",
    x"191690E",
    x"19166B4",
    x"191645B",
    x"1916202",
    x"1915FAA",
    x"1915D52",
    x"1915AFB",
    x"19158A5",
    x"191564F",
    x"19153FA",
    x"19151A5",
    x"1914F51",
    x"1914CFD",
    x"1914AAA",
    x"1914858",
    x"1914606",
    x"19143B5",
    x"1914164",
    x"1913F14",
    x"1913CC5",
    x"1913A76",
    x"1913828",
    x"19135DA",
    x"191338D",
    x"1913140",
    x"1912EF4",
    x"1912CA9",
    x"1912A5E",
    x"1912813",
    x"19125CA",
    x"1912380",
    x"1912138",
    x"1911EF0",
    x"1911CA8",
    x"1911A62",
    x"191181B",
    x"19115D5",
    x"1911390",
    x"191114C",
    x"1910F08",
    x"1910CC4",
    x"1910A81",
    x"191083F",
    x"19105FD",
    x"19103BC",
    x"191017B",
    x"190FF3B",
    x"190FCFC",
    x"190FABD",
    x"190F87E",
    x"190F640",
    x"190F403",
    x"190F1C6",
    x"190EF8A",
    x"190ED4F",
    x"190EB14",
    x"190E8D9",
    x"190E69F",
    x"190E466",
    x"190E22D",
    x"190DFF5",
    x"190DDBD",
    x"190DB86",
    x"190D94F",
    x"190D719",
    x"190D4E4",
    x"190D2AF",
    x"190D07A",
    x"190CE47",
    x"190CC13",
    x"190C9E0",
    x"190C7AE",
    x"190C57D",
    x"190C34C",
    x"190C11B",
    x"190BEEB",
    x"190BCBC",
    x"190BA8D",
    x"190B85E",
    x"190B630",
    x"190B403",
    x"190B1D6",
    x"190AFAA",
    x"190AD7F",
    x"190AB53",
    x"190A929",
    x"190A6FF",
    x"190A4D5",
    x"190A2AC",
    x"190A084",
    x"1909E5C",
    x"1909C35",
    x"1909A0E",
    x"19097E8",
    x"19095C2",
    x"190939D",
    x"1909178",
    x"1908F54",
    x"1908D31",
    x"1908B0E",
    x"19088EB",
    x"19086C9",
    x"19084A8",
    x"1908287",
    x"1908067",
    x"1907E47",
    x"1907C27",
    x"1907A09",
    x"19077EA",
    x"19075CD",
    x"19073AF",
    x"1907193",
    x"1906F77",
    x"1906D5B",
    x"1906B40",
    x"1906925",
    x"190670B",
    x"19064F2",
    x"19062D9",
    x"19060C0",
    x"1905EA9",
    x"1905C91",
    x"1905A7A",
    x"1905864",
    x"190564E",
    x"1905439",
    x"1905224",
    x"1905010",
    x"1904DFC",
    x"1904BE9",
    x"19049D6",
    x"19047C4",
    x"19045B2",
    x"19043A1",
    x"1904190",
    x"1903F80",
    x"1903D71",
    x"1903B61",
    x"1903953",
    x"1903745",
    x"1903537",
    x"190332A",
    x"190311E",
    x"1902F12",
    x"1902D06",
    x"1902AFB",
    x"19028F1",
    x"19026E7",
    x"19024DD",
    x"19022D4",
    x"19020CC",
    x"1901EC4",
    x"1901CBC",
    x"1901AB5",
    x"19018AF",
    x"19016A9",
    x"19014A4",
    x"190129F",
    x"190109A",
    x"1900E96",
    x"1900C93",
    x"1900A90",
    x"190088E",
    x"190068C",
    x"190048A",
    x"190028A",
    x"1900089",
    x"18FFD13",
    x"18FF914",
    x"18FF517",
    x"18FF11A",
    x"18FED1E",
    x"18FE923",
    x"18FE529",
    x"18FE131",
    x"18FDD39",
    x"18FD942",
    x"18FD54C",
    x"18FD157",
    x"18FCD64",
    x"18FC971",
    x"18FC57F",
    x"18FC18E",
    x"18FBD9E",
    x"18FB9AF",
    x"18FB5C1",
    x"18FB1D4",
    x"18FADE8",
    x"18FA9FD",
    x"18FA613",
    x"18FA22A",
    x"18F9E42",
    x"18F9A5B",
    x"18F9675",
    x"18F9290",
    x"18F8EAC",
    x"18F8AC9",
    x"18F86E6",
    x"18F8305",
    x"18F7F25",
    x"18F7B46",
    x"18F7767",
    x"18F738A",
    x"18F6FAD",
    x"18F6BD2",
    x"18F67F8",
    x"18F641E",
    x"18F6045",
    x"18F5C6E",
    x"18F5897",
    x"18F54C2",
    x"18F50ED",
    x"18F4D19",
    x"18F4946",
    x"18F4575",
    x"18F41A4",
    x"18F3DD4",
    x"18F3A05",
    x"18F3637",
    x"18F326A",
    x"18F2E9D",
    x"18F2AD2",
    x"18F2708",
    x"18F233F",
    x"18F1F76",
    x"18F1BAF",
    x"18F17E9",
    x"18F1423",
    x"18F105F",
    x"18F0C9B",
    x"18F08D8",
    x"18F0516",
    x"18F0156",
    x"18EFD96",
    x"18EF9D7",
    x"18EF619",
    x"18EF25C",
    x"18EEEA0",
    x"18EEAE5",
    x"18EE72A",
    x"18EE371",
    x"18EDFB9",
    x"18EDC01",
    x"18ED84B",
    x"18ED495",
    x"18ED0E0",
    x"18ECD2C",
    x"18EC97A",
    x"18EC5C8",
    x"18EC217",
    x"18EBE67",
    x"18EBAB8",
    x"18EB709",
    x"18EB35C",
    x"18EAFB0",
    x"18EAC04",
    x"18EA85A",
    x"18EA4B0",
    x"18EA107",
    x"18E9D60",
    x"18E99B9",
    x"18E9613",
    x"18E926E",
    x"18E8EC9",
    x"18E8B26",
    x"18E8784",
    x"18E83E2",
    x"18E8042",
    x"18E7CA2",
    x"18E7904",
    x"18E7566",
    x"18E71C9",
    x"18E6E2D",
    x"18E6A92",
    x"18E66F8",
    x"18E635E",
    x"18E5FC6",
    x"18E5C2E",
    x"18E5898",
    x"18E5502",
    x"18E516D",
    x"18E4DD9",
    x"18E4A46",
    x"18E46B4",
    x"18E4323",
    x"18E3F93",
    x"18E3C03",
    x"18E3875",
    x"18E34E7",
    x"18E315A",
    x"18E2DCE",
    x"18E2A43",
    x"18E26B9",
    x"18E2330",
    x"18E1FA8",
    x"18E1C20",
    x"18E189A",
    x"18E1514",
    x"18E118F",
    x"18E0E0B",
    x"18E0A88",
    x"18E0706",
    x"18E0384",
    x"18E0004",
    x"18DFC84",
    x"18DF906",
    x"18DF588",
    x"18DF20B",
    x"18DEE8F",
    x"18DEB14",
    x"18DE799",
    x"18DE420",
    x"18DE0A7",
    x"18DDD30",
    x"18DD9B9",
    x"18DD643",
    x"18DD2CE",
    x"18DCF59",
    x"18DCBE6",
    x"18DC873",
    x"18DC502",
    x"18DC191",
    x"18DBE21",
    x"18DBAB2",
    x"18DB744",
    x"18DB3D6",
    x"18DB06A",
    x"18DACFE",
    x"18DA993",
    x"18DA629",
    x"18DA2C0",
    x"18D9F58",
    x"18D9BF0",
    x"18D988A",
    x"18D9524",
    x"18D91BF",
    x"18D8E5B",
    x"18D8AF8",
    x"18D8796",
    x"18D8434",
    x"18D80D4",
    x"18D7D74",
    x"18D7A15",
    x"18D76B7",
    x"18D735A",
    x"18D6FFD",
    x"18D6CA2",
    x"18D6947",
    x"18D65ED",
    x"18D6294",
    x"18D5F3C",
    x"18D5BE4",
    x"18D588E",
    x"18D5538",
    x"18D51E3",
    x"18D4E8F",
    x"18D4B3C",
    x"18D47E9",
    x"18D4498",
    x"18D4147",
    x"18D3DF7",
    x"18D3AA8",
    x"18D375A",
    x"18D340C",
    x"18D30C0",
    x"18D2D74",
    x"18D2A29",
    x"18D26DF",
    x"18D2396",
    x"18D204D",
    x"18D1D06",
    x"18D19BF",
    x"18D1679",
    x"18D1333",
    x"18D0FEF",
    x"18D0CAC",
    x"18D0969",
    x"18D0627",
    x"18D02E6",
    x"18CFFA5",
    x"18CFC66",
    x"18CF927",
    x"18CF5E9",
    x"18CF2AC",
    x"18CEF70",
    x"18CEC34",
    x"18CE8FA",
    x"18CE5C0",
    x"18CE287",
    x"18CDF4F",
    x"18CDC17",
    x"18CD8E1",
    x"18CD5AB",
    x"18CD276",
    x"18CCF42",
    x"18CCC0E",
    x"18CC8DC",
    x"18CC5AA",
    x"18CC279",
    x"18CBF49",
    x"18CBC19",
    x"18CB8EA",
    x"18CB5BD",
    x"18CB290",
    x"18CAF63",
    x"18CAC38",
    x"18CA90D",
    x"18CA5E3",
    x"18CA2BA",
    x"18C9F92",
    x"18C9C6B",
    x"18C9944",
    x"18C961E",
    x"18C92F9",
    x"18C8FD4",
    x"18C8CB1",
    x"18C898E",
    x"18C866C",
    x"18C834B",
    x"18C802A",
    x"18C7D0B",
    x"18C79EC",
    x"18C76CE",
    x"18C73B0",
    x"18C7094",
    x"18C6D78",
    x"18C6A5D",
    x"18C6743",
    x"18C642A",
    x"18C6111",
    x"18C5DF9",
    x"18C5AE2",
    x"18C57CC",
    x"18C54B6",
    x"18C51A1",
    x"18C4E8D",
    x"18C4B7A",
    x"18C4867",
    x"18C4556",
    x"18C4245",
    x"18C3F35",
    x"18C3C25",
    x"18C3917",
    x"18C3609",
    x"18C32FC",
    x"18C2FEF",
    x"18C2CE4",
    x"18C29D9",
    x"18C26CF",
    x"18C23C5",
    x"18C20BD",
    x"18C1DB5",
    x"18C1AAE",
    x"18C17A8",
    x"18C14A2",
    x"18C119D",
    x"18C0E99",
    x"18C0B96",
    x"18C0893",
    x"18C0592",
    x"18C0291",
    x"18BFF90",
    x"18BFC91",
    x"18BF992",
    x"18BF694",
    x"18BF397",
    x"18BF09A",
    x"18BED9F",
    x"18BEAA4",
    x"18BE7A9",
    x"18BE4B0",
    x"18BE1B7",
    x"18BDEBF",
    x"18BDBC8",
    x"18BD8D1",
    x"18BD5DB",
    x"18BD2E6",
    x"18BCFF2",
    x"18BCCFE",
    x"18BCA0B",
    x"18BC719",
    x"18BC428",
    x"18BC137",
    x"18BBE47",
    x"18BBB58",
    x"18BB869",
    x"18BB57C",
    x"18BB28F",
    x"18BAFA2",
    x"18BACB7",
    x"18BA9CC",
    x"18BA6E2",
    x"18BA3F9",
    x"18BA110",
    x"18B9E28",
    x"18B9B41",
    x"18B985A",
    x"18B9575",
    x"18B9290",
    x"18B8FAB",
    x"18B8CC8",
    x"18B89E5",
    x"18B8703",
    x"18B8421",
    x"18B8141",
    x"18B7E61",
    x"18B7B82",
    x"18B78A3",
    x"18B75C5",
    x"18B72E8",
    x"18B700C",
    x"18B6D30",
    x"18B6A55",
    x"18B677B",
    x"18B64A1",
    x"18B61C9",
    x"18B5EF1",
    x"18B5C19",
    x"18B5943",
    x"18B566D",
    x"18B5397",
    x"18B50C3",
    x"18B4DEF",
    x"18B4B1C",
    x"18B4849",
    x"18B4578",
    x"18B42A7",
    x"18B3FD6",
    x"18B3D07",
    x"18B3A38",
    x"18B376A",
    x"18B349C",
    x"18B31CF",
    x"18B2F03",
    x"18B2C38",
    x"18B296D",
    x"18B26A3",
    x"18B23DA",
    x"18B2111",
    x"18B1E49",
    x"18B1B82",
    x"18B18BB",
    x"18B15F6",
    x"18B1331",
    x"18B106C",
    x"18B0DA8",
    x"18B0AE5",
    x"18B0823",
    x"18B0561",
    x"18B02A0",
    x"18AFFE0",
    x"18AFD20",
    x"18AFA61",
    x"18AF7A3",
    x"18AF4E5",
    x"18AF229",
    x"18AEF6C",
    x"18AECB1",
    x"18AE9F6",
    x"18AE73C",
    x"18AE482",
    x"18AE1CA",
    x"18ADF12",
    x"18ADC5A",
    x"18AD9A3",
    x"18AD6ED",
    x"18AD438",
    x"18AD183",
    x"18ACECF",
    x"18ACC1C",
    x"18AC969",
    x"18AC6B7",
    x"18AC406",
    x"18AC155",
    x"18ABEA5",
    x"18ABBF6",
    x"18AB947",
    x"18AB699",
    x"18AB3EC",
    x"18AB13F",
    x"18AAE93",
    x"18AABE8",
    x"18AA93D",
    x"18AA693",
    x"18AA3EA",
    x"18AA141",
    x"18A9E99",
    x"18A9BF2",
    x"18A994B",
    x"18A96A5",
    x"18A9400",
    x"18A915B",
    x"18A8EB7",
    x"18A8C14",
    x"18A8971",
    x"18A86CF",
    x"18A842E",
    x"18A818D",
    x"18A7EED",
    x"18A7C4E",
    x"18A79AF",
    x"18A7711",
    x"18A7473",
    x"18A71D7",
    x"18A6F3A",
    x"18A6C9F",
    x"18A6A04",
    x"18A676A",
    x"18A64D0",
    x"18A6238",
    x"18A5F9F",
    x"18A5D08",
    x"18A5A71",
    x"18A57DB",
    x"18A5545",
    x"18A52B0",
    x"18A501C",
    x"18A4D88",
    x"18A4AF5",
    x"18A4862",
    x"18A45D1",
    x"18A433F",
    x"18A40AF",
    x"18A3E1F",
    x"18A3B90",
    x"18A3901",
    x"18A3673",
    x"18A33E6",
    x"18A3159",
    x"18A2ECD",
    x"18A2C42",
    x"18A29B7",
    x"18A272D",
    x"18A24A4",
    x"18A221B",
    x"18A1F93",
    x"18A1D0B",
    x"18A1A84",
    x"18A17FE",
    x"18A1578",
    x"18A12F3",
    x"18A106F",
    x"18A0DEB",
    x"18A0B68",
    x"18A08E5",
    x"18A0663",
    x"18A03E2",
    x"18A0161",
    x"189FEE1",
    x"189FC62",
    x"189F9E3",
    x"189F765",
    x"189F4E7",
    x"189F26A",
    x"189EFEE",
    x"189ED72",
    x"189EAF7",
    x"189E87D",
    x"189E603",
    x"189E38A",
    x"189E111",
    x"189DE99",
    x"189DC22",
    x"189D9AB",
    x"189D735",
    x"189D4C0",
    x"189D24B",
    x"189CFD7",
    x"189CD63",
    x"189CAF0",
    x"189C87E",
    x"189C60C",
    x"189C39A",
    x"189C12A",
    x"189BEBA",
    x"189BC4B",
    x"189B9DC",
    x"189B76E",
    x"189B500",
    x"189B293",
    x"189B027",
    x"189ADBB",
    x"189AB50",
    x"189A8E5",
    x"189A67B",
    x"189A412",
    x"189A1A9",
    x"1899F41",
    x"1899CDA",
    x"1899A73",
    x"189980D",
    x"18995A7",
    x"1899342",
    x"18990DD",
    x"1898E79",
    x"1898C16",
    x"18989B3",
    x"1898751",
    x"18984F0",
    x"189828F",
    x"189802E",
    x"1897DCF",
    x"1897B6F",
    x"1897911",
    x"18976B3",
    x"1897455",
    x"18971F9",
    x"1896F9D",
    x"1896D41",
    x"1896AE6",
    x"189688B",
    x"1896632",
    x"18963D8",
    x"1896180",
    x"1895F28",
    x"1895CD0",
    x"1895A79",
    x"1895823",
    x"18955CD",
    x"1895378",
    x"1895123",
    x"1894ECF",
    x"1894C7C",
    x"1894A29",
    x"18947D7",
    x"1894585",
    x"1894334",
    x"18940E4",
    x"1893E94",
    x"1893C44",
    x"18939F6",
    x"18937A7",
    x"189355A",
    x"189330D",
    x"18930C0",
    x"1892E74",
    x"1892C29",
    x"18929DE",
    x"1892794",
    x"189254A",
    x"1892301",
    x"18920B9",
    x"1891E71",
    x"1891C2A",
    x"18919E3",
    x"189179D",
    x"1891557",
    x"1891312",
    x"18910CE",
    x"1890E8A",
    x"1890C46",
    x"1890A04",
    x"18907C1",
    x"1890580",
    x"189033F",
    x"18900FE",
    x"188FEBE",
    x"188FC7F",
    x"188FA40",
    x"188F802",
    x"188F5C4",
    x"188F387",
    x"188F14A",
    x"188EF0E",
    x"188ECD3",
    x"188EA98",
    x"188E85D",
    x"188E623",
    x"188E3EA",
    x"188E1B1",
    x"188DF79",
    x"188DD42",
    x"188DB0B",
    x"188D8D4",
    x"188D69E",
    x"188D469",
    x"188D234",
    x"188D000",
    x"188CDCC",
    x"188CB99",
    x"188C966",
    x"188C734",
    x"188C503",
    x"188C2D2",
    x"188C0A1",
    x"188BE71",
    x"188BC42",
    x"188BA13",
    x"188B7E5",
    x"188B5B7",
    x"188B38A",
    x"188B15E",
    x"188AF31",
    x"188AD06",
    x"188AADB",
    x"188A8B0",
    x"188A687",
    x"188A45D",
    x"188A234",
    x"188A00C",
    x"1889DE4",
    x"1889BBD",
    x"1889997",
    x"1889770",
    x"188954B",
    x"1889326",
    x"1889101",
    x"1888EDD",
    x"1888CBA",
    x"1888A97",
    x"1888874",
    x"1888653",
    x"1888431",
    x"1888211",
    x"1887FF0",
    x"1887DD1",
    x"1887BB1",
    x"1887993",
    x"1887775",
    x"1887557",
    x"188733A",
    x"188711D",
    x"1886F01",
    x"1886CE6",
    x"1886ACB",
    x"18868B0",
    x"1886697",
    x"188647D",
    x"1886264",
    x"188604C",
    x"1885E34",
    x"1885C1D",
    x"1885A06",
    x"18857F0",
    x"18855DA",
    x"18853C5",
    x"18851B0",
    x"1884F9C",
    x"1884D88",
    x"1884B75",
    x"1884963",
    x"1884751",
    x"188453F",
    x"188432E",
    x"188411D",
    x"1883F0D",
    x"1883CFE",
    x"1883AEF",
    x"18838E0",
    x"18836D3",
    x"18834C5",
    x"18832B8",
    x"18830AC",
    x"1882EA0",
    x"1882C94",
    x"1882A8A",
    x"188287F",
    x"1882675",
    x"188246C",
    x"1882263",
    x"188205B",
    x"1881E53",
    x"1881C4C",
    x"1881A45",
    x"188183E",
    x"1881639",
    x"1881433",
    x"188122E",
    x"188102A",
    x"1880E26",
    x"1880C23",
    x"1880A20",
    x"188081E",
    x"188061C",
    x"188041B",
    x"188021A",
    x"188001A",
    x"187FC35",
    x"187F836",
    x"187F439",
    x"187F03C",
    x"187EC41",
    x"187E846",
    x"187E44C",
    x"187E054",
    x"187DC5C",
    x"187D866",
    x"187D470",
    x"187D07B",
    x"187CC88",
    x"187C895",
    x"187C4A4",
    x"187C0B3",
    x"187BCC3",
    x"187B8D5",
    x"187B4E7",
    x"187B0FA",
    x"187AD0E",
    x"187A924",
    x"187A53A",
    x"187A151",
    x"1879D69",
    x"1879982",
    x"187959C",
    x"18791B7",
    x"1878DD3",
    x"18789F0",
    x"187860E",
    x"187822D",
    x"1877E4D",
    x"1877A6E",
    x"1877690",
    x"18772B3",
    x"1876ED7",
    x"1876AFC",
    x"1876721",
    x"1876348",
    x"1875F70",
    x"1875B98",
    x"18757C2",
    x"18753EC",
    x"1875018",
    x"1874C44",
    x"1874872",
    x"18744A0",
    x"18740CF",
    x"1873D00",
    x"1873931",
    x"1873563",
    x"1873196",
    x"1872DCA",
    x"18729FF",
    x"1872635",
    x"187226C",
    x"1871EA4",
    x"1871ADD",
    x"1871717",
    x"1871351",
    x"1870F8D",
    x"1870BCA",
    x"1870807",
    x"1870446",
    x"1870085",
    x"186FCC5",
    x"186F907",
    x"186F549",
    x"186F18C",
    x"186EDD0",
    x"186EA15",
    x"186E65B",
    x"186E2A2",
    x"186DEEA",
    x"186DB32",
    x"186D77C",
    x"186D3C7",
    x"186D012",
    x"186CC5F",
    x"186C8AC",
    x"186C4FA",
    x"186C14A",
    x"186BD9A",
    x"186B9EB",
    x"186B63D",
    x"186B290",
    x"186AEE3",
    x"186AB38",
    x"186A78E",
    x"186A3E4",
    x"186A03C",
    x"1869C94",
    x"18698EE",
    x"1869548",
    x"18691A3",
    x"1868DFF",
    x"1868A5C",
    x"18686BA",
    x"1868319",
    x"1867F78",
    x"1867BD9",
    x"186783A",
    x"186749D",
    x"1867100",
    x"1866D64",
    x"18669C9",
    x"186662F",
    x"1866296",
    x"1865EFE",
    x"1865B67",
    x"18657D0",
    x"186543B",
    x"18650A6",
    x"1864D13",
    x"1864980",
    x"18645EE",
    x"186425D",
    x"1863ECD",
    x"1863B3D",
    x"18637AF",
    x"1863421",
    x"1863095",
    x"1862D09",
    x"186297E",
    x"18625F4",
    x"186226B",
    x"1861EE3",
    x"1861B5C",
    x"18617D6",
    x"1861450",
    x"18610CB",
    x"1860D48",
    x"18609C5",
    x"1860643",
    x"18602C2",
    x"185FF41",
    x"185FBC2",
    x"185F843",
    x"185F4C6",
    x"185F149",
    x"185EDCD",
    x"185EA52",
    x"185E6D8",
    x"185E35F",
    x"185DFE6",
    x"185DC6F",
    x"185D8F8",
    x"185D582",
    x"185D20D",
    x"185CE99",
    x"185CB26",
    x"185C7B4",
    x"185C442",
    x"185C0D2",
    x"185BD62",
    x"185B9F3",
    x"185B685",
    x"185B318",
    x"185AFAB",
    x"185AC40",
    x"185A8D5",
    x"185A56B",
    x"185A202",
    x"1859E9A",
    x"1859B33",
    x"18597CD",
    x"1859467",
    x"1859103",
    x"1858D9F",
    x"1858A3C",
    x"18586DA",
    x"1858378",
    x"1858018",
    x"1857CB8",
    x"185795A",
    x"18575FC",
    x"185729F",
    x"1856F42",
    x"1856BE7",
    x"185688C",
    x"1856533",
    x"18561DA",
    x"1855E82",
    x"1855B2B",
    x"18557D4",
    x"185547F",
    x"185512A",
    x"1854DD6",
    x"1854A83",
    x"1854731",
    x"18543DF",
    x"185408F",
    x"1853D3F",
    x"18539F0",
    x"18536A2",
    x"1853355",
    x"1853008",
    x"1852CBD",
    x"1852972",
    x"1852628",
    x"18522DF",
    x"1851F97",
    x"1851C4F",
    x"1851909",
    x"18515C3",
    x"185127E",
    x"1850F39",
    x"1850BF6",
    x"18508B3",
    x"1850572",
    x"1850231",
    x"184FEF1",
    x"184FBB1",
    x"184F873",
    x"184F535",
    x"184F1F8",
    x"184EEBC",
    x"184EB81",
    x"184E846",
    x"184E50D",
    x"184E1D4",
    x"184DE9C",
    x"184DB64",
    x"184D82E",
    x"184D4F8",
    x"184D1C4",
    x"184CE90",
    x"184CB5C",
    x"184C82A",
    x"184C4F8",
    x"184C1C7",
    x"184BE97",
    x"184BB68",
    x"184B83A",
    x"184B50C",
    x"184B1DF",
    x"184AEB3",
    x"184AB88",
    x"184A85D",
    x"184A534",
    x"184A20B",
    x"1849EE3",
    x"1849BBB",
    x"1849895",
    x"184956F",
    x"184924A",
    x"1848F26",
    x"1848C02",
    x"18488E0",
    x"18485BE",
    x"184829D",
    x"1847F7D",
    x"1847C5D",
    x"184793E",
    x"1847620",
    x"1847303",
    x"1846FE7",
    x"1846CCB",
    x"18469B1",
    x"1846697",
    x"184637D",
    x"1846065",
    x"1845D4D",
    x"1845A36",
    x"1845720",
    x"184540B",
    x"18450F6",
    x"1844DE2",
    x"1844ACF",
    x"18447BD",
    x"18444AB",
    x"184419A",
    x"1843E8A",
    x"1843B7B",
    x"184386D",
    x"184355F",
    x"1843252",
    x"1842F46",
    x"1842C3A",
    x"1842930",
    x"1842626",
    x"184231D",
    x"1842014",
    x"1841D0C",
    x"1841A06",
    x"18416FF",
    x"18413FA",
    x"18410F5",
    x"1840DF2",
    x"1840AEF",
    x"18407EC",
    x"18404EB",
    x"18401EA",
    x"183FEEA",
    x"183FBEA",
    x"183F8EC",
    x"183F5EE",
    x"183F2F1",
    x"183EFF4",
    x"183ECF9",
    x"183E9FE",
    x"183E704",
    x"183E40A",
    x"183E112",
    x"183DE1A",
    x"183DB23",
    x"183D82C",
    x"183D537",
    x"183D242",
    x"183CF4D",
    x"183CC5A",
    x"183C967",
    x"183C675",
    x"183C384",
    x"183C093",
    x"183BDA4",
    x"183BAB5",
    x"183B7C6",
    x"183B4D9",
    x"183B1EC",
    x"183AF00",
    x"183AC14",
    x"183A92A",
    x"183A640",
    x"183A357",
    x"183A06E",
    x"1839D86",
    x"1839A9F",
    x"18397B9",
    x"18394D4",
    x"18391EF",
    x"1838F0B",
    x"1838C27",
    x"1838945",
    x"1838663",
    x"1838381",
    x"18380A1",
    x"1837DC1",
    x"1837AE2",
    x"1837804",
    x"1837526",
    x"1837249",
    x"1836F6D",
    x"1836C91",
    x"18369B6",
    x"18366DC",
    x"1836403",
    x"183612A",
    x"1835E52",
    x"1835B7B",
    x"18358A5",
    x"18355CF",
    x"18352FA",
    x"1835025",
    x"1834D52",
    x"1834A7F",
    x"18347AD",
    x"18344DB",
    x"183420A",
    x"1833F3A",
    x"1833C6A",
    x"183399C",
    x"18336CE",
    x"1833400",
    x"1833134",
    x"1832E68",
    x"1832B9C",
    x"18328D2",
    x"1832608",
    x"183233F",
    x"1832076",
    x"1831DAF",
    x"1831AE8",
    x"1831821",
    x"183155C",
    x"1831297",
    x"1830FD2",
    x"1830D0F",
    x"1830A4C",
    x"1830789",
    x"18304C8",
    x"1830207",
    x"182FF47",
    x"182FC87",
    x"182F9C9",
    x"182F70B",
    x"182F44D",
    x"182F190",
    x"182EED4",
    x"182EC19",
    x"182E95E",
    x"182E6A4",
    x"182E3EB",
    x"182E132",
    x"182DE7A",
    x"182DBC3",
    x"182D90C",
    x"182D657",
    x"182D3A1",
    x"182D0ED",
    x"182CE39",
    x"182CB86",
    x"182C8D3",
    x"182C621",
    x"182C370",
    x"182C0BF",
    x"182BE10",
    x"182BB60",
    x"182B8B2",
    x"182B604",
    x"182B357",
    x"182B0AA",
    x"182ADFF",
    x"182AB53",
    x"182A8A9",
    x"182A5FF",
    x"182A356",
    x"182A0AD",
    x"1829E06",
    x"1829B5E",
    x"18298B8",
    x"1829612",
    x"182936D",
    x"18290C8",
    x"1828E24",
    x"1828B81",
    x"18288DF",
    x"182863D",
    x"182839C",
    x"18280FB",
    x"1827E5B",
    x"1827BBC",
    x"182791D",
    x"182767F",
    x"18273E2",
    x"1827145",
    x"1826EA9",
    x"1826C0E",
    x"1826973",
    x"18266D9",
    x"1826440",
    x"18261A7",
    x"1825F0F",
    x"1825C78",
    x"18259E1",
    x"182574B",
    x"18254B5",
    x"1825220",
    x"1824F8C",
    x"1824CF9",
    x"1824A66",
    x"18247D3",
    x"1824542",
    x"18242B1",
    x"1824020",
    x"1823D91",
    x"1823B02",
    x"1823873",
    x"18235E5",
    x"1823358",
    x"18230CC",
    x"1822E40",
    x"1822BB5",
    x"182292A",
    x"18226A0",
    x"1822417",
    x"182218E",
    x"1821F06",
    x"1821C7E",
    x"18219F8",
    x"1821771",
    x"18214EC",
    x"1821267",
    x"1820FE3",
    x"1820D5F",
    x"1820ADC",
    x"182085A",
    x"18205D8",
    x"1820357",
    x"18200D6",
    x"181FE56",
    x"181FBD7",
    x"181F958",
    x"181F6DA",
    x"181F45D",
    x"181F1E0",
    x"181EF64",
    x"181ECE8",
    x"181EA6E",
    x"181E7F3",
    x"181E57A",
    x"181E300",
    x"181E088",
    x"181DE10",
    x"181DB99",
    x"181D922",
    x"181D6AC",
    x"181D437",
    x"181D1C2",
    x"181CF4E",
    x"181CCDB",
    x"181CA68",
    x"181C7F5",
    x"181C584",
    x"181C313",
    x"181C0A2",
    x"181BE32",
    x"181BBC3",
    x"181B955",
    x"181B6E6",
    x"181B479",
    x"181B20C",
    x"181AFA0",
    x"181AD34",
    x"181AAC9",
    x"181A85F",
    x"181A5F5",
    x"181A38C",
    x"181A123",
    x"1819EBC",
    x"1819C54",
    x"18199ED",
    x"1819787",
    x"1819522",
    x"18192BD",
    x"1819058",
    x"1818DF4",
    x"1818B91",
    x"181892F",
    x"18186CD",
    x"181846B",
    x"181820A",
    x"1817FAA",
    x"1817D4B",
    x"1817AEC",
    x"181788D",
    x"181762F",
    x"18173D2",
    x"1817175",
    x"1816F19",
    x"1816CBE",
    x"1816A63",
    x"1816809",
    x"18165AF",
    x"1816356",
    x"18160FD",
    x"1815EA5",
    x"1815C4E",
    x"18159F7",
    x"18157A1",
    x"181554B",
    x"18152F6",
    x"18150A2",
    x"1814E4E",
    x"1814BFB",
    x"18149A8",
    x"1814756",
    x"1814504",
    x"18142B3",
    x"1814063",
    x"1813E13",
    x"1813BC4",
    x"1813975",
    x"1813727",
    x"18134DA",
    x"181328D",
    x"1813040",
    x"1812DF5",
    x"1812BA9",
    x"181295F",
    x"1812715",
    x"18124CB",
    x"1812282",
    x"181203A",
    x"1811DF2",
    x"1811BAB",
    x"1811964",
    x"181171E",
    x"18114D9",
    x"1811294",
    x"1811050",
    x"1810E0C",
    x"1810BC9",
    x"1810986",
    x"1810744",
    x"1810502",
    x"18102C1",
    x"1810081",
    x"180FE41",
    x"180FC02",
    x"180F9C3",
    x"180F785",
    x"180F547",
    x"180F30A",
    x"180F0CE",
    x"180EE92",
    x"180EC56",
    x"180EA1C",
    x"180E7E1",
    x"180E5A8",
    x"180E36F",
    x"180E136",
    x"180DEFE",
    x"180DCC6",
    x"180DA90",
    x"180D859",
    x"180D623",
    x"180D3EE",
    x"180D1B9",
    x"180CF85",
    x"180CD52",
    x"180CB1F",
    x"180C8EC",
    x"180C6BA",
    x"180C489",
    x"180C258",
    x"180C028",
    x"180BDF8",
    x"180BBC9",
    x"180B99A",
    x"180B76C",
    x"180B53E",
    x"180B311",
    x"180B0E5",
    x"180AEB9",
    x"180AC8D",
    x"180AA62",
    x"180A838",
    x"180A60E",
    x"180A3E5",
    x"180A1BC",
    x"1809F94",
    x"1809D6D",
    x"1809B45",
    x"180991F",
    x"18096F9",
    x"18094D3",
    x"18092AF",
    x"180908A",
    x"1808E66",
    x"1808C43",
    x"1808A20",
    x"18087FE",
    x"18085DC",
    x"18083BB",
    x"180819A",
    x"1807F7A",
    x"1807D5B",
    x"1807B3B",
    x"180791D",
    x"18076FF",
    x"18074E1",
    x"18072C4",
    x"18070A8",
    x"1806E8C",
    x"1806C71",
    x"1806A56",
    x"180683C",
    x"1806622",
    x"1806408",
    x"18061F0",
    x"1805FD8",
    x"1805DC0",
    x"1805BA9",
    x"1805992",
    x"180577C",
    x"1805566",
    x"1805351",
    x"180513D",
    x"1804F29",
    x"1804D15",
    x"1804B02",
    x"18048F0",
    x"18046DE",
    x"18044CC",
    x"18042BB",
    x"18040AB",
    x"1803E9B",
    x"1803C8B",
    x"1803A7D",
    x"180386E",
    x"1803660",
    x"1803453",
    x"1803246",
    x"180303A",
    x"1802E2E",
    x"1802C23",
    x"1802A18",
    x"180280E",
    x"1802604",
    x"18023FB",
    x"18021F2",
    x"1801FEA",
    x"1801DE2",
    x"1801BDB",
    x"18019D4",
    x"18017CE",
    x"18015C8",
    x"18013C3",
    x"18011BE",
    x"1800FBA",
    x"1800DB6",
    x"1800BB3",
    x"18009B1",
    x"18007AE",
    x"18005AD",
    x"18003AC",
    x"18001AB",
    x"17FFF56",
    x"17FFB57",
    x"17FF758",
    x"17FF35B",
    x"17FEF5F",
    x"17FEB63",
    x"17FE769",
    x"17FE36F",
    x"17FDF77",
    x"17FDB80",
    x"17FD789",
    x"17FD394",
    x"17FCFA0",
    x"17FCBAC",
    x"17FC7BA",
    x"17FC3C8",
    x"17FBFD8",
    x"17FBBE8",
    x"17FB7FA",
    x"17FB40C",
    x"17FB020",
    x"17FAC34",
    x"17FA84A",
    x"17FA460",
    x"17FA078",
    x"17F9C90",
    x"17F98A9",
    x"17F94C4",
    x"17F90DF",
    x"17F8CFB",
    x"17F8918",
    x"17F8537",
    x"17F8156",
    x"17F7D76",
    x"17F7997",
    x"17F75B9",
    x"17F71DC",
    x"17F6E00",
    x"17F6A25",
    x"17F664B",
    x"17F6272",
    x"17F5E9A",
    x"17F5AC3",
    x"17F56ED",
    x"17F5317",
    x"17F4F43",
    x"17F4B70",
    x"17F479D",
    x"17F43CC",
    x"17F3FFB",
    x"17F3C2C",
    x"17F385D",
    x"17F3490",
    x"17F30C3",
    x"17F2CF7",
    x"17F292D",
    x"17F2563",
    x"17F219A",
    x"17F1DD2",
    x"17F1A0B",
    x"17F1645",
    x"17F1280",
    x"17F0EBC",
    x"17F0AF8",
    x"17F0736",
    x"17F0375",
    x"17EFFB4",
    x"17EFBF5",
    x"17EF836",
    x"17EF479",
    x"17EF0BC",
    x"17EED00",
    x"17EE946",
    x"17EE58C",
    x"17EE1D3",
    x"17EDE1B",
    x"17EDA64",
    x"17ED6AE",
    x"17ED2F9",
    x"17ECF44",
    x"17ECB91",
    x"17EC7DE",
    x"17EC42D",
    x"17EC07C",
    x"17EBCCD",
    x"17EB91E",
    x"17EB570",
    x"17EB1C3",
    x"17EAE17",
    x"17EAA6C",
    x"17EA6C2",
    x"17EA319",
    x"17E9F71",
    x"17E9BC9",
    x"17E9823",
    x"17E947D",
    x"17E90D8",
    x"17E8D35",
    x"17E8992",
    x"17E85F0",
    x"17E824F",
    x"17E7EAF",
    x"17E7B0F",
    x"17E7771",
    x"17E73D4",
    x"17E7037",
    x"17E6C9C",
    x"17E6901",
    x"17E6567",
    x"17E61CE",
    x"17E5E36",
    x"17E5A9F",
    x"17E5709",
    x"17E5374",
    x"17E4FDF",
    x"17E4C4C",
    x"17E48B9",
    x"17E4527",
    x"17E4196",
    x"17E3E07",
    x"17E3A77",
    x"17E36E9",
    x"17E335C",
    x"17E2FD0",
    x"17E2C44",
    x"17E28B9",
    x"17E2530",
    x"17E21A7",
    x"17E1E1F",
    x"17E1A98",
    x"17E1712",
    x"17E138C",
    x"17E1008",
    x"17E0C84",
    x"17E0902",
    x"17E0580",
    x"17E01FF",
    x"17DFE7F",
    x"17DFB00",
    x"17DF781",
    x"17DF404",
    x"17DF087",
    x"17DED0C",
    x"17DE991",
    x"17DE617",
    x"17DE29E",
    x"17DDF25",
    x"17DDBAE",
    x"17DD838",
    x"17DD4C2",
    x"17DD14D",
    x"17DCDD9",
    x"17DCA66",
    x"17DC6F4",
    x"17DC383",
    x"17DC012",
    x"17DBCA3",
    x"17DB934",
    x"17DB5C6",
    x"17DB259",
    x"17DAEED",
    x"17DAB82",
    x"17DA817",
    x"17DA4AE",
    x"17DA145",
    x"17D9DDD",
    x"17D9A76",
    x"17D9710",
    x"17D93AA",
    x"17D9046",
    x"17D8CE2",
    x"17D8980",
    x"17D861E",
    x"17D82BC",
    x"17D7F5C",
    x"17D7BFD",
    x"17D789E",
    x"17D7540",
    x"17D71E4",
    x"17D6E88",
    x"17D6B2C",
    x"17D67D2",
    x"17D6478",
    x"17D6120",
    x"17D5DC8",
    x"17D5A71",
    x"17D571B",
    x"17D53C5",
    x"17D5071",
    x"17D4D1D",
    x"17D49CA",
    x"17D4678",
    x"17D4327",
    x"17D3FD7",
    x"17D3C87",
    x"17D3938",
    x"17D35EA",
    x"17D329D",
    x"17D2F51",
    x"17D2C06",
    x"17D28BB",
    x"17D2571",
    x"17D2228",
    x"17D1EE0",
    x"17D1B99",
    x"17D1852",
    x"17D150D",
    x"17D11C8",
    x"17D0E84",
    x"17D0B41",
    x"17D07FE",
    x"17D04BD",
    x"17D017C",
    x"17CFE3C",
    x"17CFAFD",
    x"17CF7BE",
    x"17CF481",
    x"17CF144",
    x"17CEE08",
    x"17CEACD",
    x"17CE793",
    x"17CE459",
    x"17CE121",
    x"17CDDE9",
    x"17CDAB2",
    x"17CD77B",
    x"17CD446",
    x"17CD111",
    x"17CCDDD",
    x"17CCAAA",
    x"17CC778",
    x"17CC447",
    x"17CC116",
    x"17CBDE6",
    x"17CBAB7",
    x"17CB789",
    x"17CB45B",
    x"17CB12F",
    x"17CAE03",
    x"17CAAD8",
    x"17CA7AD",
    x"17CA484",
    x"17CA15B",
    x"17C9E33",
    x"17C9B0C",
    x"17C97E5",
    x"17C94C0",
    x"17C919B",
    x"17C8E77",
    x"17C8B54",
    x"17C8831",
    x"17C8510",
    x"17C81EF",
    x"17C7ECF",
    x"17C7BB0",
    x"17C7891",
    x"17C7573",
    x"17C7256",
    x"17C6F3A",
    x"17C6C1F",
    x"17C6904",
    x"17C65EA",
    x"17C62D1",
    x"17C5FB9",
    x"17C5CA1",
    x"17C598A",
    x"17C5674",
    x"17C535F",
    x"17C504B",
    x"17C4D37",
    x"17C4A24",
    x"17C4712",
    x"17C4401",
    x"17C40F0",
    x"17C3DE0",
    x"17C3AD1",
    x"17C37C3",
    x"17C34B5",
    x"17C31A8",
    x"17C2E9C",
    x"17C2B91",
    x"17C2887",
    x"17C257D",
    x"17C2274",
    x"17C1F6C",
    x"17C1C64",
    x"17C195D",
    x"17C1657",
    x"17C1352",
    x"17C104E",
    x"17C0D4A",
    x"17C0A47",
    x"17C0745",
    x"17C0443",
    x"17C0143",
    x"17BFE43",
    x"17BFB44",
    x"17BF845",
    x"17BF547",
    x"17BF24B",
    x"17BEF4E",
    x"17BEC53",
    x"17BE958",
    x"17BE65E",
    x"17BE365",
    x"17BE06D",
    x"17BDD75",
    x"17BDA7E",
    x"17BD788",
    x"17BD492",
    x"17BD19D",
    x"17BCEA9",
    x"17BCBB6",
    x"17BC8C3",
    x"17BC5D2",
    x"17BC2E0",
    x"17BBFF0",
    x"17BBD00",
    x"17BBA12",
    x"17BB723",
    x"17BB436",
    x"17BB149",
    x"17BAE5D",
    x"17BAB72",
    x"17BA888",
    x"17BA59E",
    x"17BA2B5",
    x"17B9FCD",
    x"17B9CE5",
    x"17B99FE",
    x"17B9718",
    x"17B9433",
    x"17B914E",
    x"17B8E6A",
    x"17B8B87",
    x"17B88A4",
    x"17B85C2",
    x"17B82E1",
    x"17B8001",
    x"17B7D21",
    x"17B7A42",
    x"17B7764",
    x"17B7487",
    x"17B71AA",
    x"17B6ECE",
    x"17B6BF2",
    x"17B6918",
    x"17B663E",
    x"17B6365",
    x"17B608C",
    x"17B5DB4",
    x"17B5ADD",
    x"17B5807",
    x"17B5531",
    x"17B525C",
    x"17B4F88",
    x"17B4CB5",
    x"17B49E2",
    x"17B4710",
    x"17B443E",
    x"17B416E",
    x"17B3E9E",
    x"17B3BCE",
    x"17B3900",
    x"17B3632",
    x"17B3365",
    x"17B3098",
    x"17B2DCC",
    x"17B2B01",
    x"17B2837",
    x"17B256D",
    x"17B22A4",
    x"17B1FDC",
    x"17B1D14",
    x"17B1A4D",
    x"17B1787",
    x"17B14C1",
    x"17B11FD",
    x"17B0F38",
    x"17B0C75",
    x"17B09B2",
    x"17B06F0",
    x"17B042F",
    x"17B016E",
    x"17AFEAE",
    x"17AFBEF",
    x"17AF930",
    x"17AF672",
    x"17AF3B5",
    x"17AF0F8",
    x"17AEE3C",
    x"17AEB81",
    x"17AE8C7",
    x"17AE60D",
    x"17AE354",
    x"17AE09B",
    x"17ADDE3",
    x"17ADB2C",
    x"17AD876",
    x"17AD5C0",
    x"17AD30B",
    x"17AD056",
    x"17ACDA3",
    x"17ACAF0",
    x"17AC83D",
    x"17AC58B",
    x"17AC2DA",
    x"17AC02A",
    x"17ABD7A",
    x"17ABACB",
    x"17AB81D",
    x"17AB56F",
    x"17AB2C2",
    x"17AB016",
    x"17AAD6A",
    x"17AAABF",
    x"17AA815",
    x"17AA56B",
    x"17AA2C2",
    x"17AA01A",
    x"17A9D72",
    x"17A9ACB",
    x"17A9825",
    x"17A957F",
    x"17A92DA",
    x"17A9035",
    x"17A8D92",
    x"17A8AEF",
    x"17A884C",
    x"17A85AB",
    x"17A8309",
    x"17A8069",
    x"17A7DC9",
    x"17A7B2A",
    x"17A788C",
    x"17A75EE",
    x"17A7351",
    x"17A70B4",
    x"17A6E18",
    x"17A6B7D",
    x"17A68E3",
    x"17A6649",
    x"17A63AF",
    x"17A6117",
    x"17A5E7F",
    x"17A5BE8",
    x"17A5951",
    x"17A56BB",
    x"17A5426",
    x"17A5191",
    x"17A4EFD",
    x"17A4C69",
    x"17A49D7",
    x"17A4744",
    x"17A44B3",
    x"17A4222",
    x"17A3F92",
    x"17A3D02",
    x"17A3A73",
    x"17A37E5",
    x"17A3557",
    x"17A32CA",
    x"17A303E",
    x"17A2DB2",
    x"17A2B27",
    x"17A289D",
    x"17A2613",
    x"17A238A",
    x"17A2101",
    x"17A1E79",
    x"17A1BF2",
    x"17A196B",
    x"17A16E5",
    x"17A1460",
    x"17A11DB",
    x"17A0F57",
    x"17A0CD3",
    x"17A0A50",
    x"17A07CE",
    x"17A054C",
    x"17A02CB",
    x"17A004B",
    x"179FDCB",
    x"179FB4C",
    x"179F8CE",
    x"179F650",
    x"179F3D3",
    x"179F156",
    x"179EEDA",
    x"179EC5E",
    x"179E9E4",
    x"179E769",
    x"179E4F0",
    x"179E277",
    x"179DFFF",
    x"179DD87",
    x"179DB10",
    x"179D899",
    x"179D624",
    x"179D3AE",
    x"179D13A",
    x"179CEC6",
    x"179CC52",
    x"179C9E0",
    x"179C76D",
    x"179C4FC",
    x"179C28B",
    x"179C01B",
    x"179BDAB",
    x"179BB3C",
    x"179B8CD",
    x"179B65F",
    x"179B3F2",
    x"179B185",
    x"179AF19",
    x"179ACAE",
    x"179AA43",
    x"179A7D9",
    x"179A56F",
    x"179A306",
    x"179A09E",
    x"1799E36",
    x"1799BCE",
    x"1799968",
    x"1799702",
    x"179949C",
    x"1799237",
    x"1798FD3",
    x"1798D70",
    x"1798B0C",
    x"17988AA",
    x"1798648",
    x"17983E7",
    x"1798186",
    x"1797F26",
    x"1797CC7",
    x"1797A68",
    x"1797809",
    x"17975AC",
    x"179734F",
    x"17970F2",
    x"1796E96",
    x"1796C3B",
    x"17969E0",
    x"1796786",
    x"179652C",
    x"17962D3",
    x"179607B",
    x"1795E23",
    x"1795BCC",
    x"1795975",
    x"179571F",
    x"17954CA",
    x"1795275",
    x"1795020",
    x"1794DCD",
    x"1794B79",
    x"1794927",
    x"17946D5",
    x"1794483",
    x"1794233",
    x"1793FE2",
    x"1793D93",
    x"1793B44",
    x"17938F5",
    x"17936A7",
    x"179345A",
    x"179320D",
    x"1792FC1",
    x"1792D75",
    x"1792B2A",
    x"17928DF",
    x"1792695",
    x"179244C",
    x"1792203",
    x"1791FBB",
    x"1791D73",
    x"1791B2C",
    x"17918E6",
    x"17916A0",
    x"179145B",
    x"1791216",
    x"1790FD2",
    x"1790D8E",
    x"1790B4B",
    x"1790908",
    x"17906C6",
    x"1790485",
    x"1790244",
    x"1790004",
    x"178FDC4",
    x"178FB85",
    x"178F946",
    x"178F708",
    x"178F4CB",
    x"178F28E",
    x"178F051",
    x"178EE16",
    x"178EBDA",
    x"178E9A0",
    x"178E766",
    x"178E52C",
    x"178E2F3",
    x"178E0BA",
    x"178DE83",
    x"178DC4B",
    x"178DA14",
    x"178D7DE",
    x"178D5A9",
    x"178D373",
    x"178D13F",
    x"178CF0B",
    x"178CCD7",
    x"178CAA4",
    x"178C872",
    x"178C640",
    x"178C40F",
    x"178C1DE",
    x"178BFAE",
    x"178BD7E",
    x"178BB4F",
    x"178B921",
    x"178B6F3",
    x"178B4C5",
    x"178B298",
    x"178B06C",
    x"178AE40",
    x"178AC15",
    x"178A9EA",
    x"178A7C0",
    x"178A596",
    x"178A36D",
    x"178A144",
    x"1789F1C",
    x"1789CF5",
    x"1789ACE",
    x"17898A7",
    x"1789681",
    x"178945C",
    x"1789237",
    x"1789013",
    x"1788DEF",
    x"1788BCC",
    x"17889A9",
    x"1788787",
    x"1788566",
    x"1788345",
    x"1788124",
    x"1787F04",
    x"1787CE4",
    x"1787AC5",
    x"17878A7",
    x"1787689",
    x"178746C",
    x"178724F",
    x"1787033",
    x"1786E17",
    x"1786BFC",
    x"17869E1",
    x"17867C7",
    x"17865AD",
    x"1786394",
    x"178617B",
    x"1785F63",
    x"1785D4B",
    x"1785B34",
    x"178591E",
    x"1785708",
    x"17854F2",
    x"17852DD",
    x"17850C9",
    x"1784EB5",
    x"1784CA2",
    x"1784A8F",
    x"178487C",
    x"178466A",
    x"1784459",
    x"1784248",
    x"1784038",
    x"1783E28",
    x"1783C19",
    x"1783A0A",
    x"17837FC",
    x"17835EE",
    x"17833E1",
    x"17831D4",
    x"1782FC8",
    x"1782DBC",
    x"1782BB1",
    x"17829A6",
    x"178279C",
    x"1782593",
    x"1782389",
    x"1782181",
    x"1781F79",
    x"1781D71",
    x"1781B6A",
    x"1781963",
    x"178175D",
    x"1781558",
    x"1781353",
    x"178114E",
    x"1780F4A",
    x"1780D46",
    x"1780B43",
    x"1780941",
    x"178073F",
    x"178053D",
    x"178033C",
    x"178013C",
    x"177FE77",
    x"177FA78",
    x"177F67A",
    x"177F27D",
    x"177EE81",
    x"177EA86",
    x"177E68C",
    x"177E293",
    x"177DE9A",
    x"177DAA3",
    x"177D6AD",
    x"177D2B8",
    x"177CEC4",
    x"177CAD1",
    x"177C6DE",
    x"177C2ED",
    x"177BEFD",
    x"177BB0E",
    x"177B71F",
    x"177B332",
    x"177AF46",
    x"177AB5A",
    x"177A770",
    x"177A387",
    x"1779F9E",
    x"1779BB7",
    x"17797D0",
    x"17793EB",
    x"1779006",
    x"1778C23",
    x"1778840",
    x"177845F",
    x"177807E",
    x"1777C9F",
    x"17778C0",
    x"17774E2",
    x"1777105",
    x"1776D2A",
    x"177694F",
    x"1776575",
    x"177619C",
    x"1775DC4",
    x"17759ED",
    x"1775617",
    x"1775242",
    x"1774E6E",
    x"1774A9B",
    x"17746C9",
    x"17742F8",
    x"1773F27",
    x"1773B58",
    x"177378A",
    x"17733BC",
    x"1772FF0",
    x"1772C24",
    x"177285A",
    x"1772490",
    x"17720C7",
    x"1771D00",
    x"1771939",
    x"1771573",
    x"17711AE",
    x"1770DEA",
    x"1770A27",
    x"1770665",
    x"17702A4",
    x"176FEE4",
    x"176FB25",
    x"176F766",
    x"176F3A9",
    x"176EFEC",
    x"176EC31",
    x"176E876",
    x"176E4BD",
    x"176E104",
    x"176DD4C",
    x"176D995",
    x"176D5DF",
    x"176D22A",
    x"176CE76",
    x"176CAC3",
    x"176C711",
    x"176C360",
    x"176BFAF",
    x"176BC00",
    x"176B851",
    x"176B4A4",
    x"176B0F7",
    x"176AD4B",
    x"176A9A0",
    x"176A5F6",
    x"176A24D",
    x"1769EA5",
    x"1769AFE",
    x"1769758",
    x"17693B2",
    x"176900E",
    x"1768C6A",
    x"17688C8",
    x"1768526",
    x"1768185",
    x"1767DE5",
    x"1767A46",
    x"17676A8",
    x"176730B",
    x"1766F6E",
    x"1766BD3",
    x"1766839",
    x"176649F",
    x"1766106",
    x"1765D6E",
    x"17659D8",
    x"1765642",
    x"17652AC",
    x"1764F18",
    x"1764B85",
    x"17647F2",
    x"1764461",
    x"17640D0",
    x"1763D40",
    x"17639B2",
    x"1763624",
    x"1763297",
    x"1762F0A",
    x"1762B7F",
    x"17627F5",
    x"176246B",
    x"17620E2",
    x"1761D5B",
    x"17619D4",
    x"176164E",
    x"17612C9",
    x"1760F44",
    x"1760BC1",
    x"176083E",
    x"17604BD",
    x"176013C",
    x"175FDBC",
    x"175FA3D",
    x"175F6BF",
    x"175F342",
    x"175EFC5",
    x"175EC4A",
    x"175E8CF",
    x"175E555",
    x"175E1DD",
    x"175DE65",
    x"175DAED",
    x"175D777",
    x"175D402",
    x"175D08D",
    x"175CD19",
    x"175C9A7",
    x"175C635",
    x"175C2C3",
    x"175BF53",
    x"175BBE4",
    x"175B875",
    x"175B508",
    x"175B19B",
    x"175AE2F",
    x"175AAC4",
    x"175A759",
    x"175A3F0",
    x"175A087",
    x"1759D20",
    x"17599B9",
    x"1759653",
    x"17592EE",
    x"1758F89",
    x"1758C26",
    x"17588C3",
    x"1758562",
    x"1758201",
    x"1757EA1",
    x"1757B41",
    x"17577E3",
    x"1757485",
    x"1757129",
    x"1756DCD",
    x"1756A72",
    x"1756718",
    x"17563BE",
    x"1756066",
    x"1755D0E",
    x"17559B7",
    x"1755661",
    x"175530C",
    x"1754FB8",
    x"1754C64",
    x"1754911",
    x"17545C0",
    x"175426F",
    x"1753F1E",
    x"1753BCF",
    x"1753880",
    x"1753533",
    x"17531E6",
    x"1752E9A",
    x"1752B4F",
    x"1752804",
    x"17524BB",
    x"1752172",
    x"1751E2A",
    x"1751AE3",
    x"175179C",
    x"1751457",
    x"1751112",
    x"1750DCE",
    x"1750A8B",
    x"1750749",
    x"1750408",
    x"17500C7",
    x"174FD87",
    x"174FA48",
    x"174F70A",
    x"174F3CD",
    x"174F090",
    x"174ED54",
    x"174EA1A",
    x"174E6DF",
    x"174E3A6",
    x"174E06E",
    x"174DD36",
    x"174D9FF",
    x"174D6C9",
    x"174D394",
    x"174D05F",
    x"174CD2B",
    x"174C9F8",
    x"174C6C6",
    x"174C395",
    x"174C065",
    x"174BD35",
    x"174BA06",
    x"174B6D8",
    x"174B3AB",
    x"174B07E",
    x"174AD52",
    x"174AA27",
    x"174A6FD",
    x"174A3D4",
    x"174A0AB",
    x"1749D84",
    x"1749A5D",
    x"1749736",
    x"1749411",
    x"17490EC",
    x"1748DC9",
    x"1748AA5",
    x"1748783",
    x"1748462",
    x"1748141",
    x"1747E21",
    x"1747B02",
    x"17477E4",
    x"17474C6",
    x"17471A9",
    x"1746E8D",
    x"1746B72",
    x"1746857",
    x"174653E",
    x"1746225",
    x"1745F0D",
    x"1745BF5",
    x"17458DF",
    x"17455C9",
    x"17452B4",
    x"1744F9F",
    x"1744C8C",
    x"1744979",
    x"1744667",
    x"1744356",
    x"1744046",
    x"1743D36",
    x"1743A27",
    x"1743719",
    x"174340B",
    x"17430FF",
    x"1742DF3",
    x"1742AE8",
    x"17427DD",
    x"17424D4",
    x"17421CB",
    x"1741EC3",
    x"1741BBC",
    x"17418B5",
    x"17415AF",
    x"17412AA",
    x"1740FA6",
    x"1740CA2",
    x"17409A0",
    x"174069E",
    x"174039C",
    x"174009C",
    x"173FD9C",
    x"173FA9D",
    x"173F79F",
    x"173F4A1",
    x"173F1A4",
    x"173EEA8",
    x"173EBAD",
    x"173E8B3",
    x"173E5B9",
    x"173E2C0",
    x"173DFC7",
    x"173DCD0",
    x"173D9D9",
    x"173D6E3",
    x"173D3EE",
    x"173D0F9",
    x"173CE05",
    x"173CB12",
    x"173C81F",
    x"173C52E",
    x"173C23D",
    x"173BF4D",
    x"173BC5D",
    x"173B96F",
    x"173B681",
    x"173B393",
    x"173B0A7",
    x"173ADBB",
    x"173AAD0",
    x"173A7E6",
    x"173A4FC",
    x"173A213",
    x"1739F2B",
    x"1739C43",
    x"173995D",
    x"1739677",
    x"1739392",
    x"17390AD",
    x"1738DC9",
    x"1738AE6",
    x"1738804",
    x"1738522",
    x"1738241",
    x"1737F61",
    x"1737C81",
    x"17379A3",
    x"17376C5",
    x"17373E7",
    x"173710B",
    x"1736E2F",
    x"1736B54",
    x"1736879",
    x"173659F",
    x"17362C6",
    x"1735FEE",
    x"1735D16",
    x"1735A3F",
    x"1735769",
    x"1735494",
    x"17351BF",
    x"1734EEB",
    x"1734C17",
    x"1734945",
    x"1734673",
    x"17343A2",
    x"17340D1",
    x"1733E01",
    x"1733B32",
    x"1733864",
    x"1733596",
    x"17332C9",
    x"1732FFC",
    x"1732D31",
    x"1732A66",
    x"173279C",
    x"17324D2",
    x"1732209",
    x"1731F41",
    x"1731C7A",
    x"17319B3",
    x"17316ED",
    x"1731427",
    x"1731163",
    x"1730E9F",
    x"1730BDB",
    x"1730919",
    x"1730657",
    x"1730396",
    x"17300D5",
    x"172FE15",
    x"172FB56",
    x"172F897",
    x"172F5DA",
    x"172F31D",
    x"172F060",
    x"172EDA4",
    x"172EAE9",
    x"172E82F",
    x"172E575",
    x"172E2BC",
    x"172E004",
    x"172DD4C",
    x"172DA95",
    x"172D7DF",
    x"172D529",
    x"172D274",
    x"172CFC0",
    x"172CD0C",
    x"172CA59",
    x"172C7A7",
    x"172C4F6",
    x"172C245",
    x"172BF94",
    x"172BCE5",
    x"172BA36",
    x"172B788",
    x"172B4DA",
    x"172B22D",
    x"172AF81",
    x"172ACD6",
    x"172AA2B",
    x"172A781",
    x"172A4D7",
    x"172A22E",
    x"1729F86",
    x"1729CDE",
    x"1729A37",
    x"1729791",
    x"17294EC",
    x"1729247",
    x"1728FA3",
    x"1728CFF",
    x"1728A5C",
    x"17287BA",
    x"1728518",
    x"1728277",
    x"1727FD7",
    x"1727D37",
    x"1727A98",
    x"17277FA",
    x"172755C",
    x"17272BF",
    x"1727023",
    x"1726D87",
    x"1726AEC",
    x"1726852",
    x"17265B8",
    x"172631F",
    x"1726086",
    x"1725DEF",
    x"1725B58",
    x"17258C1",
    x"172562B",
    x"1725396",
    x"1725101",
    x"1724E6D",
    x"1724BDA",
    x"1724947",
    x"17246B6",
    x"1724424",
    x"1724193",
    x"1723F03",
    x"1723C74",
    x"17239E5",
    x"1723757",
    x"17234C9",
    x"172323D",
    x"1722FB0",
    x"1722D25",
    x"1722A9A",
    x"172280F",
    x"1722586",
    x"17222FD",
    x"1722074",
    x"1721DEC",
    x"1721B65",
    x"17218DF",
    x"1721659",
    x"17213D4",
    x"172114F",
    x"1720ECB",
    x"1720C48",
    x"17209C5",
    x"1720743",
    x"17204C1",
    x"1720240",
    x"171FFC0",
    x"171FD40",
    x"171FAC1",
    x"171F843",
    x"171F5C5",
    x"171F348",
    x"171F0CC",
    x"171EE50",
    x"171EBD4",
    x"171E95A",
    x"171E6E0",
    x"171E466",
    x"171E1EE",
    x"171DF75",
    x"171DCFE",
    x"171DA87",
    x"171D811",
    x"171D59B",
    x"171D326",
    x"171D0B1",
    x"171CE3D",
    x"171CBCA",
    x"171C958",
    x"171C6E6",
    x"171C474",
    x"171C203",
    x"171BF93",
    x"171BD23",
    x"171BAB5",
    x"171B846",
    x"171B5D8",
    x"171B36B",
    x"171B0FF",
    x"171AE93",
    x"171AC27",
    x"171A9BD",
    x"171A753",
    x"171A4E9",
    x"171A280",
    x"171A018",
    x"1719DB0",
    x"1719B49",
    x"17198E2",
    x"171967C",
    x"1719417",
    x"17191B2",
    x"1718F4E",
    x"1718CEB",
    x"1718A88",
    x"1718825",
    x"17185C4",
    x"1718363",
    x"1718102",
    x"1717EA2",
    x"1717C43",
    x"17179E4",
    x"1717786",
    x"1717528",
    x"17172CB",
    x"171706F",
    x"1716E13",
    x"1716BB8",
    x"171695D",
    x"1716703",
    x"17164AA",
    x"1716251",
    x"1715FF8",
    x"1715DA1",
    x"1715B4A",
    x"17158F3",
    x"171569D",
    x"1715448",
    x"17151F3",
    x"1714F9F",
    x"1714D4B",
    x"1714AF8",
    x"17148A6",
    x"1714654",
    x"1714403",
    x"17141B2",
    x"1713F62",
    x"1713D12",
    x"1713AC3",
    x"1713875",
    x"1713627",
    x"17133DA",
    x"171318D",
    x"1712F41",
    x"1712CF5",
    x"1712AAA",
    x"1712860",
    x"1712616",
    x"17123CD",
    x"1712184",
    x"1711F3C",
    x"1711CF5",
    x"1711AAE",
    x"1711867",
    x"1711622",
    x"17113DC",
    x"1711198",
    x"1710F54",
    x"1710D10",
    x"1710ACD",
    x"171088B",
    x"1710649",
    x"1710407",
    x"17101C7",
    x"170FF87",
    x"170FD47",
    x"170FB08",
    x"170F8C9",
    x"170F68C",
    x"170F44E",
    x"170F211",
    x"170EFD5",
    x"170ED99",
    x"170EB5E",
    x"170E924",
    x"170E6EA",
    x"170E4B0",
    x"170E277",
    x"170E03F",
    x"170DE07",
    x"170DBD0",
    x"170D999",
    x"170D763",
    x"170D52E",
    x"170D2F9",
    x"170D0C4",
    x"170CE90",
    x"170CC5D",
    x"170CA2A",
    x"170C7F8",
    x"170C5C6",
    x"170C395",
    x"170C164",
    x"170BF34",
    x"170BD05",
    x"170BAD6",
    x"170B8A7",
    x"170B679",
    x"170B44C",
    x"170B21F",
    x"170AFF3",
    x"170ADC7",
    x"170AB9C",
    x"170A971",
    x"170A747",
    x"170A51E",
    x"170A2F5",
    x"170A0CC",
    x"1709EA4",
    x"1709C7D",
    x"1709A56",
    x"1709830",
    x"170960A",
    x"17093E5",
    x"17091C0",
    x"1708F9C",
    x"1708D78",
    x"1708B55",
    x"1708933",
    x"1708711",
    x"17084EF",
    x"17082CE",
    x"17080AE",
    x"1707E8E",
    x"1707C6E",
    x"1707A50",
    x"1707831",
    x"1707613",
    x"17073F6",
    x"17071DA",
    x"1706FBD",
    x"1706DA2",
    x"1706B86",
    x"170696C",
    x"1706752",
    x"1706538",
    x"170631F",
    x"1706107",
    x"1705EEF",
    x"1705CD7",
    x"1705AC0",
    x"17058AA",
    x"1705694",
    x"170547F",
    x"170526A",
    x"1705055",
    x"1704E41",
    x"1704C2E",
    x"1704A1B",
    x"1704809",
    x"17045F7",
    x"17043E6",
    x"17041D5",
    x"1703FC5",
    x"1703DB6",
    x"1703BA6",
    x"1703998",
    x"170378A",
    x"170357C",
    x"170336F",
    x"1703162",
    x"1702F56",
    x"1702D4B",
    x"1702B3F",
    x"1702935",
    x"170272B",
    x"1702521",
    x"1702318",
    x"1702110",
    x"1701F08",
    x"1701D00",
    x"1701AF9",
    x"17018F3",
    x"17016ED",
    x"17014E7",
    x"17012E2",
    x"17010DE",
    x"1700EDA",
    x"1700CD6",
    x"1700AD4",
    x"17008D1",
    x"17006CF",
    x"17004CE",
    x"17002CD",
    x"17000CC",
    x"16FFD99",
    x"16FF99A",
    x"16FF59C",
    x"16FF19F",
    x"16FEDA3",
    x"16FE9A9",
    x"16FE5AF",
    x"16FE1B6",
    x"16FDDBE",
    x"16FD9C7",
    x"16FD5D1",
    x"16FD1DC",
    x"16FCDE8",
    x"16FC9F5",
    x"16FC603",
    x"16FC212",
    x"16FBE22",
    x"16FBA33",
    x"16FB645",
    x"16FB258",
    x"16FAE6C",
    x"16FAA81",
    x"16FA696",
    x"16FA2AD",
    x"16F9EC5",
    x"16F9ADE",
    x"16F96F8",
    x"16F9312",
    x"16F8F2E",
    x"16F8B4B",
    x"16F8768",
    x"16F8387",
    x"16F7FA7",
    x"16F7BC7",
    x"16F77E9",
    x"16F740B",
    x"16F702F",
    x"16F6C53",
    x"16F6879",
    x"16F649F",
    x"16F60C6",
    x"16F5CEF",
    x"16F5918",
    x"16F5542",
    x"16F516D",
    x"16F4D99",
    x"16F49C6",
    x"16F45F4",
    x"16F4223",
    x"16F3E53",
    x"16F3A84",
    x"16F36B6",
    x"16F32E9",
    x"16F2F1D",
    x"16F2B51",
    x"16F2787",
    x"16F23BE",
    x"16F1FF5",
    x"16F1C2E",
    x"16F1867",
    x"16F14A1",
    x"16F10DD",
    x"16F0D19",
    x"16F0956",
    x"16F0594",
    x"16F01D3",
    x"16EFE13",
    x"16EFA54",
    x"16EF696",
    x"16EF2D9",
    x"16EEF1D",
    x"16EEB61",
    x"16EE7A7",
    x"16EE3EE",
    x"16EE035",
    x"16EDC7E",
    x"16ED8C7",
    x"16ED511",
    x"16ED15C",
    x"16ECDA8",
    x"16EC9F5",
    x"16EC643",
    x"16EC292",
    x"16EBEE2",
    x"16EBB33",
    x"16EB785",
    x"16EB3D7",
    x"16EB02B",
    x"16EAC7F",
    x"16EA8D4",
    x"16EA52B",
    x"16EA182",
    x"16E9DDA",
    x"16E9A33",
    x"16E968D",
    x"16E92E8",
    x"16E8F43",
    x"16E8BA0",
    x"16E87FE",
    x"16E845C",
    x"16E80BB",
    x"16E7D1C",
    x"16E797D",
    x"16E75DF",
    x"16E7242",
    x"16E6EA6",
    x"16E6B0B",
    x"16E6770",
    x"16E63D7",
    x"16E603E",
    x"16E5CA7",
    x"16E5910",
    x"16E557A",
    x"16E51E5",
    x"16E4E51",
    x"16E4ABE",
    x"16E472C",
    x"16E439A",
    x"16E400A",
    x"16E3C7A",
    x"16E38EC",
    x"16E355E",
    x"16E31D1",
    x"16E2E45",
    x"16E2ABA",
    x"16E2730",
    x"16E23A6",
    x"16E201E",
    x"16E1C96",
    x"16E1910",
    x"16E158A",
    x"16E1205",
    x"16E0E81",
    x"16E0AFE",
    x"16E077B",
    x"16E03FA",
    x"16E0079",
    x"16DFCFA",
    x"16DF97B",
    x"16DF5FD",
    x"16DF280",
    x"16DEF04",
    x"16DEB88",
    x"16DE80E",
    x"16DE494",
    x"16DE11C",
    x"16DDDA4",
    x"16DDA2D",
    x"16DD6B7",
    x"16DD341",
    x"16DCFCD",
    x"16DCC59",
    x"16DC8E7",
    x"16DC575",
    x"16DC204",
    x"16DBE94",
    x"16DBB25",
    x"16DB7B6",
    x"16DB449",
    x"16DB0DC",
    x"16DAD71",
    x"16DAA06",
    x"16DA69C",
    x"16DA332",
    x"16D9FCA",
    x"16D9C62",
    x"16D98FC",
    x"16D9596",
    x"16D9231",
    x"16D8ECD",
    x"16D8B6A",
    x"16D8807",
    x"16D84A6",
    x"16D8145",
    x"16D7DE5",
    x"16D7A86",
    x"16D7728",
    x"16D73CA",
    x"16D706E",
    x"16D6D12",
    x"16D69B7",
    x"16D665D",
    x"16D6304",
    x"16D5FAC",
    x"16D5C54",
    x"16D58FD",
    x"16D55A8",
    x"16D5253",
    x"16D4EFE",
    x"16D4BAB",
    x"16D4859",
    x"16D4507",
    x"16D41B6",
    x"16D3E66",
    x"16D3B17",
    x"16D37C9",
    x"16D347B",
    x"16D312E",
    x"16D2DE2",
    x"16D2A97",
    x"16D274D",
    x"16D2404",
    x"16D20BB",
    x"16D1D73",
    x"16D1A2C",
    x"16D16E6",
    x"16D13A1",
    x"16D105C",
    x"16D0D19",
    x"16D09D6",
    x"16D0694",
    x"16D0353",
    x"16D0012",
    x"16CFCD3",
    x"16CF994",
    x"16CF656",
    x"16CF319",
    x"16CEFDC",
    x"16CECA1",
    x"16CE966",
    x"16CE62C",
    x"16CE2F3",
    x"16CDFBB",
    x"16CDC83",
    x"16CD94C",
    x"16CD616",
    x"16CD2E1",
    x"16CCFAD",
    x"16CCC79",
    x"16CC947",
    x"16CC615",
    x"16CC2E4",
    x"16CBFB3",
    x"16CBC84",
    x"16CB955",
    x"16CB627",
    x"16CB2FA",
    x"16CAFCE",
    x"16CACA2",
    x"16CA977",
    x"16CA64D",
    x"16CA324",
    x"16C9FFC",
    x"16C9CD4",
    x"16C99AD",
    x"16C9687",
    x"16C9362",
    x"16C903E",
    x"16C8D1A",
    x"16C89F7",
    x"16C86D5",
    x"16C83B4",
    x"16C8093",
    x"16C7D73",
    x"16C7A54",
    x"16C7736",
    x"16C7419",
    x"16C70FC",
    x"16C6DE0",
    x"16C6AC5",
    x"16C67AB",
    x"16C6491",
    x"16C6179",
    x"16C5E61",
    x"16C5B49",
    x"16C5833",
    x"16C551D",
    x"16C5208",
    x"16C4EF4",
    x"16C4BE1",
    x"16C48CE",
    x"16C45BD",
    x"16C42AB",
    x"16C3F9B",
    x"16C3C8C",
    x"16C397D",
    x"16C366F",
    x"16C3362",
    x"16C3055",
    x"16C2D4A",
    x"16C2A3F",
    x"16C2734",
    x"16C242B",
    x"16C2122",
    x"16C1E1A",
    x"16C1B13",
    x"16C180D",
    x"16C1507",
    x"16C1202",
    x"16C0EFE",
    x"16C0BFB",
    x"16C08F8",
    x"16C05F6",
    x"16C02F5",
    x"16BFFF5",
    x"16BFCF5",
    x"16BF9F6",
    x"16BF6F8",
    x"16BF3FB",
    x"16BF0FE",
    x"16BEE02",
    x"16BEB07",
    x"16BE80D",
    x"16BE513",
    x"16BE21A",
    x"16BDF22",
    x"16BDC2B",
    x"16BD934",
    x"16BD63E",
    x"16BD349",
    x"16BD055",
    x"16BCD61",
    x"16BCA6E",
    x"16BC77C",
    x"16BC48A",
    x"16BC199",
    x"16BBEA9",
    x"16BBBBA",
    x"16BB8CB",
    x"16BB5DE",
    x"16BB2F1",
    x"16BB004",
    x"16BAD19",
    x"16BAA2E",
    x"16BA743",
    x"16BA45A",
    x"16BA171",
    x"16B9E89",
    x"16B9BA2",
    x"16B98BB",
    x"16B95D6",
    x"16B92F1",
    x"16B900C",
    x"16B8D29",
    x"16B8A46",
    x"16B8763",
    x"16B8482",
    x"16B81A1",
    x"16B7EC1",
    x"16B7BE2",
    x"16B7903",
    x"16B7625",
    x"16B7348",
    x"16B706C",
    x"16B6D90",
    x"16B6AB5",
    x"16B67DA",
    x"16B6501",
    x"16B6228",
    x"16B5F50",
    x"16B5C78",
    x"16B59A2",
    x"16B56CC",
    x"16B53F6",
    x"16B5122",
    x"16B4E4E",
    x"16B4B7A",
    x"16B48A8",
    x"16B45D6",
    x"16B4305",
    x"16B4035",
    x"16B3D65",
    x"16B3A96",
    x"16B37C8",
    x"16B34FA",
    x"16B322D",
    x"16B2F61",
    x"16B2C95",
    x"16B29CB",
    x"16B2700",
    x"16B2437",
    x"16B216E",
    x"16B1EA6",
    x"16B1BDF",
    x"16B1918",
    x"16B1652",
    x"16B138D",
    x"16B10C9",
    x"16B0E05",
    x"16B0B42",
    x"16B087F",
    x"16B05BD",
    x"16B02FC",
    x"16B003C",
    x"16AFD7C",
    x"16AFABD",
    x"16AF7FF",
    x"16AF541",
    x"16AF284",
    x"16AEFC8",
    x"16AED0C",
    x"16AEA51",
    x"16AE797",
    x"16AE4DE",
    x"16AE225",
    x"16ADF6D",
    x"16ADCB5",
    x"16AD9FE",
    x"16AD748",
    x"16AD493",
    x"16AD1DE",
    x"16ACF2A",
    x"16ACC76",
    x"16AC9C3",
    x"16AC711",
    x"16AC460",
    x"16AC1AF",
    x"16ABEFF",
    x"16ABC50",
    x"16AB9A1",
    x"16AB6F3",
    x"16AB445",
    x"16AB199",
    x"16AAEED",
    x"16AAC41",
    x"16AA996",
    x"16AA6EC",
    x"16AA443",
    x"16AA19A",
    x"16A9EF2",
    x"16A9C4B",
    x"16A99A4",
    x"16A96FE",
    x"16A9459",
    x"16A91B4",
    x"16A8F10",
    x"16A8C6C",
    x"16A89C9",
    x"16A8727",
    x"16A8486",
    x"16A81E5",
    x"16A7F45",
    x"16A7CA5",
    x"16A7A07",
    x"16A7768",
    x"16A74CB",
    x"16A722E",
    x"16A6F92",
    x"16A6CF6",
    x"16A6A5B",
    x"16A67C1",
    x"16A6527",
    x"16A628F",
    x"16A5FF6",
    x"16A5D5F",
    x"16A5AC8",
    x"16A5831",
    x"16A559B",
    x"16A5306",
    x"16A5072",
    x"16A4DDE",
    x"16A4B4B",
    x"16A48B8",
    x"16A4627",
    x"16A4395",
    x"16A4105",
    x"16A3E75",
    x"16A3BE6",
    x"16A3957",
    x"16A36C9",
    x"16A343C",
    x"16A31AF",
    x"16A2F23",
    x"16A2C97",
    x"16A2A0C",
    x"16A2782",
    x"16A24F9",
    x"16A2270",
    x"16A1FE7",
    x"16A1D60",
    x"16A1AD9",
    x"16A1852",
    x"16A15CD",
    x"16A1347",
    x"16A10C3",
    x"16A0E3F",
    x"16A0BBC",
    x"16A0939",
    x"16A06B7",
    x"16A0436",
    x"16A01B5",
    x"169FF35",
    x"169FCB5",
    x"169FA37",
    x"169F7B8",
    x"169F53B",
    x"169F2BE",
    x"169F041",
    x"169EDC6",
    x"169EB4B",
    x"169E8D0",
    x"169E656",
    x"169E3DD",
    x"169E164",
    x"169DEEC",
    x"169DC75",
    x"169D9FE",
    x"169D788",
    x"169D512",
    x"169D29D",
    x"169D029",
    x"169CDB5",
    x"169CB42",
    x"169C8CF",
    x"169C65E",
    x"169C3EC",
    x"169C17C",
    x"169BF0C",
    x"169BC9C",
    x"169BA2D",
    x"169B7BF",
    x"169B551",
    x"169B2E4",
    x"169B078",
    x"169AE0C",
    x"169ABA1",
    x"169A936",
    x"169A6CC",
    x"169A463",
    x"169A1FA",
    x"1699F92",
    x"1699D2A",
    x"1699AC3",
    x"169985D",
    x"16995F7",
    x"1699392",
    x"169912D",
    x"1698EC9",
    x"1698C66",
    x"1698A03",
    x"16987A1",
    x"169853F",
    x"16982DE",
    x"169807E",
    x"1697E1E",
    x"1697BBF",
    x"1697960",
    x"1697702",
    x"16974A5",
    x"1697248",
    x"1696FEC",
    x"1696D90",
    x"1696B35",
    x"16968DA",
    x"1696680",
    x"1696427",
    x"16961CE",
    x"1695F76",
    x"1695D1F",
    x"1695AC8",
    x"1695871",
    x"169561B",
    x"16953C6",
    x"1695171",
    x"1694F1D",
    x"1694CCA",
    x"1694A77",
    x"1694825",
    x"16945D3",
    x"1694382",
    x"1694131",
    x"1693EE1",
    x"1693C92",
    x"1693A43",
    x"16937F5",
    x"16935A7",
    x"169335A",
    x"169310D",
    x"1692EC1",
    x"1692C76",
    x"1692A2B",
    x"16927E1",
    x"1692597",
    x"169234E",
    x"1692105",
    x"1691EBD",
    x"1691C76",
    x"1691A2F",
    x"16917E9",
    x"16915A3",
    x"169135E",
    x"169111A",
    x"1690ED6",
    x"1690C92",
    x"1690A4F",
    x"169080D",
    x"16905CB",
    x"169038A",
    x"1690149",
    x"168FF09",
    x"168FCCA",
    x"168FA8B",
    x"168F84D",
    x"168F60F",
    x"168F3D2",
    x"168F195",
    x"168EF59",
    x"168ED1D",
    x"168EAE2",
    x"168E8A8",
    x"168E66E",
    x"168E435",
    x"168E1FC",
    x"168DFC4",
    x"168DD8C",
    x"168DB55",
    x"168D91E",
    x"168D6E8",
    x"168D4B3",
    x"168D27E",
    x"168D04A",
    x"168CE16",
    x"168CBE3",
    x"168C9B0",
    x"168C77E",
    x"168C54C",
    x"168C31B",
    x"168C0EB",
    x"168BEBB",
    x"168BC8B",
    x"168BA5C",
    x"168B82E",
    x"168B600",
    x"168B3D3",
    x"168B1A6",
    x"168AF7A",
    x"168AD4F",
    x"168AB24",
    x"168A8F9",
    x"168A6CF",
    x"168A4A6",
    x"168A27D",
    x"168A054",
    x"1689E2D",
    x"1689C05",
    x"16899DF",
    x"16897B8",
    x"1689593",
    x"168936E",
    x"1689149",
    x"1688F25",
    x"1688D01",
    x"1688ADE",
    x"16888BC",
    x"168869A",
    x"1688479",
    x"1688258",
    x"1688037",
    x"1687E18",
    x"1687BF8",
    x"16879DA",
    x"16877BC",
    x"168759E",
    x"1687381",
    x"1687164",
    x"1686F48",
    x"1686D2C",
    x"1686B11",
    x"16868F7",
    x"16866DD",
    x"16864C3",
    x"16862AB",
    x"1686092",
    x"1685E7A",
    x"1685C63",
    x"1685A4C",
    x"1685836",
    x"1685620",
    x"168540B",
    x"16851F6",
    x"1684FE2",
    x"1684DCE",
    x"1684BBB",
    x"16849A8",
    x"1684796",
    x"1684584",
    x"1684373",
    x"1684163",
    x"1683F53",
    x"1683D43",
    x"1683B34",
    x"1683925",
    x"1683717",
    x"168350A",
    x"16832FD",
    x"16830F0",
    x"1682EE4",
    x"1682CD9",
    x"1682ACE",
    x"16828C3",
    x"16826BA",
    x"16824B0",
    x"16822A7",
    x"168209F",
    x"1681E97",
    x"1681C8F",
    x"1681A89",
    x"1681882",
    x"168167C",
    x"1681477",
    x"1681272",
    x"168106E",
    x"1680E6A",
    x"1680C67",
    x"1680A64",
    x"1680861",
    x"168065F",
    x"168045E",
    x"168025D",
    x"168005D",
    x"167FCBB",
    x"167F8BC",
    x"167F4BE",
    x"167F0C2",
    x"167ECC6",
    x"167E8CB",
    x"167E4D2",
    x"167E0D9",
    x"167DCE1",
    x"167D8EA",
    x"167D4F5",
    x"167D100",
    x"167CD0C",
    x"167C919",
    x"167C528",
    x"167C137",
    x"167BD47",
    x"167B958",
    x"167B56A",
    x"167B17D",
    x"167AD92",
    x"167A9A7",
    x"167A5BD",
    x"167A1D4",
    x"1679DEC",
    x"1679A05",
    x"167961F",
    x"167923A",
    x"1678E56",
    x"1678A73",
    x"1678690",
    x"16782AF",
    x"1677ECF",
    x"1677AF0",
    x"1677712",
    x"1677334",
    x"1676F58",
    x"1676B7D",
    x"16767A2",
    x"16763C9",
    x"1675FF0",
    x"1675C19",
    x"1675842",
    x"167546D",
    x"1675098",
    x"1674CC5",
    x"16748F2",
    x"1674520",
    x"167414F",
    x"1673D7F",
    x"16739B0",
    x"16735E3",
    x"1673216",
    x"1672E49",
    x"1672A7E",
    x"16726B4",
    x"16722EB",
    x"1671F23",
    x"1671B5B",
    x"1671795",
    x"16713D0",
    x"167100B",
    x"1670C48",
    x"1670885",
    x"16704C3",
    x"1670103",
    x"166FD43",
    x"166F984",
    x"166F5C6",
    x"166F209",
    x"166EE4D",
    x"166EA92",
    x"166E6D8",
    x"166E31F",
    x"166DF66",
    x"166DBAF",
    x"166D7F8",
    x"166D443",
    x"166D08E",
    x"166CCDB",
    x"166C928",
    x"166C576",
    x"166C1C5",
    x"166BE15",
    x"166BA66",
    x"166B6B8",
    x"166B30B",
    x"166AF5E",
    x"166ABB3",
    x"166A809",
    x"166A45F",
    x"166A0B6",
    x"1669D0F",
    x"1669968",
    x"16695C2",
    x"166921D",
    x"1668E79",
    x"1668AD6",
    x"1668733",
    x"1668392",
    x"1667FF2",
    x"1667C52",
    x"16678B4",
    x"1667516",
    x"1667179",
    x"1666DDD",
    x"1666A42",
    x"16666A8",
    x"166630F",
    x"1665F76",
    x"1665BDF",
    x"1665848",
    x"16654B3",
    x"166511E",
    x"1664D8A",
    x"16649F7",
    x"1664665",
    x"16642D4",
    x"1663F44",
    x"1663BB5",
    x"1663826",
    x"1663498",
    x"166310C",
    x"1662D80",
    x"16629F5",
    x"166266B",
    x"16622E2",
    x"1661F5A",
    x"1661BD2",
    x"166184C",
    x"16614C6",
    x"1661141",
    x"1660DBD",
    x"1660A3A",
    x"16606B8",
    x"1660337",
    x"165FFB7",
    x"165FC37",
    x"165F8B8",
    x"165F53B",
    x"165F1BE",
    x"165EE42",
    x"165EAC7",
    x"165E74C",
    x"165E3D3",
    x"165E05B",
    x"165DCE3",
    x"165D96C",
    x"165D5F6",
    x"165D281",
    x"165CF0D",
    x"165CB9A",
    x"165C827",
    x"165C4B6",
    x"165C145",
    x"165BDD5",
    x"165BA66",
    x"165B6F8",
    x"165B38A",
    x"165B01E",
    x"165ACB2",
    x"165A948",
    x"165A5DE",
    x"165A275",
    x"1659F0C",
    x"1659BA5",
    x"165983F",
    x"16594D9",
    x"1659174",
    x"1658E10",
    x"1658AAD",
    x"165874B",
    x"16583EA",
    x"1658089",
    x"1657D29",
    x"16579CA",
    x"165766C",
    x"165730F",
    x"1656FB3",
    x"1656C57",
    x"16568FD",
    x"16565A3",
    x"165624A",
    x"1655EF2",
    x"1655B9A",
    x"1655844",
    x"16554EE",
    x"1655199",
    x"1654E45",
    x"1654AF2",
    x"16547A0",
    x"165444E",
    x"16540FE",
    x"1653DAE",
    x"1653A5F",
    x"1653711",
    x"16533C3",
    x"1653077",
    x"1652D2B",
    x"16529E0",
    x"1652696",
    x"165234D",
    x"1652005",
    x"1651CBD",
    x"1651976",
    x"1651630",
    x"16512EB",
    x"1650FA7",
    x"1650C63",
    x"1650921",
    x"16505DF",
    x"165029E",
    x"164FF5D",
    x"164FC1E",
    x"164F8DF",
    x"164F5A2",
    x"164F265",
    x"164EF28",
    x"164EBED",
    x"164E8B2",
    x"164E579",
    x"164E240",
    x"164DF08",
    x"164DBD0",
    x"164D89A",
    x"164D564",
    x"164D22F",
    x"164CEFB",
    x"164CBC7",
    x"164C895",
    x"164C563",
    x"164C232",
    x"164BF02",
    x"164BBD3",
    x"164B8A4",
    x"164B576",
    x"164B249",
    x"164AF1D",
    x"164ABF2",
    x"164A8C7",
    x"164A59D",
    x"164A274",
    x"1649F4C",
    x"1649C25",
    x"16498FE",
    x"16495D8",
    x"16492B3",
    x"1648F8F",
    x"1648C6B",
    x"1648949",
    x"1648627",
    x"1648306",
    x"1647FE5",
    x"1647CC6",
    x"16479A7",
    x"1647689",
    x"164736C",
    x"164704F",
    x"1646D33",
    x"1646A19",
    x"16466FE",
    x"16463E5",
    x"16460CC",
    x"1645DB5",
    x"1645A9E",
    x"1645787",
    x"1645472",
    x"164515D",
    x"1644E49",
    x"1644B36",
    x"1644824",
    x"1644512",
    x"1644201",
    x"1643EF1",
    x"1643BE2",
    x"16438D3",
    x"16435C5",
    x"16432B8",
    x"1642FAC",
    x"1642CA0",
    x"1642995",
    x"164268B",
    x"1642382",
    x"164207A",
    x"1641D72",
    x"1641A6B",
    x"1641765",
    x"164145F",
    x"164115B",
    x"1640E57",
    x"1640B53",
    x"1640851",
    x"164054F",
    x"164024E",
    x"163FF4E",
    x"163FC4F",
    x"163F950",
    x"163F652",
    x"163F355",
    x"163F058",
    x"163ED5D",
    x"163EA62",
    x"163E767",
    x"163E46E",
    x"163E175",
    x"163DE7D",
    x"163DB86",
    x"163D88F",
    x"163D59A",
    x"163D2A5",
    x"163CFB0",
    x"163CCBD",
    x"163C9CA",
    x"163C6D8",
    x"163C3E7",
    x"163C0F6",
    x"163BE06",
    x"163BB17",
    x"163B828",
    x"163B53B",
    x"163B24E",
    x"163AF62",
    x"163AC76",
    x"163A98B",
    x"163A6A1",
    x"163A3B8",
    x"163A0D0",
    x"1639DE8",
    x"1639B01",
    x"163981A",
    x"1639535",
    x"1639250",
    x"1638F6B",
    x"1638C88",
    x"16389A5",
    x"16386C3",
    x"16383E2",
    x"1638101",
    x"1637E21",
    x"1637B42",
    x"1637864",
    x"1637586",
    x"16372A9",
    x"1636FCD",
    x"1636CF1",
    x"1636A16",
    x"163673C",
    x"1636462",
    x"163618A",
    x"1635EB2",
    x"1635BDA",
    x"1635904",
    x"163562E",
    x"1635359",
    x"1635084",
    x"1634DB0",
    x"1634ADD",
    x"163480B",
    x"1634539",
    x"1634268",
    x"1633F98",
    x"1633CC9",
    x"16339FA",
    x"163372C",
    x"163345E",
    x"1633191",
    x"1632EC5",
    x"1632BFA",
    x"163292F",
    x"1632665",
    x"163239C",
    x"16320D4",
    x"1631E0C",
    x"1631B45",
    x"163187E",
    x"16315B8",
    x"16312F3",
    x"163102F",
    x"1630D6B",
    x"1630AA8",
    x"16307E6",
    x"1630524",
    x"1630263",
    x"162FFA3",
    x"162FCE3",
    x"162FA25",
    x"162F766",
    x"162F4A9",
    x"162F1EC",
    x"162EF30",
    x"162EC74",
    x"162E9BA",
    x"162E700",
    x"162E446",
    x"162E18D",
    x"162DED5",
    x"162DC1E",
    x"162D967",
    x"162D6B1",
    x"162D3FC",
    x"162D147",
    x"162CE93",
    x"162CBE0",
    x"162C92D",
    x"162C67B",
    x"162C3CA",
    x"162C11A",
    x"162BE6A",
    x"162BBBA",
    x"162B90C",
    x"162B65E",
    x"162B3B1",
    x"162B104",
    x"162AE58",
    x"162ABAD",
    x"162A902",
    x"162A658",
    x"162A3AF",
    x"162A106",
    x"1629E5F",
    x"1629BB7",
    x"1629911",
    x"162966B",
    x"16293C5",
    x"1629121",
    x"1628E7D",
    x"1628BDA",
    x"1628937",
    x"1628695",
    x"16283F4",
    x"1628153",
    x"1627EB3",
    x"1627C14",
    x"1627975",
    x"16276D7",
    x"162743A",
    x"162719D",
    x"1626F01",
    x"1626C65",
    x"16269CB",
    x"1626730",
    x"1626497",
    x"16261FE",
    x"1625F66",
    x"1625CCE",
    x"1625A38",
    x"16257A1",
    x"162550C",
    x"1625277",
    x"1624FE2",
    x"1624D4F",
    x"1624ABC",
    x"1624829",
    x"1624598",
    x"1624307",
    x"1624076",
    x"1623DE6",
    x"1623B57",
    x"16238C9",
    x"162363B",
    x"16233AE",
    x"1623121",
    x"1622E95",
    x"1622C0A",
    x"162297F",
    x"16226F5",
    x"162246C",
    x"16221E3",
    x"1621F5B",
    x"1621CD3",
    x"1621A4C",
    x"16217C6",
    x"1621540",
    x"16212BB",
    x"1621037",
    x"1620DB3",
    x"1620B30",
    x"16208AE",
    x"162062C",
    x"16203AB",
    x"162012A",
    x"161FEAA",
    x"161FC2B",
    x"161F9AC",
    x"161F72E",
    x"161F4B0",
    x"161F233",
    x"161EFB7",
    x"161ED3C",
    x"161EAC1",
    x"161E846",
    x"161E5CC",
    x"161E353",
    x"161E0DB",
    x"161DE63",
    x"161DBEC",
    x"161D975",
    x"161D6FF",
    x"161D489",
    x"161D215",
    x"161CFA0",
    x"161CD2D",
    x"161CABA",
    x"161C847",
    x"161C5D6",
    x"161C364",
    x"161C0F4",
    x"161BE84",
    x"161BC15",
    x"161B9A6",
    x"161B738",
    x"161B4CA",
    x"161B25D",
    x"161AFF1",
    x"161AD85",
    x"161AB1A",
    x"161A8B0",
    x"161A646",
    x"161A3DD",
    x"161A174",
    x"1619F0C",
    x"1619CA5",
    x"1619A3E",
    x"16197D7",
    x"1619572",
    x"161930D",
    x"16190A8",
    x"1618E44",
    x"1618BE1",
    x"161897E",
    x"161871C",
    x"16184BB",
    x"161825A",
    x"1617FFA",
    x"1617D9A",
    x"1617B3B",
    x"16178DC",
    x"161767F",
    x"1617421",
    x"16171C4",
    x"1616F68",
    x"1616D0D",
    x"1616AB2",
    x"1616857",
    x"16165FE",
    x"16163A4",
    x"161614C",
    x"1615EF4",
    x"1615C9C",
    x"1615A45",
    x"16157EF",
    x"1615599",
    x"1615344",
    x"16150F0",
    x"1614E9C",
    x"1614C49",
    x"16149F6",
    x"16147A4",
    x"1614552",
    x"1614301",
    x"16140B0",
    x"1613E61",
    x"1613C11",
    x"16139C3",
    x"1613774",
    x"1613527",
    x"16132DA",
    x"161308D",
    x"1612E42",
    x"1612BF6",
    x"16129AC",
    x"1612761",
    x"1612518",
    x"16122CF",
    x"1612086",
    x"1611E3F",
    x"1611BF7",
    x"16119B1",
    x"161176A",
    x"1611525",
    x"16112E0",
    x"161109B",
    x"1610E58",
    x"1610C14",
    x"16109D2",
    x"161078F",
    x"161054E",
    x"161030D",
    x"16100CC",
    x"160FE8C",
    x"160FC4D",
    x"160FA0E",
    x"160F7D0",
    x"160F592",
    x"160F355",
    x"160F119",
    x"160EEDD",
    x"160ECA1",
    x"160EA66",
    x"160E82C",
    x"160E5F2",
    x"160E3B9",
    x"160E180",
    x"160DF48",
    x"160DD11",
    x"160DADA",
    x"160D8A3",
    x"160D66D",
    x"160D438",
    x"160D203",
    x"160CFCF",
    x"160CD9B",
    x"160CB68",
    x"160C936",
    x"160C704",
    x"160C4D2",
    x"160C2A1",
    x"160C071",
    x"160BE41",
    x"160BC12",
    x"160B9E3",
    x"160B7B5",
    x"160B587",
    x"160B35A",
    x"160B12D",
    x"160AF01",
    x"160ACD6",
    x"160AAAB",
    x"160A881",
    x"160A657",
    x"160A42D",
    x"160A205",
    x"1609FDC",
    x"1609DB5",
    x"1609B8E",
    x"1609967",
    x"1609741",
    x"160951B",
    x"16092F6",
    x"16090D2",
    x"1608EAE",
    x"1608C8A",
    x"1608A68",
    x"1608845",
    x"1608623",
    x"1608402",
    x"16081E1",
    x"1607FC1",
    x"1607DA2",
    x"1607B82",
    x"1607964",
    x"1607746",
    x"1607528",
    x"160730B",
    x"16070EF",
    x"1606ED3",
    x"1606CB7",
    x"1606A9C",
    x"1606882",
    x"1606668",
    x"160644F",
    x"1606236",
    x"160601E",
    x"1605E06",
    x"1605BEF",
    x"16059D8",
    x"16057C2",
    x"16055AC",
    x"1605397",
    x"1605182",
    x"1604F6E",
    x"1604D5B",
    x"1604B47",
    x"1604935",
    x"1604723",
    x"1604511",
    x"1604300",
    x"16040F0",
    x"1603EE0",
    x"1603CD0",
    x"1603AC1",
    x"16038B3",
    x"16036A5",
    x"1603498",
    x"160328B",
    x"160307E",
    x"1602E73",
    x"1602C67",
    x"1602A5C",
    x"1602852",
    x"1602648",
    x"160243F",
    x"1602236",
    x"160202E",
    x"1601E26",
    x"1601C1F",
    x"1601A18",
    x"1601812",
    x"160160C",
    x"1601407",
    x"1601202",
    x"1600FFE",
    x"1600DFA",
    x"1600BF7",
    x"16009F4",
    x"16007F2",
    x"16005F0",
    x"16003EF",
    x"16001EE",
    x"15FFFDC",
    x"15FFBDC",
    x"15FF7DE",
    x"15FF3E0",
    x"15FEFE4",
    x"15FEBE9",
    x"15FE7EE",
    x"15FE3F5",
    x"15FDFFC",
    x"15FDC05",
    x"15FD80E",
    x"15FD419",
    x"15FD024",
    x"15FCC30",
    x"15FC83E",
    x"15FC44C",
    x"15FC05C",
    x"15FBC6C",
    x"15FB87E",
    x"15FB490",
    x"15FB0A3",
    x"15FACB8",
    x"15FA8CD",
    x"15FA4E3",
    x"15FA0FA",
    x"15F9D13",
    x"15F992C",
    x"15F9546",
    x"15F9161",
    x"15F8D7D",
    x"15F899B",
    x"15F85B9",
    x"15F81D8",
    x"15F7DF8",
    x"15F7A19",
    x"15F763B",
    x"15F725E",
    x"15F6E81",
    x"15F6AA6",
    x"15F66CC",
    x"15F62F3",
    x"15F5F1B",
    x"15F5B43",
    x"15F576D",
    x"15F5398",
    x"15F4FC3",
    x"15F4BF0",
    x"15F481D",
    x"15F444C",
    x"15F407B",
    x"15F3CAB",
    x"15F38DD",
    x"15F350F",
    x"15F3142",
    x"15F2D76",
    x"15F29AC",
    x"15F25E2",
    x"15F2219",
    x"15F1E51",
    x"15F1A89",
    x"15F16C3",
    x"15F12FE",
    x"15F0F3A",
    x"15F0B76",
    x"15F07B4",
    x"15F03F3",
    x"15F0032",
    x"15EFC72",
    x"15EF8B4",
    x"15EF4F6",
    x"15EF139",
    x"15EED7D",
    x"15EE9C3",
    x"15EE609",
    x"15EE250",
    x"15EDE97",
    x"15EDAE0",
    x"15ED72A",
    x"15ED375",
    x"15ECFC0",
    x"15ECC0D",
    x"15EC85A",
    x"15EC4A9",
    x"15EC0F8",
    x"15EBD48",
    x"15EB999",
    x"15EB5EB",
    x"15EB23E",
    x"15EAE92",
    x"15EAAE7",
    x"15EA73D",
    x"15EA393",
    x"15E9FEB",
    x"15E9C43",
    x"15E989D",
    x"15E94F7",
    x"15E9152",
    x"15E8DAE",
    x"15E8A0C",
    x"15E8669",
    x"15E82C8",
    x"15E7F28",
    x"15E7B89",
    x"15E77EA",
    x"15E744D",
    x"15E70B0",
    x"15E6D14",
    x"15E697A",
    x"15E65E0",
    x"15E6247",
    x"15E5EAF",
    x"15E5B17",
    x"15E5781",
    x"15E53EC",
    x"15E5057",
    x"15E4CC3",
    x"15E4931",
    x"15E459F",
    x"15E420E",
    x"15E3E7E",
    x"15E3AEF",
    x"15E3760",
    x"15E33D3",
    x"15E3046",
    x"15E2CBB",
    x"15E2930",
    x"15E25A6",
    x"15E221D",
    x"15E1E95",
    x"15E1B0E",
    x"15E1788",
    x"15E1402",
    x"15E107E",
    x"15E0CFA",
    x"15E0977",
    x"15E05F5",
    x"15E0274",
    x"15DFEF4",
    x"15DFB75",
    x"15DF7F6",
    x"15DF479",
    x"15DF0FC",
    x"15DED80",
    x"15DEA05",
    x"15DE68B",
    x"15DE312",
    x"15DDF9A",
    x"15DDC22",
    x"15DD8AC",
    x"15DD536",
    x"15DD1C1",
    x"15DCE4D",
    x"15DCADA",
    x"15DC768",
    x"15DC3F6",
    x"15DC086",
    x"15DBD16",
    x"15DB9A7",
    x"15DB639",
    x"15DB2CC",
    x"15DAF60",
    x"15DABF4",
    x"15DA88A",
    x"15DA520",
    x"15DA1B7",
    x"15D9E4F",
    x"15D9AE8",
    x"15D9782",
    x"15D941C",
    x"15D90B8",
    x"15D8D54",
    x"15D89F1",
    x"15D868F",
    x"15D832E",
    x"15D7FCD",
    x"15D7C6E",
    x"15D790F",
    x"15D75B1",
    x"15D7254",
    x"15D6EF8",
    x"15D6B9D",
    x"15D6842",
    x"15D64E9",
    x"15D6190",
    x"15D5E38",
    x"15D5AE1",
    x"15D578A",
    x"15D5435",
    x"15D50E0",
    x"15D4D8C",
    x"15D4A39",
    x"15D46E7",
    x"15D4396",
    x"15D4046",
    x"15D3CF6",
    x"15D39A7",
    x"15D3659",
    x"15D330C",
    x"15D2FC0",
    x"15D2C74",
    x"15D2929",
    x"15D25DF",
    x"15D2296",
    x"15D1F4E",
    x"15D1C07",
    x"15D18C0",
    x"15D157A",
    x"15D1235",
    x"15D0EF1",
    x"15D0BAE",
    x"15D086B",
    x"15D052A",
    x"15D01E9",
    x"15CFEA9",
    x"15CFB69",
    x"15CF82B",
    x"15CF4ED",
    x"15CF1B1",
    x"15CEE75",
    x"15CEB39",
    x"15CE7FF",
    x"15CE4C5",
    x"15CE18D",
    x"15CDE55",
    x"15CDB1D",
    x"15CD7E7",
    x"15CD4B1",
    x"15CD17D",
    x"15CCE49",
    x"15CCB15",
    x"15CC7E3",
    x"15CC4B2",
    x"15CC181",
    x"15CBE51",
    x"15CBB22",
    x"15CB7F3",
    x"15CB4C6",
    x"15CB199",
    x"15CAE6D",
    x"15CAB42",
    x"15CA817",
    x"15CA4EE",
    x"15CA1C5",
    x"15C9E9D",
    x"15C9B75",
    x"15C984F",
    x"15C9529",
    x"15C9204",
    x"15C8EE0",
    x"15C8BBD",
    x"15C889A",
    x"15C8579",
    x"15C8258",
    x"15C7F37",
    x"15C7C18",
    x"15C78F9",
    x"15C75DC",
    x"15C72BE",
    x"15C6FA2",
    x"15C6C87",
    x"15C696C",
    x"15C6652",
    x"15C6339",
    x"15C6020",
    x"15C5D09",
    x"15C59F2",
    x"15C56DC",
    x"15C53C6",
    x"15C50B2",
    x"15C4D9E",
    x"15C4A8B",
    x"15C4779",
    x"15C4467",
    x"15C4157",
    x"15C3E47",
    x"15C3B37",
    x"15C3829",
    x"15C351B",
    x"15C320E",
    x"15C2F02",
    x"15C2BF7",
    x"15C28EC",
    x"15C25E2",
    x"15C22D9",
    x"15C1FD1",
    x"15C1CC9",
    x"15C19C3",
    x"15C16BD",
    x"15C13B7",
    x"15C10B3",
    x"15C0DAF",
    x"15C0AAC",
    x"15C07AA",
    x"15C04A8",
    x"15C01A7",
    x"15BFEA7",
    x"15BFBA8",
    x"15BF8A9",
    x"15BF5AC",
    x"15BF2AF",
    x"15BEFB2",
    x"15BECB7",
    x"15BE9BC",
    x"15BE6C2",
    x"15BE3C9",
    x"15BE0D0",
    x"15BDDD8",
    x"15BDAE1",
    x"15BD7EB",
    x"15BD4F5",
    x"15BD200",
    x"15BCF0C",
    x"15BCC19",
    x"15BC926",
    x"15BC634",
    x"15BC343",
    x"15BC052",
    x"15BBD63",
    x"15BBA74",
    x"15BB786",
    x"15BB498",
    x"15BB1AB",
    x"15BAEBF",
    x"15BABD4",
    x"15BA8E9",
    x"15BA5FF",
    x"15BA316",
    x"15BA02E",
    x"15B9D46",
    x"15B9A5F",
    x"15B9779",
    x"15B9493",
    x"15B91AF",
    x"15B8ECB",
    x"15B8BE7",
    x"15B8905",
    x"15B8623",
    x"15B8342",
    x"15B8061",
    x"15B7D81",
    x"15B7AA2",
    x"15B77C4",
    x"15B74E7",
    x"15B720A",
    x"15B6F2E",
    x"15B6C52",
    x"15B6977",
    x"15B669D",
    x"15B63C4",
    x"15B60EB",
    x"15B5E14",
    x"15B5B3C",
    x"15B5866",
    x"15B5590",
    x"15B52BB",
    x"15B4FE7",
    x"15B4D13",
    x"15B4A40",
    x"15B476E",
    x"15B449D",
    x"15B41CC",
    x"15B3EFC",
    x"15B3C2C",
    x"15B395E",
    x"15B3690",
    x"15B33C2",
    x"15B30F6",
    x"15B2E2A",
    x"15B2B5F",
    x"15B2894",
    x"15B25CA",
    x"15B2301",
    x"15B2039",
    x"15B1D71",
    x"15B1AAA",
    x"15B17E4",
    x"15B151E",
    x"15B1259",
    x"15B0F95",
    x"15B0CD1",
    x"15B0A0F",
    x"15B074C",
    x"15B048B",
    x"15B01CA",
    x"15AFF0A",
    x"15AFC4B",
    x"15AF98C",
    x"15AF6CE",
    x"15AF411",
    x"15AF154",
    x"15AEE98",
    x"15AEBDD",
    x"15AE922",
    x"15AE668",
    x"15AE3AF",
    x"15AE0F6",
    x"15ADE3E",
    x"15ADB87",
    x"15AD8D0",
    x"15AD61B",
    x"15AD365",
    x"15AD0B1",
    x"15ACDFD",
    x"15ACB4A",
    x"15AC897",
    x"15AC5E6",
    x"15AC334",
    x"15AC084",
    x"15ABDD4",
    x"15ABB25",
    x"15AB877",
    x"15AB5C9",
    x"15AB31C",
    x"15AB06F",
    x"15AADC4",
    x"15AAB18",
    x"15AA86E",
    x"15AA5C4",
    x"15AA31B",
    x"15AA073",
    x"15A9DCB",
    x"15A9B24",
    x"15A987D",
    x"15A95D8",
    x"15A9332",
    x"15A908E",
    x"15A8DEA",
    x"15A8B47",
    x"15A88A4",
    x"15A8603",
    x"15A8361",
    x"15A80C1",
    x"15A7E21",
    x"15A7B82",
    x"15A78E3",
    x"15A7645",
    x"15A73A8",
    x"15A710C",
    x"15A6E70",
    x"15A6BD4",
    x"15A693A",
    x"15A66A0",
    x"15A6406",
    x"15A616E",
    x"15A5ED6",
    x"15A5C3E",
    x"15A59A8",
    x"15A5711",
    x"15A547C",
    x"15A51E7",
    x"15A4F53",
    x"15A4CC0",
    x"15A4A2D",
    x"15A479B",
    x"15A4509",
    x"15A4278",
    x"15A3FE8",
    x"15A3D58",
    x"15A3AC9",
    x"15A383B",
    x"15A35AD",
    x"15A3320",
    x"15A3093",
    x"15A2E08",
    x"15A2B7C",
    x"15A28F2",
    x"15A2668",
    x"15A23DF",
    x"15A2156",
    x"15A1ECE",
    x"15A1C47",
    x"15A19C0",
    x"15A173A",
    x"15A14B4",
    x"15A122F",
    x"15A0FAB",
    x"15A0D27",
    x"15A0AA4",
    x"15A0822",
    x"15A05A0",
    x"15A031F",
    x"15A009F",
    x"159FE1F",
    x"159FBA0",
    x"159F921",
    x"159F6A3",
    x"159F426",
    x"159F1A9",
    x"159EF2D",
    x"159ECB2",
    x"159EA37",
    x"159E7BC",
    x"159E543",
    x"159E2CA",
    x"159E051",
    x"159DDDA",
    x"159DB62",
    x"159D8EC",
    x"159D676",
    x"159D401",
    x"159D18C",
    x"159CF18",
    x"159CCA4",
    x"159CA32",
    x"159C7BF",
    x"159C54E",
    x"159C2DD",
    x"159C06C",
    x"159BDFD",
    x"159BB8D",
    x"159B91F",
    x"159B6B1",
    x"159B443",
    x"159B1D7",
    x"159AF6A",
    x"159ACFF",
    x"159AA94",
    x"159A82A",
    x"159A5C0",
    x"159A357",
    x"159A0EE",
    x"1599E86",
    x"1599C1F",
    x"15999B8",
    x"1599752",
    x"15994ED",
    x"1599288",
    x"1599023",
    x"1598DC0",
    x"1598B5C",
    x"15988FA",
    x"1598698",
    x"1598437",
    x"15981D6",
    x"1597F76",
    x"1597D16",
    x"1597AB7",
    x"1597859",
    x"15975FB",
    x"159739E",
    x"1597141",
    x"1596EE5",
    x"1596C8A",
    x"1596A2F",
    x"15967D5",
    x"159657B",
    x"1596322",
    x"15960C9",
    x"1595E71",
    x"1595C1A",
    x"15959C3",
    x"159576D",
    x"1595518",
    x"15952C3",
    x"159506E",
    x"1594E1A",
    x"1594BC7",
    x"1594975",
    x"1594723",
    x"15944D1",
    x"1594280",
    x"1594030",
    x"1593DE0",
    x"1593B91",
    x"1593942",
    x"15936F4",
    x"15934A7",
    x"159325A",
    x"159300E",
    x"1592DC2",
    x"1592B77",
    x"159292C",
    x"15926E2",
    x"1592499",
    x"1592250",
    x"1592008",
    x"1591DC0",
    x"1591B79",
    x"1591932",
    x"15916EC",
    x"15914A7",
    x"1591262",
    x"159101D",
    x"1590DDA",
    x"1590B96",
    x"1590954",
    x"1590712",
    x"15904D0",
    x"159028F",
    x"159004F",
    x"158FE0F",
    x"158FBD0",
    x"158F991",
    x"158F753",
    x"158F516",
    x"158F2D9",
    x"158F09C",
    x"158EE60",
    x"158EC25",
    x"158E9EA",
    x"158E7B0",
    x"158E576",
    x"158E33D",
    x"158E105",
    x"158DECD",
    x"158DC95",
    x"158DA5F",
    x"158D828",
    x"158D5F3",
    x"158D3BD",
    x"158D189",
    x"158CF55",
    x"158CD21",
    x"158CAEE",
    x"158C8BB",
    x"158C68A",
    x"158C458",
    x"158C227",
    x"158BFF7",
    x"158BDC7",
    x"158BB98",
    x"158B96A",
    x"158B73C",
    x"158B50E",
    x"158B2E1",
    x"158B0B5",
    x"158AE89",
    x"158AC5D",
    x"158AA32",
    x"158A808",
    x"158A5DE",
    x"158A3B5",
    x"158A18D",
    x"1589F64",
    x"1589D3D",
    x"1589B16",
    x"15898EF",
    x"15896C9",
    x"15894A4",
    x"158927F",
    x"158905B",
    x"1588E37",
    x"1588C14",
    x"15889F1",
    x"15887CF",
    x"15885AD",
    x"158838C",
    x"158816B",
    x"1587F4B",
    x"1587D2C",
    x"1587B0D",
    x"15878EE",
    x"15876D0",
    x"15874B3",
    x"1587296",
    x"1587079",
    x"1586E5D",
    x"1586C42",
    x"1586A27",
    x"158680D",
    x"15865F3",
    x"15863DA",
    x"15861C1",
    x"1585FA9",
    x"1585D92",
    x"1585B7A",
    x"1585964",
    x"158574E",
    x"1585538",
    x"1585323",
    x"158510F",
    x"1584EFB",
    x"1584CE7",
    x"1584AD4",
    x"15848C2",
    x"15846B0",
    x"158449E",
    x"158428D",
    x"158407D",
    x"1583E6D",
    x"1583C5E",
    x"1583A4F",
    x"1583841",
    x"1583633",
    x"1583426",
    x"1583219",
    x"158300D",
    x"1582E01",
    x"1582BF6",
    x"15829EB",
    x"15827E1",
    x"15825D7",
    x"15823CE",
    x"15821C5",
    x"1581FBD",
    x"1581DB5",
    x"1581BAE",
    x"15819A7",
    x"15817A1",
    x"158159B",
    x"1581396",
    x"1581192",
    x"1580F8D",
    x"1580D8A",
    x"1580B87",
    x"1580984",
    x"1580782",
    x"1580580",
    x"158037F",
    x"158017F",
    x"157FEFD",
    x"157FAFE",
    x"157F700",
    x"157F303",
    x"157EF06",
    x"157EB0B",
    x"157E711",
    x"157E318",
    x"157DF1F",
    x"157DB28",
    x"157D732",
    x"157D33C",
    x"157CF48",
    x"157CB55",
    x"157C762",
    x"157C371",
    x"157BF81",
    x"157BB91",
    x"157B7A3",
    x"157B3B6",
    x"157AFC9",
    x"157ABDE",
    x"157A7F3",
    x"157A40A",
    x"157A021",
    x"1579C3A",
    x"1579853",
    x"157946D",
    x"1579089",
    x"1578CA5",
    x"15788C2",
    x"15784E1",
    x"1578100",
    x"1577D20",
    x"1577941",
    x"1577564",
    x"1577187",
    x"1576DAB",
    x"15769D0",
    x"15765F6",
    x"157621D",
    x"1575E45",
    x"1575A6E",
    x"1575698",
    x"15752C3",
    x"1574EEE",
    x"1574B1B",
    x"1574749",
    x"1574377",
    x"1573FA7",
    x"1573BD8",
    x"1573809",
    x"157343C",
    x"157306F",
    x"1572CA3",
    x"15728D9",
    x"157250F",
    x"1572146",
    x"1571D7E",
    x"15719B7",
    x"15715F1",
    x"157122C",
    x"1570E68",
    x"1570AA5",
    x"15706E3",
    x"1570322",
    x"156FF61",
    x"156FBA2",
    x"156F7E4",
    x"156F426",
    x"156F06A",
    x"156ECAE",
    x"156E8F3",
    x"156E539",
    x"156E181",
    x"156DDC9",
    x"156DA12",
    x"156D65C",
    x"156D2A7",
    x"156CEF2",
    x"156CB3F",
    x"156C78D",
    x"156C3DB",
    x"156C02B",
    x"156BC7B",
    x"156B8CD",
    x"156B51F",
    x"156B172",
    x"156ADC6",
    x"156AA1B",
    x"156A671",
    x"156A2C8",
    x"1569F20",
    x"1569B78",
    x"15697D2",
    x"156942C",
    x"1569088",
    x"1568CE4",
    x"1568941",
    x"15685A0",
    x"15681FF",
    x"1567E5F",
    x"1567ABF",
    x"1567721",
    x"1567384",
    x"1566FE7",
    x"1566C4C",
    x"15668B1",
    x"1566517",
    x"156617F",
    x"1565DE7",
    x"1565A50",
    x"15656BA",
    x"1565324",
    x"1564F90",
    x"1564BFD",
    x"156486A",
    x"15644D8",
    x"1564148",
    x"1563DB8",
    x"1563A29",
    x"156369B",
    x"156330D",
    x"1562F81",
    x"1562BF6",
    x"156286B",
    x"15624E1",
    x"1562159",
    x"1561DD1",
    x"1561A4A",
    x"15616C4",
    x"156133E",
    x"1560FBA",
    x"1560C37",
    x"15608B4",
    x"1560532",
    x"15601B1",
    x"155FE31",
    x"155FAB2",
    x"155F734",
    x"155F3B7",
    x"155F03A",
    x"155ECBF",
    x"155E944",
    x"155E5CA",
    x"155E251",
    x"155DED9",
    x"155DB61",
    x"155D7EB",
    x"155D475",
    x"155D101",
    x"155CD8D",
    x"155CA1A",
    x"155C6A8",
    x"155C337",
    x"155BFC6",
    x"155BC57",
    x"155B8E8",
    x"155B57A",
    x"155B20D",
    x"155AEA1",
    x"155AB36",
    x"155A7CC",
    x"155A462",
    x"155A0FA",
    x"1559D92",
    x"1559A2B",
    x"15596C5",
    x"155935F",
    x"1558FFB",
    x"1558C97",
    x"1558935",
    x"15585D3",
    x"1558272",
    x"1557F12",
    x"1557BB2",
    x"1557854",
    x"15574F6",
    x"1557199",
    x"1556E3D",
    x"1556AE2",
    x"1556788",
    x"155642E",
    x"15560D6",
    x"1555D7E",
    x"1555A27",
    x"15556D1",
    x"155537C",
    x"1555027",
    x"1554CD3",
    x"1554981",
    x"155462F",
    x"15542DE",
    x"1553F8D",
    x"1553C3E",
    x"15538EF",
    x"15535A1",
    x"1553254",
    x"1552F08",
    x"1552BBD",
    x"1552872",
    x"1552529",
    x"15521E0",
    x"1551E98",
    x"1551B50",
    x"155180A",
    x"15514C4",
    x"1551180",
    x"1550E3C",
    x"1550AF8",
    x"15507B6",
    x"1550475",
    x"1550134",
    x"154FDF4",
    x"154FAB5",
    x"154F777",
    x"154F439",
    x"154F0FD",
    x"154EDC1",
    x"154EA86",
    x"154E74B",
    x"154E412",
    x"154E0D9",
    x"154DDA2",
    x"154DA6B",
    x"154D734",
    x"154D3FF",
    x"154D0CA",
    x"154CD97",
    x"154CA64",
    x"154C731",
    x"154C400",
    x"154C0CF",
    x"154BDA0",
    x"154BA71",
    x"154B742",
    x"154B415",
    x"154B0E8",
    x"154ADBD",
    x"154AA91",
    x"154A767",
    x"154A43E",
    x"154A115",
    x"1549DED",
    x"1549AC6",
    x"15497A0",
    x"154947A",
    x"1549156",
    x"1548E32",
    x"1548B0E",
    x"15487EC",
    x"15484CB",
    x"15481AA",
    x"1547E8A",
    x"1547B6A",
    x"154784C",
    x"154752E",
    x"1547211",
    x"1546EF5",
    x"1546BDA",
    x"15468BF",
    x"15465A6",
    x"154628D",
    x"1545F74",
    x"1545C5D",
    x"1545946",
    x"1545630",
    x"154531B",
    x"1545007",
    x"1544CF3",
    x"15449E0",
    x"15446CE",
    x"15443BD",
    x"15440AC",
    x"1543D9C",
    x"1543A8D",
    x"154377F",
    x"1543472",
    x"1543165",
    x"1542E59",
    x"1542B4E",
    x"1542843",
    x"154253A",
    x"1542231",
    x"1541F28",
    x"1541C21",
    x"154191A",
    x"1541615",
    x"154130F",
    x"154100B",
    x"1540D07",
    x"1540A04",
    x"1540702",
    x"1540401",
    x"1540100",
    x"153FE00",
    x"153FB01",
    x"153F803",
    x"153F505",
    x"153F208",
    x"153EF0C",
    x"153EC11",
    x"153E916",
    x"153E61C",
    x"153E323",
    x"153E02B",
    x"153DD33",
    x"153DA3C",
    x"153D746",
    x"153D451",
    x"153D15C",
    x"153CE68",
    x"153CB75",
    x"153C882",
    x"153C590",
    x"153C29F",
    x"153BFAF",
    x"153BCC0",
    x"153B9D1",
    x"153B6E3",
    x"153B3F5",
    x"153B109",
    x"153AE1D",
    x"153AB32",
    x"153A847",
    x"153A55D",
    x"153A274",
    x"1539F8C",
    x"1539CA5",
    x"15399BE",
    x"15396D8",
    x"15393F2",
    x"153910E",
    x"1538E2A",
    x"1538B47",
    x"1538864",
    x"1538583",
    x"15382A2",
    x"1537FC1",
    x"1537CE2",
    x"1537A03",
    x"1537725",
    x"1537447",
    x"153716B",
    x"1536E8F",
    x"1536BB3",
    x"15368D9",
    x"15365FF",
    x"1536326",
    x"153604D",
    x"1535D76",
    x"1535A9F",
    x"15357C8",
    x"15354F3",
    x"153521E",
    x"1534F4A",
    x"1534C76",
    x"15349A3",
    x"15346D1",
    x"1534400",
    x"153412F",
    x"1533E5F",
    x"1533B90",
    x"15338C2",
    x"15335F4",
    x"1533327",
    x"153305A",
    x"1532D8E",
    x"1532AC3",
    x"15327F9",
    x"153252F",
    x"1532266",
    x"1531F9E",
    x"1531CD7",
    x"1531A10",
    x"153174A",
    x"1531484",
    x"15311BF",
    x"1530EFB",
    x"1530C38",
    x"1530975",
    x"15306B3",
    x"15303F2",
    x"1530131",
    x"152FE71",
    x"152FBB2",
    x"152F8F3",
    x"152F635",
    x"152F378",
    x"152F0BC",
    x"152EE00",
    x"152EB45",
    x"152E88A",
    x"152E5D0",
    x"152E317",
    x"152E05F",
    x"152DDA7",
    x"152DAF0",
    x"152D83A",
    x"152D584",
    x"152D2CF",
    x"152D01B",
    x"152CD67",
    x"152CAB4",
    x"152C801",
    x"152C550",
    x"152C29F",
    x"152BFEE",
    x"152BD3F",
    x"152BA90",
    x"152B7E2",
    x"152B534",
    x"152B287",
    x"152AFDB",
    x"152AD2F",
    x"152AA84",
    x"152A7DA",
    x"152A530",
    x"152A287",
    x"1529FDF",
    x"1529D37",
    x"1529A90",
    x"15297EA",
    x"1529544",
    x"152929F",
    x"1528FFB",
    x"1528D57",
    x"1528AB4",
    x"1528812",
    x"1528570",
    x"15282CF",
    x"152802F",
    x"1527D8F",
    x"1527AF0",
    x"1527852",
    x"15275B4",
    x"1527317",
    x"152707A",
    x"1526DDF",
    x"1526B43",
    x"15268A9",
    x"152660F",
    x"1526376",
    x"15260DD",
    x"1525E46",
    x"1525BAE",
    x"1525918",
    x"1525682",
    x"15253EC",
    x"1525158",
    x"1524EC4",
    x"1524C30",
    x"152499E",
    x"152470C",
    x"152447A",
    x"15241E9",
    x"1523F59",
    x"1523CCA",
    x"1523A3B",
    x"15237AD",
    x"152351F",
    x"1523292",
    x"1523006",
    x"1522D7A",
    x"1522AEF",
    x"1522864",
    x"15225DB",
    x"1522352",
    x"15220C9",
    x"1521E41",
    x"1521BBA",
    x"1521933",
    x"15216AD",
    x"1521428",
    x"15211A3",
    x"1520F1F",
    x"1520C9C",
    x"1520A19",
    x"1520797",
    x"1520515",
    x"1520294",
    x"1520014",
    x"151FD94",
    x"151FB15",
    x"151F897",
    x"151F619",
    x"151F39B",
    x"151F11F",
    x"151EEA3",
    x"151EC28",
    x"151E9AD",
    x"151E733",
    x"151E4B9",
    x"151E240",
    x"151DFC8",
    x"151DD50",
    x"151DAD9",
    x"151D863",
    x"151D5ED",
    x"151D378",
    x"151D104",
    x"151CE90",
    x"151CC1C",
    x"151C9A9",
    x"151C737",
    x"151C4C6",
    x"151C255",
    x"151BFE5",
    x"151BD75",
    x"151BB06",
    x"151B898",
    x"151B62A",
    x"151B3BC",
    x"151B150",
    x"151AEE4",
    x"151AC78",
    x"151AA0E",
    x"151A7A3",
    x"151A53A",
    x"151A2D1",
    x"151A068",
    x"1519E01",
    x"1519B99",
    x"1519933",
    x"15196CD",
    x"1519467",
    x"1519203",
    x"1518F9E",
    x"1518D3B",
    x"1518AD8",
    x"1518875",
    x"1518613",
    x"15183B2",
    x"1518152",
    x"1517EF2",
    x"1517C92",
    x"1517A33",
    x"15177D5",
    x"1517577",
    x"151731A",
    x"15170BE",
    x"1516E62",
    x"1516C07",
    x"15169AC",
    x"1516752",
    x"15164F8",
    x"151629F",
    x"1516047",
    x"1515DEF",
    x"1515B98",
    x"1515941",
    x"15156EB",
    x"1515496",
    x"1515241",
    x"1514FED",
    x"1514D99",
    x"1514B46",
    x"15148F3",
    x"15146A2",
    x"1514450",
    x"15141FF",
    x"1513FAF",
    x"1513D60",
    x"1513B10",
    x"15138C2",
    x"1513674",
    x"1513427",
    x"15131DA",
    x"1512F8E",
    x"1512D42",
    x"1512AF7",
    x"15128AD",
    x"1512663",
    x"151241A",
    x"15121D1",
    x"1511F89",
    x"1511D41",
    x"1511AFA",
    x"15118B4",
    x"151166E",
    x"1511428",
    x"15111E4",
    x"1510F9F",
    x"1510D5C",
    x"1510B19",
    x"15108D6",
    x"1510694",
    x"1510453",
    x"1510212",
    x"150FFD2",
    x"150FD92",
    x"150FB53",
    x"150F915",
    x"150F6D7",
    x"150F499",
    x"150F25C",
    x"150F020",
    x"150EDE4",
    x"150EBA9",
    x"150E96E",
    x"150E734",
    x"150E4FB",
    x"150E2C2",
    x"150E089",
    x"150DE52",
    x"150DC1A",
    x"150D9E3",
    x"150D7AD",
    x"150D578",
    x"150D343",
    x"150D10E",
    x"150CEDA",
    x"150CCA7",
    x"150CA74",
    x"150C841",
    x"150C610",
    x"150C3DE",
    x"150C1AE",
    x"150BF7D",
    x"150BD4E",
    x"150BB1F",
    x"150B8F0",
    x"150B6C2",
    x"150B495",
    x"150B268",
    x"150B03C",
    x"150AE10",
    x"150ABE5",
    x"150A9BA",
    x"150A790",
    x"150A566",
    x"150A33D",
    x"150A115",
    x"1509EED",
    x"1509CC5",
    x"1509A9E",
    x"1509878",
    x"1509652",
    x"150942D",
    x"1509208",
    x"1508FE4",
    x"1508DC0",
    x"1508B9D",
    x"150897A",
    x"1508758",
    x"1508536",
    x"1508315",
    x"15080F5",
    x"1507ED5",
    x"1507CB6",
    x"1507A97",
    x"1507878",
    x"150765A",
    x"150743D",
    x"1507220",
    x"1507004",
    x"1506DE8",
    x"1506BCD",
    x"15069B2",
    x"1506798",
    x"150657F",
    x"1506365",
    x"150614D",
    x"1505F35",
    x"1505D1D",
    x"1505B06",
    x"15058F0",
    x"15056DA",
    x"15054C4",
    x"15052AF",
    x"150509B",
    x"1504E87",
    x"1504C74",
    x"1504A61",
    x"150484E",
    x"150463D",
    x"150442B",
    x"150421B",
    x"150400A",
    x"1503DFB",
    x"1503BEB",
    x"15039DD",
    x"15037CE",
    x"15035C1",
    x"15033B4",
    x"15031A7",
    x"1502F9B",
    x"1502D8F",
    x"1502B84",
    x"1502979",
    x"150276F",
    x"1502566",
    x"150235C",
    x"1502154",
    x"1501F4C",
    x"1501D44",
    x"1501B3D",
    x"1501937",
    x"1501731",
    x"150152B",
    x"1501326",
    x"1501121",
    x"1500F1D",
    x"1500D1A",
    x"1500B17",
    x"1500914",
    x"1500712",
    x"1500511",
    x"1500310",
    x"150010F",
    x"14FFE1F",
    x"14FFA20",
    x"14FF622",
    x"14FF225",
    x"14FEE29",
    x"14FEA2E",
    x"14FE634",
    x"14FE23B",
    x"14FDE43",
    x"14FDA4C",
    x"14FD655",
    x"14FD260",
    x"14FCE6C",
    x"14FCA79",
    x"14FC687",
    x"14FC296",
    x"14FBEA6",
    x"14FBAB7",
    x"14FB6C8",
    x"14FB2DB",
    x"14FAEEF",
    x"14FAB04",
    x"14FA719",
    x"14FA330",
    x"14F9F48",
    x"14F9B61",
    x"14F977A",
    x"14F9395",
    x"14F8FB0",
    x"14F8BCD",
    x"14F87EA",
    x"14F8409",
    x"14F8028",
    x"14F7C49",
    x"14F786A",
    x"14F748D",
    x"14F70B0",
    x"14F6CD4",
    x"14F68FA",
    x"14F6520",
    x"14F6147",
    x"14F5D6F",
    x"14F5998",
    x"14F55C2",
    x"14F51ED",
    x"14F4E19",
    x"14F4A46",
    x"14F4674",
    x"14F42A3",
    x"14F3ED3",
    x"14F3B04",
    x"14F3735",
    x"14F3368",
    x"14F2F9C",
    x"14F2BD0",
    x"14F2806",
    x"14F243C",
    x"14F2074",
    x"14F1CAC",
    x"14F18E5",
    x"14F1520",
    x"14F115B",
    x"14F0D97",
    x"14F09D4",
    x"14F0612",
    x"14F0251",
    x"14EFE91",
    x"14EFAD2",
    x"14EF714",
    x"14EF356",
    x"14EEF9A",
    x"14EEBDE",
    x"14EE824",
    x"14EE46A",
    x"14EE0B2",
    x"14EDCFA",
    x"14ED943",
    x"14ED58D",
    x"14ED1D8",
    x"14ECE24",
    x"14ECA71",
    x"14EC6BF",
    x"14EC30E",
    x"14EBF5E",
    x"14EBBAE",
    x"14EB800",
    x"14EB452",
    x"14EB0A6",
    x"14EACFA",
    x"14EA94F",
    x"14EA5A5",
    x"14EA1FC",
    x"14E9E54",
    x"14E9AAD",
    x"14E9707",
    x"14E9362",
    x"14E8FBD",
    x"14E8C1A",
    x"14E8877",
    x"14E84D6",
    x"14E8135",
    x"14E7D95",
    x"14E79F6",
    x"14E7658",
    x"14E72BB",
    x"14E6F1F",
    x"14E6B83",
    x"14E67E9",
    x"14E644F",
    x"14E60B7",
    x"14E5D1F",
    x"14E5988",
    x"14E55F2",
    x"14E525D",
    x"14E4EC9",
    x"14E4B36",
    x"14E47A3",
    x"14E4412",
    x"14E4081",
    x"14E3CF2",
    x"14E3963",
    x"14E35D5",
    x"14E3248",
    x"14E2EBC",
    x"14E2B31",
    x"14E27A6",
    x"14E241D",
    x"14E2094",
    x"14E1D0D",
    x"14E1986",
    x"14E1600",
    x"14E127B",
    x"14E0EF7",
    x"14E0B73",
    x"14E07F1",
    x"14E046F",
    x"14E00EF",
    x"14DFD6F",
    x"14DF9F0",
    x"14DF672",
    x"14DF2F5",
    x"14DEF78",
    x"14DEBFD",
    x"14DE882",
    x"14DE509",
    x"14DE190",
    x"14DDE18",
    x"14DDAA1",
    x"14DD72B",
    x"14DD3B5",
    x"14DD041",
    x"14DCCCD",
    x"14DC95A",
    x"14DC5E8",
    x"14DC277",
    x"14DBF07",
    x"14DBB98",
    x"14DB829",
    x"14DB4BC",
    x"14DB14F",
    x"14DADE3",
    x"14DAA78",
    x"14DA70E",
    x"14DA3A4",
    x"14DA03C",
    x"14D9CD4",
    x"14D996E",
    x"14D9608",
    x"14D92A3",
    x"14D8F3E",
    x"14D8BDB",
    x"14D8878",
    x"14D8517",
    x"14D81B6",
    x"14D7E56",
    x"14D7AF7",
    x"14D7798",
    x"14D743B",
    x"14D70DE",
    x"14D6D82",
    x"14D6A28",
    x"14D66CD",
    x"14D6374",
    x"14D601C",
    x"14D5CC4",
    x"14D596D",
    x"14D5617",
    x"14D52C2",
    x"14D4F6E",
    x"14D4C1B",
    x"14D48C8",
    x"14D4576",
    x"14D4225",
    x"14D3ED5",
    x"14D3B86",
    x"14D3837",
    x"14D34EA",
    x"14D319D",
    x"14D2E51",
    x"14D2B06",
    x"14D27BB",
    x"14D2472",
    x"14D2129",
    x"14D1DE1",
    x"14D1A9A",
    x"14D1754",
    x"14D140E",
    x"14D10CA",
    x"14D0D86",
    x"14D0A43",
    x"14D0701",
    x"14D03C0",
    x"14D007F",
    x"14CFD3F",
    x"14CFA00",
    x"14CF6C2",
    x"14CF385",
    x"14CF049",
    x"14CED0D",
    x"14CE9D2",
    x"14CE698",
    x"14CE35F",
    x"14CE026",
    x"14CDCEF",
    x"14CD9B8",
    x"14CD682",
    x"14CD34D",
    x"14CD018",
    x"14CCCE5",
    x"14CC9B2",
    x"14CC680",
    x"14CC34E",
    x"14CC01E",
    x"14CBCEE",
    x"14CB9C0",
    x"14CB692",
    x"14CB364",
    x"14CB038",
    x"14CAD0C",
    x"14CA9E1",
    x"14CA6B7",
    x"14CA38E",
    x"14CA065",
    x"14C9D3E",
    x"14C9A17",
    x"14C96F1",
    x"14C93CB",
    x"14C90A7",
    x"14C8D83",
    x"14C8A60",
    x"14C873E",
    x"14C841C",
    x"14C80FC",
    x"14C7DDC",
    x"14C7ABD",
    x"14C779F",
    x"14C7481",
    x"14C7164",
    x"14C6E48",
    x"14C6B2D",
    x"14C6813",
    x"14C64F9",
    x"14C61E0",
    x"14C5EC8",
    x"14C5BB1",
    x"14C589A",
    x"14C5585",
    x"14C5270",
    x"14C4F5B",
    x"14C4C48",
    x"14C4935",
    x"14C4623",
    x"14C4312",
    x"14C4002",
    x"14C3CF2",
    x"14C39E3",
    x"14C36D5",
    x"14C33C8",
    x"14C30BB",
    x"14C2DB0",
    x"14C2AA4",
    x"14C279A",
    x"14C2491",
    x"14C2188",
    x"14C1E80",
    x"14C1B79",
    x"14C1872",
    x"14C156C",
    x"14C1267",
    x"14C0F63",
    x"14C0C60",
    x"14C095D",
    x"14C065B",
    x"14C035A",
    x"14C0059",
    x"14BFD5A",
    x"14BFA5B",
    x"14BF75D",
    x"14BF45F",
    x"14BF162",
    x"14BEE66",
    x"14BEB6B",
    x"14BE871",
    x"14BE577",
    x"14BE27E",
    x"14BDF86",
    x"14BDC8E",
    x"14BD997",
    x"14BD6A1",
    x"14BD3AC",
    x"14BD0B8",
    x"14BCDC4",
    x"14BCAD1",
    x"14BC7DE",
    x"14BC4ED",
    x"14BC1FC",
    x"14BBF0C",
    x"14BBC1C",
    x"14BB92E",
    x"14BB640",
    x"14BB353",
    x"14BB066",
    x"14BAD7A",
    x"14BAA8F",
    x"14BA7A5",
    x"14BA4BC",
    x"14BA1D3",
    x"14B9EEB",
    x"14B9C03",
    x"14B991D",
    x"14B9637",
    x"14B9351",
    x"14B906D",
    x"14B8D89",
    x"14B8AA6",
    x"14B87C4",
    x"14B84E2",
    x"14B8201",
    x"14B7F21",
    x"14B7C42",
    x"14B7963",
    x"14B7685",
    x"14B73A8",
    x"14B70CB",
    x"14B6DF0",
    x"14B6B14",
    x"14B683A",
    x"14B6560",
    x"14B6287",
    x"14B5FAF",
    x"14B5CD7",
    x"14B5A01",
    x"14B572A",
    x"14B5455",
    x"14B5180",
    x"14B4EAC",
    x"14B4BD9",
    x"14B4906",
    x"14B4634",
    x"14B4363",
    x"14B4093",
    x"14B3DC3",
    x"14B3AF4",
    x"14B3826",
    x"14B3558",
    x"14B328B",
    x"14B2FBF",
    x"14B2CF3",
    x"14B2A28",
    x"14B275E",
    x"14B2494",
    x"14B21CC",
    x"14B1F03",
    x"14B1C3C",
    x"14B1975",
    x"14B16AF",
    x"14B13EA",
    x"14B1125",
    x"14B0E61",
    x"14B0B9E",
    x"14B08DC",
    x"14B061A",
    x"14B0359",
    x"14B0098",
    x"14AFDD8",
    x"14AFB19",
    x"14AF85B",
    x"14AF59D",
    x"14AF2E0",
    x"14AF024",
    x"14AED68",
    x"14AEAAD",
    x"14AE7F3",
    x"14AE539",
    x"14AE280",
    x"14ADFC8",
    x"14ADD10",
    x"14ADA59",
    x"14AD7A3",
    x"14AD4ED",
    x"14AD238",
    x"14ACF84",
    x"14ACCD1",
    x"14ACA1E",
    x"14AC76C",
    x"14AC4BA",
    x"14AC209",
    x"14ABF59",
    x"14ABCAA",
    x"14AB9FB",
    x"14AB74D",
    x"14AB49F",
    x"14AB1F2",
    x"14AAF46",
    x"14AAC9B",
    x"14AA9F0",
    x"14AA746",
    x"14AA49C",
    x"14AA1F3",
    x"14A9F4B",
    x"14A9CA4",
    x"14A99FD",
    x"14A9757",
    x"14A94B1",
    x"14A920C",
    x"14A8F68",
    x"14A8CC5",
    x"14A8A22",
    x"14A8780",
    x"14A84DE",
    x"14A823D",
    x"14A7F9D",
    x"14A7CFD",
    x"14A7A5E",
    x"14A77C0",
    x"14A7523",
    x"14A7286",
    x"14A6FE9",
    x"14A6D4E",
    x"14A6AB3",
    x"14A6818",
    x"14A657F",
    x"14A62E5",
    x"14A604D",
    x"14A5DB5",
    x"14A5B1E",
    x"14A5888",
    x"14A55F2",
    x"14A535D",
    x"14A50C8",
    x"14A4E34",
    x"14A4BA1",
    x"14A490F",
    x"14A467D",
    x"14A43EB",
    x"14A415B",
    x"14A3ECB",
    x"14A3C3B",
    x"14A39AD",
    x"14A371E",
    x"14A3491",
    x"14A3204",
    x"14A2F78",
    x"14A2CEC",
    x"14A2A62",
    x"14A27D7",
    x"14A254E",
    x"14A22C5",
    x"14A203C",
    x"14A1DB4",
    x"14A1B2D",
    x"14A18A7",
    x"14A1621",
    x"14A139C",
    x"14A1117",
    x"14A0E93",
    x"14A0C10",
    x"14A098D",
    x"14A070B",
    x"14A048A",
    x"14A0209",
    x"149FF89",
    x"149FD09",
    x"149FA8A",
    x"149F80C",
    x"149F58E",
    x"149F311",
    x"149F095",
    x"149EE19",
    x"149EB9E",
    x"149E923",
    x"149E6A9",
    x"149E430",
    x"149E1B7",
    x"149DF3F",
    x"149DCC7",
    x"149DA50",
    x"149D7DA",
    x"149D564",
    x"149D2EF",
    x"149D07B",
    x"149CE07",
    x"149CB94",
    x"149C921",
    x"149C6AF",
    x"149C43E",
    x"149C1CD",
    x"149BF5D",
    x"149BCEE",
    x"149BA7F",
    x"149B810",
    x"149B5A3",
    x"149B336",
    x"149B0C9",
    x"149AE5D",
    x"149ABF2",
    x"149A987",
    x"149A71D",
    x"149A4B4",
    x"149A24B",
    x"1499FE2",
    x"1499D7B",
    x"1499B14",
    x"14998AD",
    x"1499647",
    x"14993E2",
    x"149917D",
    x"1498F19",
    x"1498CB6",
    x"1498A53",
    x"14987F1",
    x"149858F",
    x"149832E",
    x"14980CD",
    x"1497E6E",
    x"1497C0E",
    x"14979B0",
    x"1497751",
    x"14974F4",
    x"1497297",
    x"149703B",
    x"1496DDF",
    x"1496B84",
    x"1496929",
    x"14966CF",
    x"1496476",
    x"149621D",
    x"1495FC5",
    x"1495D6D",
    x"1495B16",
    x"14958BF",
    x"149566A",
    x"1495414",
    x"14951BF",
    x"1494F6B",
    x"1494D18",
    x"1494AC5",
    x"1494872",
    x"1494621",
    x"14943CF",
    x"149417F",
    x"1493F2F",
    x"1493CDF",
    x"1493A90",
    x"1493842",
    x"14935F4",
    x"14933A7",
    x"149315A",
    x"1492F0E",
    x"1492CC3",
    x"1492A78",
    x"149282D",
    x"14925E4",
    x"149239A",
    x"1492152",
    x"1491F0A",
    x"1491CC2",
    x"1491A7B",
    x"1491835",
    x"14915EF",
    x"14913AA",
    x"1491165",
    x"1490F21",
    x"1490CDE",
    x"1490A9B",
    x"1490859",
    x"1490617",
    x"14903D6",
    x"1490195",
    x"148FF55",
    x"148FD15",
    x"148FAD6",
    x"148F898",
    x"148F65A",
    x"148F41D",
    x"148F1E0",
    x"148EFA4",
    x"148ED68",
    x"148EB2D",
    x"148E8F2",
    x"148E6B8",
    x"148E47F",
    x"148E246",
    x"148E00E",
    x"148DDD6",
    x"148DB9F",
    x"148D968",
    x"148D732",
    x"148D4FD",
    x"148D2C8",
    x"148D093",
    x"148CE60",
    x"148CC2C",
    x"148C9F9",
    x"148C7C7",
    x"148C596",
    x"148C364",
    x"148C134",
    x"148BF04",
    x"148BCD4",
    x"148BAA5",
    x"148B877",
    x"148B649",
    x"148B41C",
    x"148B1EF",
    x"148AFC3",
    x"148AD97",
    x"148AB6C",
    x"148A942",
    x"148A718",
    x"148A4EE",
    x"148A2C5",
    x"148A09D",
    x"1489E75",
    x"1489C4D",
    x"1489A27",
    x"1489800",
    x"14895DB",
    x"14893B5",
    x"1489191",
    x"1488F6D",
    x"1488D49",
    x"1488B26",
    x"1488903",
    x"14886E1",
    x"14884C0",
    x"148829F",
    x"148807F",
    x"1487E5F",
    x"1487C3F",
    x"1487A21",
    x"1487802",
    x"14875E5",
    x"14873C7",
    x"14871AB",
    x"1486F8F",
    x"1486D73",
    x"1486B58",
    x"148693D",
    x"1486723",
    x"148650A",
    x"14862F1",
    x"14860D8",
    x"1485EC0",
    x"1485CA9",
    x"1485A92",
    x"148587C",
    x"1485666",
    x"1485450",
    x"148523C",
    x"1485027",
    x"1484E14",
    x"1484C00",
    x"14849EE",
    x"14847DB",
    x"14845CA",
    x"14843B8",
    x"14841A8",
    x"1483F98",
    x"1483D88",
    x"1483B79",
    x"148396A",
    x"148375C",
    x"148354F",
    x"1483341",
    x"1483135",
    x"1482F29",
    x"1482D1D",
    x"1482B12",
    x"1482908",
    x"14826FE",
    x"14824F4",
    x"14822EB",
    x"14820E3",
    x"1481EDB",
    x"1481CD3",
    x"1481ACC",
    x"14818C6",
    x"14816C0",
    x"14814BB",
    x"14812B6",
    x"14810B1",
    x"1480EAD",
    x"1480CAA",
    x"1480AA7",
    x"14808A5",
    x"14806A3",
    x"14804A1",
    x"14802A0",
    x"14800A0",
    x"147FD41",
    x"147F942",
    x"147F544",
    x"147F147",
    x"147ED4B",
    x"147E950",
    x"147E557",
    x"147E15E",
    x"147DD66",
    x"147D96F",
    x"147D579",
    x"147D184",
    x"147CD91",
    x"147C99E",
    x"147C5AC",
    x"147C1BB",
    x"147BDCB",
    x"147B9DC",
    x"147B5EE",
    x"147B201",
    x"147AE15",
    x"147AA2A",
    x"147A640",
    x"147A257",
    x"1479E6F",
    x"1479A88",
    x"14796A1",
    x"14792BC",
    x"1478ED8",
    x"1478AF5",
    x"1478713",
    x"1478331",
    x"1477F51",
    x"1477B72",
    x"1477793",
    x"14773B6",
    x"1476FD9",
    x"1476BFE",
    x"1476823",
    x"147644A",
    x"1476071",
    x"1475C9A",
    x"14758C3",
    x"14754ED",
    x"1475118",
    x"1474D45",
    x"1474972",
    x"14745A0",
    x"14741CF",
    x"1473DFF",
    x"1473A30",
    x"1473662",
    x"1473295",
    x"1472EC9",
    x"1472AFD",
    x"1472733",
    x"147236A",
    x"1471FA1",
    x"1471BDA",
    x"1471814",
    x"147144E",
    x"1471089",
    x"1470CC6",
    x"1470903",
    x"1470541",
    x"1470180",
    x"146FDC0",
    x"146FA01",
    x"146F643",
    x"146F286",
    x"146EECA",
    x"146EB0F",
    x"146E755",
    x"146E39B",
    x"146DFE3",
    x"146DC2B",
    x"146D875",
    x"146D4BF",
    x"146D10A",
    x"146CD57",
    x"146C9A4",
    x"146C5F2",
    x"146C241",
    x"146BE91",
    x"146BAE1",
    x"146B733",
    x"146B386",
    x"146AFD9",
    x"146AC2E",
    x"146A883",
    x"146A4DA",
    x"146A131",
    x"1469D89",
    x"14699E2",
    x"146963C",
    x"1469297",
    x"1468EF3",
    x"1468B50",
    x"14687AD",
    x"146840C",
    x"146806B",
    x"1467CCB",
    x"146792D",
    x"146758F",
    x"14671F2",
    x"1466E56",
    x"1466ABB",
    x"1466721",
    x"1466387",
    x"1465FEF",
    x"1465C57",
    x"14658C1",
    x"146552B",
    x"1465196",
    x"1464E02",
    x"1464A6F",
    x"14646DD",
    x"146434C",
    x"1463FBB",
    x"1463C2C",
    x"146389D",
    x"146350F",
    x"1463183",
    x"1462DF7",
    x"1462A6C",
    x"14626E1",
    x"1462358",
    x"1461FD0",
    x"1461C48",
    x"14618C2",
    x"146153C",
    x"14611B7",
    x"1460E33",
    x"1460AB0",
    x"146072E",
    x"14603AC",
    x"146002C",
    x"145FCAC",
    x"145F92E",
    x"145F5B0",
    x"145F233",
    x"145EEB7",
    x"145EB3B",
    x"145E7C1",
    x"145E447",
    x"145E0CF",
    x"145DD57",
    x"145D9E0",
    x"145D66A",
    x"145D2F5",
    x"145CF81",
    x"145CC0D",
    x"145C89B",
    x"145C529",
    x"145C1B8",
    x"145BE48",
    x"145BAD9",
    x"145B76B",
    x"145B3FD",
    x"145B091",
    x"145AD25",
    x"145A9BA",
    x"145A650",
    x"145A2E7",
    x"1459F7F",
    x"1459C17",
    x"14598B0",
    x"145954B",
    x"14591E6",
    x"1458E82",
    x"1458B1F",
    x"14587BC",
    x"145845B",
    x"14580FA",
    x"1457D9A",
    x"1457A3B",
    x"14576DD",
    x"1457380",
    x"1457023",
    x"1456CC8",
    x"145696D",
    x"1456613",
    x"14562BA",
    x"1455F62",
    x"1455C0A",
    x"14558B4",
    x"145555E",
    x"1455209",
    x"1454EB5",
    x"1454B62",
    x"145480F",
    x"14544BE",
    x"145416D",
    x"1453E1D",
    x"1453ACE",
    x"145377F",
    x"1453432",
    x"14530E5",
    x"1452D9A",
    x"1452A4F",
    x"1452704",
    x"14523BB",
    x"1452073",
    x"1451D2B",
    x"14519E4",
    x"145169E",
    x"1451359",
    x"1451014",
    x"1450CD1",
    x"145098E",
    x"145064C",
    x"145030B",
    x"144FFCA",
    x"144FC8B",
    x"144F94C",
    x"144F60E",
    x"144F2D1",
    x"144EF95",
    x"144EC59",
    x"144E91F",
    x"144E5E5",
    x"144E2AC",
    x"144DF73",
    x"144DC3C",
    x"144D905",
    x"144D5CF",
    x"144D29A",
    x"144CF66",
    x"144CC33",
    x"144C900",
    x"144C5CE",
    x"144C29D",
    x"144BF6D",
    x"144BC3D",
    x"144B90F",
    x"144B5E1",
    x"144B2B4",
    x"144AF87",
    x"144AC5C",
    x"144A931",
    x"144A607",
    x"144A2DE",
    x"1449FB6",
    x"1449C8E",
    x"1449968",
    x"1449642",
    x"144931D",
    x"1448FF8",
    x"1448CD5",
    x"14489B2",
    x"1448690",
    x"144836E",
    x"144804E",
    x"1447D2E",
    x"1447A0F",
    x"14476F1",
    x"14473D4",
    x"14470B7",
    x"1446D9C",
    x"1446A81",
    x"1446766",
    x"144644D",
    x"1446134",
    x"1445E1C",
    x"1445B05",
    x"14457EF",
    x"14454D9",
    x"14451C4",
    x"1444EB0",
    x"1444B9D",
    x"144488A",
    x"1444579",
    x"1444268",
    x"1443F57",
    x"1443C48",
    x"1443939",
    x"144362B",
    x"144331E",
    x"1443012",
    x"1442D06",
    x"14429FB",
    x"14426F1",
    x"14423E8",
    x"14420DF",
    x"1441DD7",
    x"1441AD0",
    x"14417CA",
    x"14414C4",
    x"14411C0",
    x"1440EBC",
    x"1440BB8",
    x"14408B6",
    x"14405B4",
    x"14402B3",
    x"143FFB3",
    x"143FCB3",
    x"143F9B4",
    x"143F6B6",
    x"143F3B9",
    x"143F0BC",
    x"143EDC0",
    x"143EAC5",
    x"143E7CB",
    x"143E4D2",
    x"143E1D9",
    x"143DEE1",
    x"143DBE9",
    x"143D8F3",
    x"143D5FD",
    x"143D308",
    x"143D013",
    x"143CD20",
    x"143CA2D",
    x"143C73B",
    x"143C449",
    x"143C158",
    x"143BE68",
    x"143BB79",
    x"143B88B",
    x"143B59D",
    x"143B2B0",
    x"143AFC4",
    x"143ACD8",
    x"143A9ED",
    x"143A703",
    x"143A41A",
    x"143A131",
    x"1439E49",
    x"1439B62",
    x"143987B",
    x"1439596",
    x"14392B1",
    x"1438FCC",
    x"1438CE9",
    x"1438A06",
    x"1438724",
    x"1438442",
    x"1438161",
    x"1437E81",
    x"1437BA2",
    x"14378C4",
    x"14375E6",
    x"1437309",
    x"143702C",
    x"1436D51",
    x"1436A76",
    x"143679B",
    x"14364C2",
    x"14361E9",
    x"1435F11",
    x"1435C39",
    x"1435963",
    x"143568D",
    x"14353B8",
    x"14350E3",
    x"1434E0F",
    x"1434B3C",
    x"1434869",
    x"1434598",
    x"14342C7",
    x"1433FF6",
    x"1433D27",
    x"1433A58",
    x"143378A",
    x"14334BC",
    x"14331EF",
    x"1432F23",
    x"1432C58",
    x"143298D",
    x"14326C3",
    x"14323F9",
    x"1432131",
    x"1431E69",
    x"1431BA2",
    x"14318DB",
    x"1431615",
    x"1431350",
    x"143108C",
    x"1430DC8",
    x"1430B05",
    x"1430842",
    x"1430580",
    x"14302BF",
    x"142FFFF",
    x"142FD3F",
    x"142FA80",
    x"142F7C2",
    x"142F505",
    x"142F248",
    x"142EF8B",
    x"142ECD0",
    x"142EA15",
    x"142E75B",
    x"142E4A1",
    x"142E1E9",
    x"142DF30",
    x"142DC79",
    x"142D9C2",
    x"142D70C",
    x"142D457",
    x"142D1A2",
    x"142CEEE",
    x"142CC3A",
    x"142C988",
    x"142C6D6",
    x"142C424",
    x"142C174",
    x"142BEC4",
    x"142BC14",
    x"142B966",
    x"142B6B8",
    x"142B40A",
    x"142B15E",
    x"142AEB1",
    x"142AC06",
    x"142A95B",
    x"142A6B1",
    x"142A408",
    x"142A15F",
    x"1429EB7",
    x"1429C10",
    x"1429969",
    x"14296C3",
    x"142941E",
    x"1429179",
    x"1428ED5",
    x"1428C32",
    x"142898F",
    x"14286ED",
    x"142844C",
    x"14281AB",
    x"1427F0B",
    x"1427C6B",
    x"14279CD",
    x"142772F",
    x"1427491",
    x"14271F4",
    x"1426F58",
    x"1426CBD",
    x"1426A22",
    x"1426788",
    x"14264EE",
    x"1426255",
    x"1425FBD",
    x"1425D25",
    x"1425A8E",
    x"14257F8",
    x"1425562",
    x"14252CD",
    x"1425039",
    x"1424DA5",
    x"1424B12",
    x"1424880",
    x"14245EE",
    x"142435D",
    x"14240CC",
    x"1423E3C",
    x"1423BAD",
    x"142391E",
    x"1423690",
    x"1423403",
    x"1423176",
    x"1422EEA",
    x"1422C5F",
    x"14229D4",
    x"142274A",
    x"14224C1",
    x"1422238",
    x"1421FAF",
    x"1421D28",
    x"1421AA1",
    x"142181A",
    x"1421595",
    x"1421310",
    x"142108B",
    x"1420E07",
    x"1420B84",
    x"1420902",
    x"1420680",
    x"14203FE",
    x"142017E",
    x"141FEFE",
    x"141FC7E",
    x"141F9FF",
    x"141F781",
    x"141F504",
    x"141F287",
    x"141F00A",
    x"141ED8F",
    x"141EB14",
    x"141E899",
    x"141E61F",
    x"141E3A6",
    x"141E12E",
    x"141DEB6",
    x"141DC3E",
    x"141D9C7",
    x"141D751",
    x"141D4DC",
    x"141D267",
    x"141CFF3",
    x"141CD7F",
    x"141CB0C",
    x"141C899",
    x"141C627",
    x"141C3B6",
    x"141C146",
    x"141BED6",
    x"141BC66",
    x"141B9F7",
    x"141B789",
    x"141B51C",
    x"141B2AF",
    x"141B042",
    x"141ADD7",
    x"141AB6B",
    x"141A901",
    x"141A697",
    x"141A42E",
    x"141A1C5",
    x"1419F5D",
    x"1419CF5",
    x"1419A8E",
    x"1419828",
    x"14195C2",
    x"141935D",
    x"14190F8",
    x"1418E94",
    x"1418C31",
    x"14189CE",
    x"141876C",
    x"141850B",
    x"14182AA",
    x"1418049",
    x"1417DEA",
    x"1417B8A",
    x"141792C",
    x"14176CE",
    x"1417470",
    x"1417214",
    x"1416FB7",
    x"1416D5C",
    x"1416B01",
    x"14168A6",
    x"141664C",
    x"14163F3",
    x"141619A",
    x"1415F42",
    x"1415CEB",
    x"1415A94",
    x"141583D",
    x"14155E8",
    x"1415392",
    x"141513E",
    x"1414EEA",
    x"1414C96",
    x"1414A44",
    x"14147F1",
    x"14145A0",
    x"141434E",
    x"14140FE",
    x"1413EAE",
    x"1413C5F",
    x"1413A10",
    x"14137C2",
    x"1413574",
    x"1413327",
    x"14130DA",
    x"1412E8E",
    x"1412C43",
    x"14129F8",
    x"14127AE",
    x"1412564",
    x"141231B",
    x"14120D3",
    x"1411E8B",
    x"1411C44",
    x"14119FD",
    x"14117B7",
    x"1411571",
    x"141132C",
    x"14110E7",
    x"1410EA3",
    x"1410C60",
    x"1410A1D",
    x"14107DB",
    x"1410599",
    x"1410358",
    x"1410118",
    x"140FED8",
    x"140FC98",
    x"140FA59",
    x"140F81B",
    x"140F5DD",
    x"140F3A0",
    x"140F163",
    x"140EF27",
    x"140ECEC",
    x"140EAB1",
    x"140E877",
    x"140E63D",
    x"140E403",
    x"140E1CB",
    x"140DF93",
    x"140DD5B",
    x"140DB24",
    x"140D8ED",
    x"140D6B7",
    x"140D482",
    x"140D24D",
    x"140D019",
    x"140CDE5",
    x"140CBB2",
    x"140C97F",
    x"140C74D",
    x"140C51C",
    x"140C2EB",
    x"140C0BA",
    x"140BE8A",
    x"140BC5B",
    x"140BA2C",
    x"140B7FE",
    x"140B5D0",
    x"140B3A3",
    x"140B176",
    x"140AF4A",
    x"140AD1F",
    x"140AAF4",
    x"140A8C9",
    x"140A69F",
    x"140A476",
    x"140A24D",
    x"140A025",
    x"1409DFD",
    x"1409BD6",
    x"14099AF",
    x"1409789",
    x"1409563",
    x"140933E",
    x"140911A",
    x"1408EF6",
    x"1408CD2",
    x"1408AAF",
    x"140888D",
    x"140866B",
    x"140844A",
    x"1408229",
    x"1408008",
    x"1407DE9",
    x"1407BCA",
    x"14079AB",
    x"140778D",
    x"140756F",
    x"1407352",
    x"1407135",
    x"1406F19",
    x"1406CFE",
    x"1406AE3",
    x"14068C8",
    x"14066AE",
    x"1406495",
    x"140627C",
    x"1406064",
    x"1405E4C",
    x"1405C35",
    x"1405A1E",
    x"1405808",
    x"14055F2",
    x"14053DD",
    x"14051C8",
    x"1404FB4",
    x"1404DA0",
    x"1404B8D",
    x"140497A",
    x"1404768",
    x"1404557",
    x"1404346",
    x"1404135",
    x"1403F25",
    x"1403D15",
    x"1403B06",
    x"14038F8",
    x"14036EA",
    x"14034DC",
    x"14032CF",
    x"14030C3",
    x"1402EB7",
    x"1402CAC",
    x"1402AA1",
    x"1402896",
    x"140268C",
    x"1402483",
    x"140227A",
    x"1402072",
    x"1401E6A",
    x"1401C63",
    x"1401A5C",
    x"1401855",
    x"1401650",
    x"140144A",
    x"1401245",
    x"1401041",
    x"1400E3D",
    x"1400C3A",
    x"1400A37",
    x"1400835",
    x"1400633",
    x"1400432",
    x"1400231",
    x"1400031",
    x"13FFC62",
    x"13FF864",
    x"13FF466",
    x"13FF069",
    x"13FEC6E",
    x"13FE873",
    x"13FE47A",
    x"13FE081",
    x"13FDC89",
    x"13FD893",
    x"13FD49D",
    x"13FD0A8",
    x"13FCCB5",
    x"13FC8C2",
    x"13FC4D0",
    x"13FC0E0",
    x"13FBCF0",
    x"13FB901",
    x"13FB513",
    x"13FB127",
    x"13FAD3B",
    x"13FA950",
    x"13FA566",
    x"13FA17D",
    x"13F9D95",
    x"13F99AF",
    x"13F95C9",
    x"13F91E4",
    x"13F8E00",
    x"13F8A1D",
    x"13F863B",
    x"13F825A",
    x"13F7E79",
    x"13F7A9A",
    x"13F76BC",
    x"13F72DF",
    x"13F6F03",
    x"13F6B27",
    x"13F674D",
    x"13F6374",
    x"13F5F9B",
    x"13F5BC4",
    x"13F57EE",
    x"13F5418",
    x"13F5043",
    x"13F4C70",
    x"13F489D",
    x"13F44CC",
    x"13F40FB",
    x"13F3D2B",
    x"13F395C",
    x"13F358E",
    x"13F31C1",
    x"13F2DF6",
    x"13F2A2B",
    x"13F2660",
    x"13F2297",
    x"13F1ECF",
    x"13F1B08",
    x"13F1742",
    x"13F137C",
    x"13F0FB8",
    x"13F0BF4",
    x"13F0832",
    x"13F0470",
    x"13F00B0",
    x"13EFCF0",
    x"13EF931",
    x"13EF573",
    x"13EF1B6",
    x"13EEDFB",
    x"13EEA3F",
    x"13EE685",
    x"13EE2CC",
    x"13EDF14",
    x"13EDB5D",
    x"13ED7A6",
    x"13ED3F1",
    x"13ED03C",
    x"13ECC89",
    x"13EC8D6",
    x"13EC524",
    x"13EC173",
    x"13EBDC4",
    x"13EBA15",
    x"13EB667",
    x"13EB2B9",
    x"13EAF0D",
    x"13EAB62",
    x"13EA7B7",
    x"13EA40E",
    x"13EA065",
    x"13E9CBE",
    x"13E9917",
    x"13E9571",
    x"13E91CC",
    x"13E8E28",
    x"13E8A85",
    x"13E86E3",
    x"13E8342",
    x"13E7FA1",
    x"13E7C02",
    x"13E7863",
    x"13E74C6",
    x"13E7129",
    x"13E6D8D",
    x"13E69F2",
    x"13E6658",
    x"13E62BF",
    x"13E5F27",
    x"13E5B90",
    x"13E57F9",
    x"13E5464",
    x"13E50CF",
    x"13E4D3B",
    x"13E49A8",
    x"13E4616",
    x"13E4285",
    x"13E3EF5",
    x"13E3B66",
    x"13E37D7",
    x"13E344A",
    x"13E30BD",
    x"13E2D31",
    x"13E29A7",
    x"13E261D",
    x"13E2294",
    x"13E1F0B",
    x"13E1B84",
    x"13E17FE",
    x"13E1478",
    x"13E10F3",
    x"13E0D70",
    x"13E09ED",
    x"13E066B",
    x"13E02E9",
    x"13DFF69",
    x"13DFBEA",
    x"13DF86B",
    x"13DF4EE",
    x"13DF171",
    x"13DEDF5",
    x"13DEA7A",
    x"13DE700",
    x"13DE386",
    x"13DE00E",
    x"13DDC96",
    x"13DD920",
    x"13DD5AA",
    x"13DD235",
    x"13DCEC1",
    x"13DCB4D",
    x"13DC7DB",
    x"13DC469",
    x"13DC0F9",
    x"13DBD89",
    x"13DBA1A",
    x"13DB6AC",
    x"13DB33F",
    x"13DAFD2",
    x"13DAC67",
    x"13DA8FC",
    x"13DA592",
    x"13DA229",
    x"13D9EC1",
    x"13D9B5A",
    x"13D97F3",
    x"13D948E",
    x"13D9129",
    x"13D8DC5",
    x"13D8A62",
    x"13D8700",
    x"13D839F",
    x"13D803E",
    x"13D7CDF",
    x"13D7980",
    x"13D7622",
    x"13D72C5",
    x"13D6F69",
    x"13D6C0D",
    x"13D68B2",
    x"13D6559",
    x"13D6200",
    x"13D5EA8",
    x"13D5B50",
    x"13D57FA",
    x"13D54A4",
    x"13D5150",
    x"13D4DFC",
    x"13D4AA9",
    x"13D4757",
    x"13D4405",
    x"13D40B4",
    x"13D3D65",
    x"13D3A16",
    x"13D36C8",
    x"13D337A",
    x"13D302E",
    x"13D2CE2",
    x"13D2998",
    x"13D264E",
    x"13D2304",
    x"13D1FBC",
    x"13D1C74",
    x"13D192E",
    x"13D15E8",
    x"13D12A3",
    x"13D0F5F",
    x"13D0C1B",
    x"13D08D9",
    x"13D0597",
    x"13D0256",
    x"13CFF16",
    x"13CFBD6",
    x"13CF898",
    x"13CF55A",
    x"13CF21D",
    x"13CEEE1",
    x"13CEBA6",
    x"13CE86B",
    x"13CE531",
    x"13CE1F8",
    x"13CDEC0",
    x"13CDB89",
    x"13CD853",
    x"13CD51D",
    x"13CD1E8",
    x"13CCEB4",
    x"13CCB81",
    x"13CC84E",
    x"13CC51C",
    x"13CC1EC",
    x"13CBEBC",
    x"13CBB8C",
    x"13CB85E",
    x"13CB530",
    x"13CB203",
    x"13CAED7",
    x"13CABAC",
    x"13CA881",
    x"13CA557",
    x"13CA22F",
    x"13C9F06",
    x"13C9BDF",
    x"13C98B8",
    x"13C9593",
    x"13C926E",
    x"13C8F49",
    x"13C8C26",
    x"13C8903",
    x"13C85E2",
    x"13C82C0",
    x"13C7FA0",
    x"13C7C81",
    x"13C7962",
    x"13C7644",
    x"13C7327",
    x"13C700A",
    x"13C6CEF",
    x"13C69D4",
    x"13C66BA",
    x"13C63A1",
    x"13C6088",
    x"13C5D70",
    x"13C5A59",
    x"13C5743",
    x"13C542E",
    x"13C5119",
    x"13C4E05",
    x"13C4AF2",
    x"13C47E0",
    x"13C44CE",
    x"13C41BD",
    x"13C3EAD",
    x"13C3B9E",
    x"13C388F",
    x"13C3582",
    x"13C3275",
    x"13C2F68",
    x"13C2C5D",
    x"13C2952",
    x"13C2648",
    x"13C233F",
    x"13C2037",
    x"13C1D2F",
    x"13C1A28",
    x"13C1722",
    x"13C141C",
    x"13C1118",
    x"13C0E14",
    x"13C0B11",
    x"13C080E",
    x"13C050D",
    x"13C020C",
    x"13BFF0C",
    x"13BFC0C",
    x"13BF90E",
    x"13BF610",
    x"13BF313",
    x"13BF016",
    x"13BED1B",
    x"13BEA20",
    x"13BE726",
    x"13BE42C",
    x"13BE133",
    x"13BDE3C",
    x"13BDB44",
    x"13BD84E",
    x"13BD558",
    x"13BD263",
    x"13BCF6F",
    x"13BCC7B",
    x"13BC989",
    x"13BC697",
    x"13BC3A5",
    x"13BC0B5",
    x"13BBDC5",
    x"13BBAD6",
    x"13BB7E8",
    x"13BB4FA",
    x"13BB20D",
    x"13BAF21",
    x"13BAC36",
    x"13BA94B",
    x"13BA661",
    x"13BA378",
    x"13BA08F",
    x"13B9DA7",
    x"13B9AC0",
    x"13B97DA",
    x"13B94F4",
    x"13B9210",
    x"13B8F2B",
    x"13B8C48",
    x"13B8965",
    x"13B8683",
    x"13B83A2",
    x"13B80C1",
    x"13B7DE2",
    x"13B7B03",
    x"13B7824",
    x"13B7546",
    x"13B726A",
    x"13B6F8D",
    x"13B6CB2",
    x"13B69D7",
    x"13B66FD",
    x"13B6423",
    x"13B614B",
    x"13B5E73",
    x"13B5B9C",
    x"13B58C5",
    x"13B55EF",
    x"13B531A",
    x"13B5046",
    x"13B4D72",
    x"13B4A9F",
    x"13B47CD",
    x"13B44FB",
    x"13B422A",
    x"13B3F5A",
    x"13B3C8A",
    x"13B39BC",
    x"13B36EE",
    x"13B3420",
    x"13B3153",
    x"13B2E87",
    x"13B2BBC",
    x"13B28F2",
    x"13B2628",
    x"13B235F",
    x"13B2096",
    x"13B1DCE",
    x"13B1B07",
    x"13B1841",
    x"13B157B",
    x"13B12B6",
    x"13B0FF2",
    x"13B0D2E",
    x"13B0A6B",
    x"13B07A9",
    x"13B04E7",
    x"13B0226",
    x"13AFF66",
    x"13AFCA7",
    x"13AF9E8",
    x"13AF72A",
    x"13AF46C",
    x"13AF1AF",
    x"13AEEF3",
    x"13AEC38",
    x"13AE97D",
    x"13AE6C3",
    x"13AE40A",
    x"13AE151",
    x"13ADE99",
    x"13ADBE2",
    x"13AD92B",
    x"13AD675",
    x"13AD3C0",
    x"13AD10B",
    x"13ACE58",
    x"13ACBA4",
    x"13AC8F2",
    x"13AC640",
    x"13AC38F",
    x"13AC0DE",
    x"13ABE2E",
    x"13ABB7F",
    x"13AB8D0",
    x"13AB623",
    x"13AB375",
    x"13AB0C9",
    x"13AAE1D",
    x"13AAB72",
    x"13AA8C7",
    x"13AA61D",
    x"13AA374",
    x"13AA0CC",
    x"13A9E24",
    x"13A9B7D",
    x"13A98D6",
    x"13A9630",
    x"13A938B",
    x"13A90E6",
    x"13A8E42",
    x"13A8B9F",
    x"13A88FD",
    x"13A865B",
    x"13A83B9",
    x"13A8119",
    x"13A7E79",
    x"13A7BDA",
    x"13A793B",
    x"13A769D",
    x"13A7400",
    x"13A7163",
    x"13A6EC7",
    x"13A6C2C",
    x"13A6991",
    x"13A66F7",
    x"13A645D",
    x"13A61C5",
    x"13A5F2D",
    x"13A5C95",
    x"13A59FE",
    x"13A5768",
    x"13A54D3",
    x"13A523E",
    x"13A4FA9",
    x"13A4D16",
    x"13A4A83",
    x"13A47F1",
    x"13A455F",
    x"13A42CE",
    x"13A403E",
    x"13A3DAE",
    x"13A3B1F",
    x"13A3890",
    x"13A3602",
    x"13A3375",
    x"13A30E9",
    x"13A2E5D",
    x"13A2BD1",
    x"13A2947",
    x"13A26BD",
    x"13A2433",
    x"13A21AB",
    x"13A1F23",
    x"13A1C9B",
    x"13A1A14",
    x"13A178E",
    x"13A1509",
    x"13A1284",
    x"13A0FFF",
    x"13A0D7C",
    x"13A0AF9",
    x"13A0876",
    x"13A05F4",
    x"13A0373",
    x"13A00F3",
    x"139FE73",
    x"139FBF3",
    x"139F975",
    x"139F6F7",
    x"139F479",
    x"139F1FC",
    x"139EF80",
    x"139ED05",
    x"139EA8A",
    x"139E80F",
    x"139E596",
    x"139E31D",
    x"139E0A4",
    x"139DE2C",
    x"139DBB5",
    x"139D93E",
    x"139D6C8",
    x"139D453",
    x"139D1DE",
    x"139CF6A",
    x"139CCF7",
    x"139CA84",
    x"139C811",
    x"139C5A0",
    x"139C32E",
    x"139C0BE",
    x"139BE4E",
    x"139BBDF",
    x"139B970",
    x"139B702",
    x"139B495",
    x"139B228",
    x"139AFBC",
    x"139AD50",
    x"139AAE5",
    x"139A87B",
    x"139A611",
    x"139A3A7",
    x"139A13F",
    x"1399ED7",
    x"1399C6F",
    x"1399A09",
    x"13997A2",
    x"139953D",
    x"13992D8",
    x"1399073",
    x"1398E10",
    x"1398BAC",
    x"139894A",
    x"13986E8",
    x"1398486",
    x"1398225",
    x"1397FC5",
    x"1397D66",
    x"1397B07",
    x"13978A8",
    x"139764A",
    x"13973ED",
    x"1397190",
    x"1396F34",
    x"1396CD9",
    x"1396A7E",
    x"1396823",
    x"13965CA",
    x"1396370",
    x"1396118",
    x"1395EC0",
    x"1395C69",
    x"1395A12",
    x"13957BB",
    x"1395566",
    x"1395311",
    x"13950BC",
    x"1394E68",
    x"1394C15",
    x"13949C2",
    x"1394770",
    x"139451F",
    x"13942CE",
    x"139407D",
    x"1393E2D",
    x"1393BDE",
    x"139398F",
    x"1393741",
    x"13934F4",
    x"13932A7",
    x"139305B",
    x"1392E0F",
    x"1392BC4",
    x"1392979",
    x"139272F",
    x"13924E5",
    x"139229C",
    x"1392054",
    x"1391E0C",
    x"1391BC5",
    x"139197E",
    x"1391738",
    x"13914F3",
    x"13912AE",
    x"1391069",
    x"1390E25",
    x"1390BE2",
    x"13909A0",
    x"139075D",
    x"139051C",
    x"13902DB",
    x"139009A",
    x"138FE5B",
    x"138FC1B",
    x"138F9DD",
    x"138F79E",
    x"138F561",
    x"138F324",
    x"138F0E7",
    x"138EEAB",
    x"138EC70",
    x"138EA35",
    x"138E7FB",
    x"138E5C1",
    x"138E388",
    x"138E14F",
    x"138DF17",
    x"138DCE0",
    x"138DAA9",
    x"138D872",
    x"138D63C",
    x"138D407",
    x"138D1D2",
    x"138CF9E",
    x"138CD6B",
    x"138CB38",
    x"138C905",
    x"138C6D3",
    x"138C4A2",
    x"138C271",
    x"138C040",
    x"138BE11",
    x"138BBE1",
    x"138B9B3",
    x"138B785",
    x"138B557",
    x"138B32A",
    x"138B0FD",
    x"138AED1",
    x"138ACA6",
    x"138AA7B",
    x"138A851",
    x"138A627",
    x"138A3FE",
    x"138A1D5",
    x"1389FAD",
    x"1389D85",
    x"1389B5E",
    x"1389937",
    x"1389711",
    x"13894EC",
    x"13892C7",
    x"13890A2",
    x"1388E7F",
    x"1388C5B",
    x"1388A38",
    x"1388816",
    x"13885F4",
    x"13883D3",
    x"13881B2",
    x"1387F92",
    x"1387D73",
    x"1387B54",
    x"1387935",
    x"1387717",
    x"13874F9",
    x"13872DC",
    x"13870C0",
    x"1386EA4",
    x"1386C89",
    x"1386A6E",
    x"1386853",
    x"138663A",
    x"1386420",
    x"1386208",
    x"1385FEF",
    x"1385DD8",
    x"1385BC0",
    x"13859AA",
    x"1385794",
    x"138557E",
    x"1385369",
    x"1385154",
    x"1384F40",
    x"1384D2D",
    x"1384B1A",
    x"1384907",
    x"13846F5",
    x"13844E4",
    x"13842D3",
    x"13840C2",
    x"1383EB2",
    x"1383CA3",
    x"1383A94",
    x"1383886",
    x"1383678",
    x"138346A",
    x"138325D",
    x"1383051",
    x"1382E45",
    x"1382C3A",
    x"1382A2F",
    x"1382825",
    x"138261B",
    x"1382412",
    x"1382209",
    x"1382001",
    x"1381DF9",
    x"1381BF2",
    x"13819EB",
    x"13817E5",
    x"13815DF",
    x"13813DA",
    x"13811D5",
    x"1380FD1",
    x"1380DCD",
    x"1380BCA",
    x"13809C7",
    x"13807C5",
    x"13805C4",
    x"13803C2",
    x"13801C2",
    x"137FF83",
    x"137FB84",
    x"137F786",
    x"137F388",
    x"137EF8C",
    x"137EB90",
    x"137E796",
    x"137E39D",
    x"137DFA4",
    x"137DBAD",
    x"137D7B6",
    x"137D3C1",
    x"137CFCD",
    x"137CBD9",
    x"137C7E7",
    x"137C3F5",
    x"137C005",
    x"137BC15",
    x"137B827",
    x"137B439",
    x"137B04C",
    x"137AC61",
    x"137A876",
    x"137A48D",
    x"137A0A4",
    x"1379CBC",
    x"13798D6",
    x"13794F0",
    x"137910B",
    x"1378D27",
    x"1378945",
    x"1378563",
    x"1378182",
    x"1377DA2",
    x"13779C3",
    x"13775E5",
    x"1377208",
    x"1376E2C",
    x"1376A51",
    x"1376677",
    x"137629E",
    x"1375EC6",
    x"1375AEE",
    x"1375718",
    x"1375343",
    x"1374F6F",
    x"1374B9B",
    x"13747C9",
    x"13743F7",
    x"1374027",
    x"1373C57",
    x"1373889",
    x"13734BB",
    x"13730EE",
    x"1372D22",
    x"1372958",
    x"137258E",
    x"13721C5",
    x"1371DFD",
    x"1371A36",
    x"1371670",
    x"13712AB",
    x"1370EE6",
    x"1370B23",
    x"1370761",
    x"13703A0",
    x"136FFDF",
    x"136FC20",
    x"136F861",
    x"136F4A3",
    x"136F0E7",
    x"136ED2B",
    x"136E970",
    x"136E5B6",
    x"136E1FD",
    x"136DE45",
    x"136DA8E",
    x"136D6D8",
    x"136D323",
    x"136CF6E",
    x"136CBBB",
    x"136C808",
    x"136C457",
    x"136C0A6",
    x"136BCF7",
    x"136B948",
    x"136B59A",
    x"136B1ED",
    x"136AE41",
    x"136AA96",
    x"136A6EC",
    x"136A342",
    x"1369F9A",
    x"1369BF3",
    x"136984C",
    x"13694A6",
    x"1369102",
    x"1368D5E",
    x"13689BB",
    x"1368619",
    x"1368278",
    x"1367ED8",
    x"1367B39",
    x"136779A",
    x"13673FD",
    x"1367060",
    x"1366CC5",
    x"136692A",
    x"1366590",
    x"13661F7",
    x"1365E5F",
    x"1365AC8",
    x"1365732",
    x"136539C",
    x"1365008",
    x"1364C74",
    x"13648E2",
    x"1364550",
    x"13641BF",
    x"1363E2F",
    x"1363AA0",
    x"1363712",
    x"1363384",
    x"1362FF8",
    x"1362C6C",
    x"13628E2",
    x"1362558",
    x"13621CF",
    x"1361E47",
    x"1361AC0",
    x"136173A",
    x"13613B4",
    x"1361030",
    x"1360CAC",
    x"1360929",
    x"13605A8",
    x"1360227",
    x"135FEA7",
    x"135FB27",
    x"135F7A9",
    x"135F42B",
    x"135F0AF",
    x"135ED33",
    x"135E9B8",
    x"135E63E",
    x"135E2C5",
    x"135DF4D",
    x"135DBD5",
    x"135D85F",
    x"135D4E9",
    x"135D175",
    x"135CE01",
    x"135CA8E",
    x"135C71B",
    x"135C3AA",
    x"135C039",
    x"135BCCA",
    x"135B95B",
    x"135B5ED",
    x"135B280",
    x"135AF14",
    x"135ABA9",
    x"135A83E",
    x"135A4D4",
    x"135A16C",
    x"1359E04",
    x"1359A9D",
    x"1359736",
    x"13593D1",
    x"135906D",
    x"1358D09",
    x"13589A6",
    x"1358644",
    x"13582E3",
    x"1357F83",
    x"1357C23",
    x"13578C4",
    x"1357567",
    x"135720A",
    x"1356EAE",
    x"1356B52",
    x"13567F8",
    x"135649E",
    x"1356146",
    x"1355DEE",
    x"1355A97",
    x"1355741",
    x"13553EB",
    x"1355097",
    x"1354D43",
    x"13549F0",
    x"135469E",
    x"135434D",
    x"1353FFC",
    x"1353CAD",
    x"135395E",
    x"1353610",
    x"13532C3",
    x"1352F77",
    x"1352C2B",
    x"13528E0",
    x"1352597",
    x"135224E",
    x"1351F06",
    x"1351BBE",
    x"1351878",
    x"1351532",
    x"13511ED",
    x"1350EA9",
    x"1350B66",
    x"1350823",
    x"13504E2",
    x"13501A1",
    x"134FE61",
    x"134FB22",
    x"134F7E3",
    x"134F4A6",
    x"134F169",
    x"134EE2D",
    x"134EAF2",
    x"134E7B8",
    x"134E47E",
    x"134E145",
    x"134DE0D",
    x"134DAD6",
    x"134D7A0",
    x"134D46A",
    x"134D136",
    x"134CE02",
    x"134CACF",
    x"134C79C",
    x"134C46B",
    x"134C13A",
    x"134BE0A",
    x"134BADB",
    x"134B7AD",
    x"134B47F",
    x"134B153",
    x"134AE27",
    x"134AAFC",
    x"134A7D1",
    x"134A4A8",
    x"134A17F",
    x"1349E57",
    x"1349B30",
    x"1349809",
    x"13494E4",
    x"13491BF",
    x"1348E9B",
    x"1348B78",
    x"1348855",
    x"1348533",
    x"1348212",
    x"1347EF2",
    x"1347BD3",
    x"13478B4",
    x"1347597",
    x"134727A",
    x"1346F5D",
    x"1346C42",
    x"1346927",
    x"134660D",
    x"13462F4",
    x"1345FDC",
    x"1345CC4",
    x"13459AE",
    x"1345697",
    x"1345382",
    x"134506E",
    x"1344D5A",
    x"1344A47",
    x"1344735",
    x"1344423",
    x"1344113",
    x"1343E03",
    x"1343AF4",
    x"13437E5",
    x"13434D8",
    x"13431CB",
    x"1342EBF",
    x"1342BB4",
    x"13428A9",
    x"134259F",
    x"1342296",
    x"1341F8E",
    x"1341C86",
    x"1341980",
    x"134167A",
    x"1341374",
    x"1341070",
    x"1340D6C",
    x"1340A69",
    x"1340767",
    x"1340466",
    x"1340165",
    x"133FE65",
    x"133FB66",
    x"133F867",
    x"133F569",
    x"133F26C",
    x"133EF70",
    x"133EC75",
    x"133E97A",
    x"133E680",
    x"133E387",
    x"133E08E",
    x"133DD96",
    x"133DA9F",
    x"133D7A9",
    x"133D4B4",
    x"133D1BF",
    x"133CECB",
    x"133CBD7",
    x"133C8E5",
    x"133C5F3",
    x"133C302",
    x"133C011",
    x"133BD22",
    x"133BA33",
    x"133B745",
    x"133B457",
    x"133B16B",
    x"133AE7F",
    x"133AB93",
    x"133A8A9",
    x"133A5BF",
    x"133A2D6",
    x"1339FEE",
    x"1339D06",
    x"1339A1F",
    x"1339739",
    x"1339453",
    x"133916F",
    x"1338E8B",
    x"1338BA7",
    x"13388C5",
    x"13385E3",
    x"1338302",
    x"1338022",
    x"1337D42",
    x"1337A63",
    x"1337785",
    x"13374A7",
    x"13371CA",
    x"1336EEE",
    x"1336C13",
    x"1336938",
    x"133665E",
    x"1336385",
    x"13360AD",
    x"1335DD5",
    x"1335AFE",
    x"1335827",
    x"1335552",
    x"133527D",
    x"1334FA8",
    x"1334CD5",
    x"1334A02",
    x"1334730",
    x"133445E",
    x"133418E",
    x"1333EBD",
    x"1333BEE",
    x"1333920",
    x"1333652",
    x"1333384",
    x"13330B8",
    x"1332DEC",
    x"1332B21",
    x"1332856",
    x"133258D",
    x"13322C4",
    x"1331FFB",
    x"1331D34",
    x"1331A6D",
    x"13317A6",
    x"13314E1",
    x"133121C",
    x"1330F58",
    x"1330C94",
    x"13309D2",
    x"133070F",
    x"133044E",
    x"133018D",
    x"132FECD",
    x"132FC0E",
    x"132F94F",
    x"132F691",
    x"132F3D4",
    x"132F117",
    x"132EE5B",
    x"132EBA0",
    x"132E8E6",
    x"132E62C",
    x"132E372",
    x"132E0BA",
    x"132DE02",
    x"132DB4B",
    x"132D894",
    x"132D5DF",
    x"132D32A",
    x"132D075",
    x"132CDC1",
    x"132CB0E",
    x"132C85C",
    x"132C5AA",
    x"132C2F9",
    x"132C049",
    x"132BD99",
    x"132BAEA",
    x"132B83B",
    x"132B58E",
    x"132B2E1",
    x"132B034",
    x"132AD88",
    x"132AADD",
    x"132A833",
    x"132A589",
    x"132A2E0",
    x"132A038",
    x"1329D90",
    x"1329AE9",
    x"1329843",
    x"132959D",
    x"13292F8",
    x"1329053",
    x"1328DB0",
    x"1328B0D",
    x"132886A",
    x"13285C8",
    x"1328327",
    x"1328087",
    x"1327DE7",
    x"1327B48",
    x"13278A9",
    x"132760C",
    x"132736E",
    x"13270D2",
    x"1326E36",
    x"1326B9B",
    x"1326900",
    x"1326666",
    x"13263CD",
    x"1326134",
    x"1325E9C",
    x"1325C05",
    x"132596E",
    x"13256D8",
    x"1325443",
    x"13251AE",
    x"1324F1A",
    x"1324C87",
    x"13249F4",
    x"1324762",
    x"13244D0",
    x"132423F",
    x"1323FAF",
    x"1323D1F",
    x"1323A90",
    x"1323802",
    x"1323574",
    x"13232E7",
    x"132305B",
    x"1322DCF",
    x"1322B44",
    x"13228BA",
    x"1322630",
    x"13223A6",
    x"132211E",
    x"1321E96",
    x"1321C0F",
    x"1321988",
    x"1321702",
    x"132147C",
    x"13211F8",
    x"1320F73",
    x"1320CF0",
    x"1320A6D",
    x"13207EB",
    x"1320569",
    x"13202E8",
    x"1320068",
    x"131FDE8",
    x"131FB69",
    x"131F8EA",
    x"131F66C",
    x"131F3EF",
    x"131F172",
    x"131EEF6",
    x"131EC7B",
    x"131EA00",
    x"131E786",
    x"131E50C",
    x"131E293",
    x"131E01B",
    x"131DDA3",
    x"131DB2C",
    x"131D8B5",
    x"131D640",
    x"131D3CA",
    x"131D156",
    x"131CEE2",
    x"131CC6E",
    x"131C9FB",
    x"131C789",
    x"131C518",
    x"131C2A7",
    x"131C036",
    x"131BDC7",
    x"131BB57",
    x"131B8E9",
    x"131B67B",
    x"131B40E",
    x"131B1A1",
    x"131AF35",
    x"131ACC9",
    x"131AA5F",
    x"131A7F4",
    x"131A58B",
    x"131A321",
    x"131A0B9",
    x"1319E51",
    x"1319BEA",
    x"1319983",
    x"131971D",
    x"13194B8",
    x"1319253",
    x"1318FEE",
    x"1318D8B",
    x"1318B28",
    x"13188C5",
    x"1318663",
    x"1318402",
    x"13181A1",
    x"1317F41",
    x"1317CE2",
    x"1317A83",
    x"1317824",
    x"13175C7",
    x"1317369",
    x"131710D",
    x"1316EB1",
    x"1316C56",
    x"13169FB",
    x"13167A1",
    x"1316547",
    x"13162EE",
    x"1316095",
    x"1315E3E",
    x"1315BE6",
    x"1315990",
    x"131573A",
    x"13154E4",
    x"131528F",
    x"131503B",
    x"1314DE7",
    x"1314B94",
    x"1314941",
    x"13146EF",
    x"131449E",
    x"131424D",
    x"1313FFD",
    x"1313DAD",
    x"1313B5E",
    x"131390F",
    x"13136C1",
    x"1313474",
    x"1313227",
    x"1312FDB",
    x"1312D8F",
    x"1312B44",
    x"13128F9",
    x"13126AF",
    x"1312466",
    x"131221D",
    x"1311FD5",
    x"1311D8D",
    x"1311B46",
    x"1311900",
    x"13116BA",
    x"1311474",
    x"1311230",
    x"1310FEB",
    x"1310DA8",
    x"1310B64",
    x"1310922",
    x"13106E0",
    x"131049E",
    x"131025E",
    x"131001D",
    x"130FDDE",
    x"130FB9E",
    x"130F960",
    x"130F722",
    x"130F4E4",
    x"130F2A7",
    x"130F06B",
    x"130EE2F",
    x"130EBF4",
    x"130E9B9",
    x"130E77F",
    x"130E545",
    x"130E30C",
    x"130E0D4",
    x"130DE9C",
    x"130DC64",
    x"130DA2E",
    x"130D7F7",
    x"130D5C2",
    x"130D38C",
    x"130D158",
    x"130CF24",
    x"130CCF0",
    x"130CABD",
    x"130C88B",
    x"130C659",
    x"130C428",
    x"130C1F7",
    x"130BFC7",
    x"130BD97",
    x"130BB68",
    x"130B939",
    x"130B70B",
    x"130B4DE",
    x"130B2B1",
    x"130B085",
    x"130AE59",
    x"130AC2D",
    x"130AA03",
    x"130A7D8",
    x"130A5AF",
    x"130A385",
    x"130A15D",
    x"1309F35",
    x"1309D0D",
    x"1309AE6",
    x"13098C0",
    x"130969A",
    x"1309475",
    x"1309250",
    x"130902B",
    x"1308E08",
    x"1308BE4",
    x"13089C2",
    x"130879F",
    x"130857E",
    x"130835D",
    x"130813C",
    x"1307F1C",
    x"1307CFD",
    x"1307ADE",
    x"13078BF",
    x"13076A1",
    x"1307484",
    x"1307267",
    x"130704B",
    x"1306E2F",
    x"1306C14",
    x"13069F9",
    x"13067DF",
    x"13065C5",
    x"13063AC",
    x"1306193",
    x"1305F7B",
    x"1305D63",
    x"1305B4C",
    x"1305936",
    x"1305720",
    x"130550A",
    x"13052F5",
    x"13050E1",
    x"1304ECD",
    x"1304CB9",
    x"1304AA6",
    x"1304894",
    x"1304682",
    x"1304471",
    x"1304260",
    x"130404F",
    x"1303E40",
    x"1303C30",
    x"1303A21",
    x"1303813",
    x"1303605",
    x"13033F8",
    x"13031EB",
    x"1302FDF",
    x"1302DD4",
    x"1302BC8",
    x"13029BE",
    x"13027B3",
    x"13025AA",
    x"13023A1",
    x"1302198",
    x"1301F90",
    x"1301D88",
    x"1301B81",
    x"130197A",
    x"1301774",
    x"130156F",
    x"130136A",
    x"1301165",
    x"1300F61",
    x"1300D5D",
    x"1300B5A",
    x"1300958",
    x"1300756",
    x"1300554",
    x"1300353",
    x"1300152",
    x"12FFEA5",
    x"12FFAA6",
    x"12FF6A8",
    x"12FF2AA",
    x"12FEEAE",
    x"12FEAB3",
    x"12FE6B9",
    x"12FE2C0",
    x"12FDEC8",
    x"12FDAD0",
    x"12FD6DA",
    x"12FD2E5",
    x"12FCEF1",
    x"12FCAFD",
    x"12FC70B",
    x"12FC31A",
    x"12FBF2A",
    x"12FBB3A",
    x"12FB74C",
    x"12FB35F",
    x"12FAF72",
    x"12FAB87",
    x"12FA79D",
    x"12FA3B3",
    x"12F9FCB",
    x"12F9BE3",
    x"12F97FD",
    x"12F9417",
    x"12F9033",
    x"12F8C4F",
    x"12F886D",
    x"12F848B",
    x"12F80AA",
    x"12F7CCB",
    x"12F78EC",
    x"12F750E",
    x"12F7131",
    x"12F6D56",
    x"12F697B",
    x"12F65A1",
    x"12F61C8",
    x"12F5DF0",
    x"12F5A19",
    x"12F5643",
    x"12F526E",
    x"12F4E9A",
    x"12F4AC6",
    x"12F46F4",
    x"12F4323",
    x"12F3F53",
    x"12F3B83",
    x"12F37B5",
    x"12F33E7",
    x"12F301B",
    x"12F2C4F",
    x"12F2885",
    x"12F24BB",
    x"12F20F2",
    x"12F1D2B",
    x"12F1964",
    x"12F159E",
    x"12F11D9",
    x"12F0E15",
    x"12F0A52",
    x"12F0690",
    x"12F02CF",
    x"12EFF0E",
    x"12EFB4F",
    x"12EF791",
    x"12EF3D3",
    x"12EF017",
    x"12EEC5B",
    x"12EE8A1",
    x"12EE4E7",
    x"12EE12E",
    x"12EDD76",
    x"12ED9C0",
    x"12ED60A",
    x"12ED255",
    x"12ECEA0",
    x"12ECAED",
    x"12EC73B",
    x"12EC38A",
    x"12EBFD9",
    x"12EBC2A",
    x"12EB87B",
    x"12EB4CD",
    x"12EB121",
    x"12EAD75",
    x"12EA9CA",
    x"12EA620",
    x"12EA277",
    x"12E9ECF",
    x"12E9B28",
    x"12E9781",
    x"12E93DC",
    x"12E9037",
    x"12E8C94",
    x"12E88F1",
    x"12E854F",
    x"12E81AE",
    x"12E7E0E",
    x"12E7A6F",
    x"12E76D1",
    x"12E7334",
    x"12E6F98",
    x"12E6BFC",
    x"12E6862",
    x"12E64C8",
    x"12E612F",
    x"12E5D97",
    x"12E5A00",
    x"12E566A",
    x"12E52D5",
    x"12E4F41",
    x"12E4BAD",
    x"12E481B",
    x"12E4489",
    x"12E40F9",
    x"12E3D69",
    x"12E39DA",
    x"12E364C",
    x"12E32BF",
    x"12E2F33",
    x"12E2BA7",
    x"12E281D",
    x"12E2493",
    x"12E210B",
    x"12E1D83",
    x"12E19FC",
    x"12E1676",
    x"12E12F1",
    x"12E0F6C",
    x"12E0BE9",
    x"12E0866",
    x"12E04E5",
    x"12E0164",
    x"12DFDE4",
    x"12DFA65",
    x"12DF6E7",
    x"12DF369",
    x"12DEFED",
    x"12DEC71",
    x"12DE8F7",
    x"12DE57D",
    x"12DE204",
    x"12DDE8C",
    x"12DDB15",
    x"12DD79E",
    x"12DD429",
    x"12DD0B4",
    x"12DCD41",
    x"12DC9CE",
    x"12DC65C",
    x"12DC2EB",
    x"12DBF7A",
    x"12DBC0B",
    x"12DB89C",
    x"12DB52F",
    x"12DB1C2",
    x"12DAE56",
    x"12DAAEA",
    x"12DA780",
    x"12DA417",
    x"12DA0AE",
    x"12D9D46",
    x"12D99DF",
    x"12D9679",
    x"12D9314",
    x"12D8FB0",
    x"12D8C4C",
    x"12D88EA",
    x"12D8588",
    x"12D8227",
    x"12D7EC7",
    x"12D7B68",
    x"12D7809",
    x"12D74AC",
    x"12D714F",
    x"12D6DF3",
    x"12D6A98",
    x"12D673E",
    x"12D63E4",
    x"12D608C",
    x"12D5D34",
    x"12D59DD",
    x"12D5687",
    x"12D5332",
    x"12D4FDD",
    x"12D4C8A",
    x"12D4937",
    x"12D45E5",
    x"12D4294",
    x"12D3F44",
    x"12D3BF5",
    x"12D38A6",
    x"12D3558",
    x"12D320B",
    x"12D2EBF",
    x"12D2B74",
    x"12D2829",
    x"12D24E0",
    x"12D2197",
    x"12D1E4F",
    x"12D1B08",
    x"12D17C2",
    x"12D147C",
    x"12D1137",
    x"12D0DF3",
    x"12D0AB0",
    x"12D076E",
    x"12D042D",
    x"12D00EC",
    x"12CFDAC",
    x"12CFA6D",
    x"12CF72F",
    x"12CF3F2",
    x"12CF0B5",
    x"12CED79",
    x"12CEA3E",
    x"12CE704",
    x"12CE3CB",
    x"12CE092",
    x"12CDD5A",
    x"12CDA24",
    x"12CD6ED",
    x"12CD3B8",
    x"12CD084",
    x"12CCD50",
    x"12CCA1D",
    x"12CC6EB",
    x"12CC3B9",
    x"12CC089",
    x"12CBD59",
    x"12CBA2A",
    x"12CB6FC",
    x"12CB3CF",
    x"12CB0A2",
    x"12CAD76",
    x"12CAA4B",
    x"12CA721",
    x"12CA3F8",
    x"12CA0CF",
    x"12C9DA7",
    x"12C9A80",
    x"12C975A",
    x"12C9435",
    x"12C9110",
    x"12C8DEC",
    x"12C8AC9",
    x"12C87A7",
    x"12C8485",
    x"12C8165",
    x"12C7E45",
    x"12C7B25",
    x"12C7807",
    x"12C74E9",
    x"12C71CD",
    x"12C6EB0",
    x"12C6B95",
    x"12C687B",
    x"12C6561",
    x"12C6248",
    x"12C5F30",
    x"12C5C18",
    x"12C5902",
    x"12C55EC",
    x"12C52D7",
    x"12C4FC2",
    x"12C4CAF",
    x"12C499C",
    x"12C468A",
    x"12C4379",
    x"12C4068",
    x"12C3D59",
    x"12C3A4A",
    x"12C373C",
    x"12C342E",
    x"12C3121",
    x"12C2E16",
    x"12C2B0A",
    x"12C2800",
    x"12C24F6",
    x"12C21EE",
    x"12C1EE5",
    x"12C1BDE",
    x"12C18D7",
    x"12C15D2",
    x"12C12CD",
    x"12C0FC8",
    x"12C0CC5",
    x"12C09C2",
    x"12C06C0",
    x"12C03BE",
    x"12C00BE",
    x"12BFDBE",
    x"12BFABF",
    x"12BF7C1",
    x"12BF4C3",
    x"12BF1C6",
    x"12BEECA",
    x"12BEBCF",
    x"12BE8D4",
    x"12BE5DB",
    x"12BE2E1",
    x"12BDFE9",
    x"12BDCF2",
    x"12BD9FB",
    x"12BD705",
    x"12BD40F",
    x"12BD11A",
    x"12BCE27",
    x"12BCB33",
    x"12BC841",
    x"12BC54F",
    x"12BC25E",
    x"12BBF6E",
    x"12BBC7F",
    x"12BB990",
    x"12BB6A2",
    x"12BB3B5",
    x"12BB0C8",
    x"12BADDC",
    x"12BAAF1",
    x"12BA807",
    x"12BA51D",
    x"12BA234",
    x"12B9F4C",
    x"12B9C64",
    x"12B997E",
    x"12B9698",
    x"12B93B2",
    x"12B90CE",
    x"12B8DEA",
    x"12B8B07",
    x"12B8825",
    x"12B8543",
    x"12B8262",
    x"12B7F82",
    x"12B7CA2",
    x"12B79C3",
    x"12B76E5",
    x"12B7408",
    x"12B712B",
    x"12B6E4F",
    x"12B6B74",
    x"12B689A",
    x"12B65C0",
    x"12B62E7",
    x"12B600E",
    x"12B5D37",
    x"12B5A60",
    x"12B5789",
    x"12B54B4",
    x"12B51DF",
    x"12B4F0B",
    x"12B4C38",
    x"12B4965",
    x"12B4693",
    x"12B43C2",
    x"12B40F1",
    x"12B3E21",
    x"12B3B52",
    x"12B3883",
    x"12B35B6",
    x"12B32E9",
    x"12B301C",
    x"12B2D51",
    x"12B2A86",
    x"12B27BB",
    x"12B24F2",
    x"12B2229",
    x"12B1F61",
    x"12B1C99",
    x"12B19D2",
    x"12B170C",
    x"12B1447",
    x"12B1182",
    x"12B0EBE",
    x"12B0BFB",
    x"12B0938",
    x"12B0676",
    x"12B03B5",
    x"12B00F4",
    x"12AFE34",
    x"12AFB75",
    x"12AF8B7",
    x"12AF5F9",
    x"12AF33C",
    x"12AF07F",
    x"12AEDC3",
    x"12AEB08",
    x"12AE84E",
    x"12AE594",
    x"12AE2DB",
    x"12AE023",
    x"12ADD6B",
    x"12ADAB4",
    x"12AD7FE",
    x"12AD548",
    x"12AD293",
    x"12ACFDF",
    x"12ACD2B",
    x"12ACA78",
    x"12AC7C6",
    x"12AC514",
    x"12AC263",
    x"12ABFB3",
    x"12ABD03",
    x"12ABA55",
    x"12AB7A6",
    x"12AB4F9",
    x"12AB24C",
    x"12AAFA0",
    x"12AACF4",
    x"12AAA49",
    x"12AA79F",
    x"12AA4F5",
    x"12AA24C",
    x"12A9FA4",
    x"12A9CFD",
    x"12A9A56",
    x"12A97AF",
    x"12A950A",
    x"12A9265",
    x"12A8FC1",
    x"12A8D1D",
    x"12A8A7A",
    x"12A87D8",
    x"12A8536",
    x"12A8295",
    x"12A7FF5",
    x"12A7D55",
    x"12A7AB6",
    x"12A7818",
    x"12A757A",
    x"12A72DD",
    x"12A7041",
    x"12A6DA5",
    x"12A6B0A",
    x"12A686F",
    x"12A65D6",
    x"12A633C",
    x"12A60A4",
    x"12A5E0C",
    x"12A5B75",
    x"12A58DE",
    x"12A5649",
    x"12A53B3",
    x"12A511F",
    x"12A4E8B",
    x"12A4BF7",
    x"12A4965",
    x"12A46D3",
    x"12A4441",
    x"12A41B1",
    x"12A3F20",
    x"12A3C91",
    x"12A3A02",
    x"12A3774",
    x"12A34E6",
    x"12A325A",
    x"12A2FCD",
    x"12A2D42",
    x"12A2AB7",
    x"12A282C",
    x"12A25A3",
    x"12A2319",
    x"12A2091",
    x"12A1E09",
    x"12A1B82",
    x"12A18FB",
    x"12A1676",
    x"12A13F0",
    x"12A116C",
    x"12A0EE8",
    x"12A0C64",
    x"12A09E1",
    x"12A075F",
    x"12A04DE",
    x"12A025D",
    x"129FFDC",
    x"129FD5D",
    x"129FADE",
    x"129F85F",
    x"129F5E2",
    x"129F364",
    x"129F0E8",
    x"129EE6C",
    x"129EBF1",
    x"129E976",
    x"129E6FC",
    x"129E482",
    x"129E20A",
    x"129DF91",
    x"129DD1A",
    x"129DAA3",
    x"129D82D",
    x"129D5B7",
    x"129D342",
    x"129D0CD",
    x"129CE59",
    x"129CBE6",
    x"129C973",
    x"129C701",
    x"129C490",
    x"129C21F",
    x"129BFAF",
    x"129BD3F",
    x"129BAD0",
    x"129B862",
    x"129B5F4",
    x"129B387",
    x"129B11A",
    x"129AEAE",
    x"129AC43",
    x"129A9D8",
    x"129A76E",
    x"129A504",
    x"129A29B",
    x"129A033",
    x"1299DCB",
    x"1299B64",
    x"12998FE",
    x"1299698",
    x"1299432",
    x"12991CE",
    x"1298F69",
    x"1298D06",
    x"1298AA3",
    x"1298841",
    x"12985DF",
    x"129837E",
    x"129811D",
    x"1297EBD",
    x"1297C5E",
    x"12979FF",
    x"12977A1",
    x"1297543",
    x"12972E6",
    x"129708A",
    x"1296E2E",
    x"1296BD3",
    x"1296978",
    x"129671E",
    x"12964C4",
    x"129626B",
    x"1296013",
    x"1295DBB",
    x"1295B64",
    x"129590E",
    x"12956B8",
    x"1295462",
    x"129520E",
    x"1294FB9",
    x"1294D66",
    x"1294B13",
    x"12948C0",
    x"129466E",
    x"129441D",
    x"12941CC",
    x"1293F7C",
    x"1293D2C",
    x"1293ADD",
    x"129388F",
    x"1293641",
    x"12933F4",
    x"12931A7",
    x"1292F5B",
    x"1292D0F",
    x"1292AC4",
    x"129287A",
    x"1292630",
    x"12923E7",
    x"129219E",
    x"1291F56",
    x"1291D0F",
    x"1291AC8",
    x"1291881",
    x"129163B",
    x"12913F6",
    x"12911B1",
    x"1290F6D",
    x"1290D2A",
    x"1290AE7",
    x"12908A4",
    x"1290662",
    x"1290421",
    x"12901E0",
    x"128FFA0",
    x"128FD60",
    x"128FB21",
    x"128F8E3",
    x"128F6A5",
    x"128F468",
    x"128F22B",
    x"128EFEF",
    x"128EDB3",
    x"128EB78",
    x"128E93D",
    x"128E703",
    x"128E4CA",
    x"128E291",
    x"128E058",
    x"128DE20",
    x"128DBE9",
    x"128D9B3",
    x"128D77C",
    x"128D547",
    x"128D312",
    x"128D0DD",
    x"128CEA9",
    x"128CC76",
    x"128CA43",
    x"128C811",
    x"128C5DF",
    x"128C3AE",
    x"128C17D",
    x"128BF4D",
    x"128BD1E",
    x"128BAEF",
    x"128B8C0",
    x"128B692",
    x"128B465",
    x"128B238",
    x"128B00C",
    x"128ADE0",
    x"128ABB5",
    x"128A98A",
    x"128A760",
    x"128A536",
    x"128A30D",
    x"128A0E5",
    x"1289EBD",
    x"1289C95",
    x"1289A6F",
    x"1289848",
    x"1289622",
    x"12893FD",
    x"12891D8",
    x"1288FB4",
    x"1288D91",
    x"1288B6E",
    x"128894B",
    x"1288729",
    x"1288507",
    x"12882E6",
    x"12880C6",
    x"1287EA6",
    x"1287C87",
    x"1287A68",
    x"1287849",
    x"128762C",
    x"128740E",
    x"12871F2",
    x"1286FD5",
    x"1286DBA",
    x"1286B9E",
    x"1286984",
    x"128676A",
    x"1286550",
    x"1286337",
    x"128611E",
    x"1285F06",
    x"1285CEF",
    x"1285AD8",
    x"12858C2",
    x"12856AC",
    x"1285496",
    x"1285281",
    x"128506D",
    x"1284E59",
    x"1284C46",
    x"1284A33",
    x"1284821",
    x"128460F",
    x"12843FE",
    x"12841ED",
    x"1283FDD",
    x"1283DCD",
    x"1283BBE",
    x"12839AF",
    x"12837A1",
    x"1283593",
    x"1283386",
    x"128317A",
    x"1282F6D",
    x"1282D62",
    x"1282B57",
    x"128294C",
    x"1282742",
    x"1282539",
    x"128232F",
    x"1282127",
    x"1281F1F",
    x"1281D17",
    x"1281B10",
    x"128190A",
    x"1281704",
    x"12814FE",
    x"12812F9",
    x"12810F5",
    x"1280EF1",
    x"1280CED",
    x"1280AEA",
    x"12808E8",
    x"12806E6",
    x"12804E4",
    x"12802E3",
    x"12800E3",
    x"127FDC7",
    x"127F9C8",
    x"127F5CA",
    x"127F1CD",
    x"127EDD1",
    x"127E9D6",
    x"127E5DC",
    x"127E1E3",
    x"127DDEB",
    x"127D9F4",
    x"127D5FE",
    x"127D209",
    x"127CE15",
    x"127CA22",
    x"127C630",
    x"127C23F",
    x"127BE4F",
    x"127BA60",
    x"127B671",
    x"127B284",
    x"127AE98",
    x"127AAAD",
    x"127A6C3",
    x"127A2DA",
    x"1279EF1",
    x"1279B0A",
    x"1279724",
    x"127933F",
    x"1278F5A",
    x"1278B77",
    x"1278795",
    x"12783B3",
    x"1277FD3",
    x"1277BF3",
    x"1277815",
    x"1277437",
    x"127705B",
    x"1276C7F",
    x"12768A4",
    x"12764CB",
    x"12760F2",
    x"1275D1A",
    x"1275943",
    x"127556E",
    x"1275199",
    x"1274DC5",
    x"12749F2",
    x"1274620",
    x"127424F",
    x"1273E7F",
    x"1273AB0",
    x"12736E1",
    x"1273314",
    x"1272F48",
    x"1272B7C",
    x"12727B2",
    x"12723E9",
    x"1272020",
    x"1271C59",
    x"1271892",
    x"12714CC",
    x"1271108",
    x"1270D44",
    x"1270981",
    x"12705BF",
    x"12701FE",
    x"126FE3E",
    x"126FA7F",
    x"126F6C1",
    x"126F304",
    x"126EF47",
    x"126EB8C",
    x"126E7D1",
    x"126E418",
    x"126E05F",
    x"126DCA8",
    x"126D8F1",
    x"126D53B",
    x"126D186",
    x"126CDD3",
    x"126CA20",
    x"126C66D",
    x"126C2BC",
    x"126BF0C",
    x"126BB5D",
    x"126B7AE",
    x"126B401",
    x"126B054",
    x"126ACA9",
    x"126A8FE",
    x"126A554",
    x"126A1AB",
    x"1269E03",
    x"1269A5C",
    x"12696B6",
    x"1269311",
    x"1268F6D",
    x"1268BC9",
    x"1268827",
    x"1268485",
    x"12680E5",
    x"1267D45",
    x"12679A6",
    x"1267608",
    x"126726B",
    x"1266ECF",
    x"1266B34",
    x"1266799",
    x"1266400",
    x"1266067",
    x"1265CD0",
    x"1265939",
    x"12655A3",
    x"126520E",
    x"1264E7A",
    x"1264AE7",
    x"1264754",
    x"12643C3",
    x"1264033",
    x"1263CA3",
    x"1263914",
    x"1263586",
    x"12631F9",
    x"1262E6D",
    x"1262AE2",
    x"1262758",
    x"12623CF",
    x"1262046",
    x"1261CBE",
    x"1261938",
    x"12615B2",
    x"126122D",
    x"1260EA9",
    x"1260B26",
    x"12607A3",
    x"1260422",
    x"12600A1",
    x"125FD21",
    x"125F9A3",
    x"125F625",
    x"125F2A7",
    x"125EF2B",
    x"125EBB0",
    x"125E835",
    x"125E4BC",
    x"125E143",
    x"125DDCB",
    x"125DA54",
    x"125D6DE",
    x"125D369",
    x"125CFF4",
    x"125CC81",
    x"125C90E",
    x"125C59C",
    x"125C22B",
    x"125BEBB",
    x"125BB4C",
    x"125B7DD",
    x"125B470",
    x"125B103",
    x"125AD97",
    x"125AA2C",
    x"125A6C2",
    x"125A359",
    x"1259FF1",
    x"1259C89",
    x"1259922",
    x"12595BD",
    x"1259257",
    x"1258EF3",
    x"1258B90",
    x"125882E",
    x"12584CC",
    x"125816B",
    x"1257E0B",
    x"1257AAC",
    x"125774E",
    x"12573F0",
    x"1257094",
    x"1256D38",
    x"12569DD",
    x"1256683",
    x"125632A",
    x"1255FD2",
    x"1255C7A",
    x"1255923",
    x"12555CE",
    x"1255279",
    x"1254F24",
    x"1254BD1",
    x"125487E",
    x"125452D",
    x"12541DC",
    x"1253E8C",
    x"1253B3D",
    x"12537EE",
    x"12534A1",
    x"1253154",
    x"1252E08",
    x"1252ABD",
    x"1252773",
    x"1252429",
    x"12520E0",
    x"1251D99",
    x"1251A52",
    x"125170C",
    x"12513C6",
    x"1251082",
    x"1250D3E",
    x"12509FB",
    x"12506B9",
    x"1250378",
    x"1250037",
    x"124FCF8",
    x"124F9B9",
    x"124F67B",
    x"124F33D",
    x"124F001",
    x"124ECC5",
    x"124E98B",
    x"124E651",
    x"124E317",
    x"124DFDF",
    x"124DCA8",
    x"124D971",
    x"124D63B",
    x"124D306",
    x"124CFD1",
    x"124CC9E",
    x"124C96B",
    x"124C639",
    x"124C308",
    x"124BFD8",
    x"124BCA8",
    x"124B979",
    x"124B64B",
    x"124B31E",
    x"124AFF2",
    x"124ACC6",
    x"124A99B",
    x"124A671",
    x"124A348",
    x"124A020",
    x"1249CF8",
    x"12499D1",
    x"12496AB",
    x"1249386",
    x"1249061",
    x"1248D3E",
    x"1248A1B",
    x"12486F9",
    x"12483D7",
    x"12480B7",
    x"1247D97",
    x"1247A78",
    x"124775A",
    x"124743C",
    x"1247120",
    x"1246E04",
    x"1246AE9",
    x"12467CE",
    x"12464B5",
    x"124619C",
    x"1245E84",
    x"1245B6D",
    x"1245856",
    x"1245540",
    x"124522B",
    x"1244F17",
    x"1244C04",
    x"12448F1",
    x"12445DF",
    x"12442CE",
    x"1243FBE",
    x"1243CAE",
    x"12439A0",
    x"1243692",
    x"1243384",
    x"1243078",
    x"1242D6C",
    x"1242A61",
    x"1242757",
    x"124244E",
    x"1242145",
    x"1241E3D",
    x"1241B36",
    x"124182F",
    x"124152A",
    x"1241225",
    x"1240F21",
    x"1240C1D",
    x"124091A",
    x"1240619",
    x"1240317",
    x"1240017",
    x"123FD17",
    x"123FA18",
    x"123F71A",
    x"123F41D",
    x"123F120",
    x"123EE24",
    x"123EB29",
    x"123E82F",
    x"123E535",
    x"123E23C",
    x"123DF44",
    x"123DC4D",
    x"123D956",
    x"123D660",
    x"123D36B",
    x"123D076",
    x"123CD82",
    x"123CA8F",
    x"123C79D",
    x"123C4AC",
    x"123C1BB",
    x"123BECB",
    x"123BBDB",
    x"123B8ED",
    x"123B5FF",
    x"123B312",
    x"123B025",
    x"123AD3A",
    x"123AA4F",
    x"123A765",
    x"123A47B",
    x"123A192",
    x"1239EAA",
    x"1239BC3",
    x"12398DC",
    x"12395F7",
    x"1239311",
    x"123902D",
    x"1238D49",
    x"1238A66",
    x"1238784",
    x"12384A3",
    x"12381C2",
    x"1237EE2",
    x"1237C02",
    x"1237924",
    x"1237646",
    x"1237369",
    x"123708C",
    x"1236DB0",
    x"1236AD5",
    x"12367FB",
    x"1236521",
    x"1236248",
    x"1235F70",
    x"1235C99",
    x"12359C2",
    x"12356EC",
    x"1235416",
    x"1235142",
    x"1234E6E",
    x"1234B9A",
    x"12348C8",
    x"12345F6",
    x"1234325",
    x"1234055",
    x"1233D85",
    x"1233AB6",
    x"12337E7",
    x"123351A",
    x"123324D",
    x"1232F81",
    x"1232CB5",
    x"12329EA",
    x"1232720",
    x"1232457",
    x"123218E",
    x"1231EC6",
    x"1231BFF",
    x"1231938",
    x"1231672",
    x"12313AD",
    x"12310E8",
    x"1230E24",
    x"1230B61",
    x"123089F",
    x"12305DD",
    x"123031C",
    x"123005B",
    x"122FD9B",
    x"122FADC",
    x"122F81E",
    x"122F560",
    x"122F2A3",
    x"122EFE7",
    x"122ED2B",
    x"122EA70",
    x"122E7B6",
    x"122E4FD",
    x"122E244",
    x"122DF8B",
    x"122DCD4",
    x"122DA1D",
    x"122D767",
    x"122D4B1",
    x"122D1FD",
    x"122CF48",
    x"122CC95",
    x"122C9E2",
    x"122C730",
    x"122C47E",
    x"122C1CE",
    x"122BF1E",
    x"122BC6E",
    x"122B9BF",
    x"122B711",
    x"122B464",
    x"122B1B7",
    x"122AF0B",
    x"122AC60",
    x"122A9B5",
    x"122A70B",
    x"122A461",
    x"122A1B8",
    x"1229F10",
    x"1229C69",
    x"12299C2",
    x"122971C",
    x"1229477",
    x"12291D2",
    x"1228F2E",
    x"1228C8A",
    x"12289E7",
    x"1228745",
    x"12284A4",
    x"1228203",
    x"1227F63",
    x"1227CC3",
    x"1227A24",
    x"1227786",
    x"12274E9",
    x"122724C",
    x"1226FB0",
    x"1226D14",
    x"1226A79",
    x"12267DF",
    x"1226545",
    x"12262AC",
    x"1226014",
    x"1225D7C",
    x"1225AE5",
    x"122584F",
    x"12255B9",
    x"1225324",
    x"122508F",
    x"1224DFB",
    x"1224B68",
    x"12248D6",
    x"1224644",
    x"12243B3",
    x"1224122",
    x"1223E92",
    x"1223C03",
    x"1223974",
    x"12236E6",
    x"1223459",
    x"12231CC",
    x"1222F40",
    x"1222CB4",
    x"1222A29",
    x"122279F",
    x"1222515",
    x"122228D",
    x"1222004",
    x"1221D7D",
    x"1221AF5",
    x"122186F",
    x"12215E9",
    x"1221364",
    x"12210E0",
    x"1220E5C",
    x"1220BD8",
    x"1220956",
    x"12206D4",
    x"1220452",
    x"12201D2",
    x"121FF51",
    x"121FCD2",
    x"121FA53",
    x"121F7D5",
    x"121F557",
    x"121F2DA",
    x"121F05E",
    x"121EDE2",
    x"121EB67",
    x"121E8EC",
    x"121E672",
    x"121E3F9",
    x"121E180",
    x"121DF08",
    x"121DC91",
    x"121DA1A",
    x"121D7A4",
    x"121D52E",
    x"121D2B9",
    x"121D045",
    x"121CDD1",
    x"121CB5E",
    x"121C8EB",
    x"121C679",
    x"121C408",
    x"121C197",
    x"121BF27",
    x"121BCB8",
    x"121BA49",
    x"121B7DB",
    x"121B56D",
    x"121B300",
    x"121B093",
    x"121AE28",
    x"121ABBC",
    x"121A952",
    x"121A6E8",
    x"121A47E",
    x"121A215",
    x"1219FAD",
    x"1219D46",
    x"1219ADF",
    x"1219878",
    x"1219612",
    x"12193AD",
    x"1219149",
    x"1218EE5",
    x"1218C81",
    x"1218A1E",
    x"12187BC",
    x"121855A",
    x"12182F9",
    x"1218099",
    x"1217E39",
    x"1217BDA",
    x"121797B",
    x"121771D",
    x"12174C0",
    x"1217263",
    x"1217006",
    x"1216DAB",
    x"1216B50",
    x"12168F5",
    x"121669B",
    x"1216442",
    x"12161E9",
    x"1215F91",
    x"1215D39",
    x"1215AE2",
    x"121588C",
    x"1215636",
    x"12153E1",
    x"121518C",
    x"1214F38",
    x"1214CE4",
    x"1214A91",
    x"121483F",
    x"12145ED",
    x"121439C",
    x"121414B",
    x"1213EFB",
    x"1213CAC",
    x"1213A5D",
    x"121380F",
    x"12135C1",
    x"1213374",
    x"1213127",
    x"1212EDB",
    x"1212C90",
    x"1212A45",
    x"12127FB",
    x"12125B1",
    x"1212368",
    x"121211F",
    x"1211ED7",
    x"1211C90",
    x"1211A49",
    x"1211803",
    x"12115BD",
    x"1211378",
    x"1211133",
    x"1210EEF",
    x"1210CAC",
    x"1210A69",
    x"1210827",
    x"12105E5",
    x"12103A4",
    x"1210163",
    x"120FF23",
    x"120FCE3",
    x"120FAA5",
    x"120F866",
    x"120F628",
    x"120F3EB",
    x"120F1AE",
    x"120EF72",
    x"120ED37",
    x"120EAFC",
    x"120E8C1",
    x"120E687",
    x"120E44E",
    x"120E215",
    x"120DFDD",
    x"120DDA5",
    x"120DB6E",
    x"120D937",
    x"120D701",
    x"120D4CC",
    x"120D297",
    x"120D063",
    x"120CE2F",
    x"120CBFC",
    x"120C9C9",
    x"120C797",
    x"120C565",
    x"120C334",
    x"120C103",
    x"120BED3",
    x"120BCA4",
    x"120BA75",
    x"120B847",
    x"120B619",
    x"120B3EC",
    x"120B1BF",
    x"120AF93",
    x"120AD67",
    x"120AB3C",
    x"120A912",
    x"120A6E8",
    x"120A4BE",
    x"120A295",
    x"120A06D",
    x"1209E45",
    x"1209C1E",
    x"12099F7",
    x"12097D1",
    x"12095AB",
    x"1209386",
    x"1209161",
    x"1208F3D",
    x"1208D1A",
    x"1208AF7",
    x"12088D4",
    x"12086B2",
    x"1208491",
    x"1208270",
    x"1208050",
    x"1207E30",
    x"1207C11",
    x"12079F2",
    x"12077D4",
    x"12075B6",
    x"1207399",
    x"120717C",
    x"1206F60",
    x"1206D44",
    x"1206B29",
    x"120690F",
    x"12066F5",
    x"12064DB",
    x"12062C2",
    x"12060AA",
    x"1205E92",
    x"1205C7B",
    x"1205A64",
    x"120584D",
    x"1205638",
    x"1205422",
    x"120520E",
    x"1204FF9",
    x"1204DE6",
    x"1204BD2",
    x"12049C0",
    x"12047AE",
    x"120459C",
    x"120438B",
    x"120417A",
    x"1203F6A",
    x"1203D5A",
    x"1203B4B",
    x"120393D",
    x"120372F",
    x"1203521",
    x"1203314",
    x"1203108",
    x"1202EFC",
    x"1202CF0",
    x"1202AE5",
    x"12028DB",
    x"12026D1",
    x"12024C7",
    x"12022BE",
    x"12020B6",
    x"1201EAE",
    x"1201CA7",
    x"1201AA0",
    x"1201899",
    x"1201693",
    x"120148E",
    x"1201289",
    x"1201085",
    x"1200E81",
    x"1200C7D",
    x"1200A7B",
    x"1200878",
    x"1200676",
    x"1200475",
    x"1200274",
    x"1200074",
    x"11FFCE8",
    x"11FF8E9",
    x"11FF4EC",
    x"11FF0EF",
    x"11FECF3",
    x"11FE8F8",
    x"11FE4FF",
    x"11FE106",
    x"11FDD0E",
    x"11FD917",
    x"11FD522",
    x"11FD12D",
    x"11FCD39",
    x"11FC946",
    x"11FC554",
    x"11FC164",
    x"11FBD74",
    x"11FB985",
    x"11FB597",
    x"11FB1AA",
    x"11FADBE",
    x"11FA9D3",
    x"11FA5E9",
    x"11FA200",
    x"11F9E18",
    x"11F9A31",
    x"11F964B",
    x"11F9266",
    x"11F8E82",
    x"11F8A9F",
    x"11F86BD",
    x"11F82DB",
    x"11F7EFB",
    x"11F7B1C",
    x"11F773E",
    x"11F7360",
    x"11F6F84",
    x"11F6BA9",
    x"11F67CE",
    x"11F63F5",
    x"11F601C",
    x"11F5C45",
    x"11F586E",
    x"11F5498",
    x"11F50C4",
    x"11F4CF0",
    x"11F491D",
    x"11F454B",
    x"11F417B",
    x"11F3DAB",
    x"11F39DC",
    x"11F360E",
    x"11F3241",
    x"11F2E75",
    x"11F2AAA",
    x"11F26DF",
    x"11F2316",
    x"11F1F4E",
    x"11F1B86",
    x"11F17C0",
    x"11F13FB",
    x"11F1036",
    x"11F0C72",
    x"11F08B0",
    x"11F04EE",
    x"11F012D",
    x"11EFD6D",
    x"11EF9AF",
    x"11EF5F1",
    x"11EF234",
    x"11EEE78",
    x"11EEABC",
    x"11EE702",
    x"11EE349",
    x"11EDF91",
    x"11EDBD9",
    x"11ED823",
    x"11ED46D",
    x"11ED0B8",
    x"11ECD05",
    x"11EC952",
    x"11EC5A0",
    x"11EC1EF",
    x"11EBE3F",
    x"11EBA90",
    x"11EB6E2",
    x"11EB335",
    x"11EAF88",
    x"11EABDD",
    x"11EA832",
    x"11EA489",
    x"11EA0E0",
    x"11E9D38",
    x"11E9991",
    x"11E95EB",
    x"11E9246",
    x"11E8EA2",
    x"11E8AFF",
    x"11E875D",
    x"11E83BB",
    x"11E801B",
    x"11E7C7B",
    x"11E78DD",
    x"11E753F",
    x"11E71A2",
    x"11E6E06",
    x"11E6A6B",
    x"11E66D1",
    x"11E6338",
    x"11E5F9F",
    x"11E5C08",
    x"11E5871",
    x"11E54DC",
    x"11E5147",
    x"11E4DB3",
    x"11E4A20",
    x"11E468E",
    x"11E42FD",
    x"11E3F6C",
    x"11E3BDD",
    x"11E384E",
    x"11E34C1",
    x"11E3134",
    x"11E2DA8",
    x"11E2A1D",
    x"11E2693",
    x"11E230A",
    x"11E1F82",
    x"11E1BFA",
    x"11E1874",
    x"11E14EE",
    x"11E1169",
    x"11E0DE5",
    x"11E0A62",
    x"11E06E0",
    x"11E035F",
    x"11DFFDE",
    x"11DFC5F",
    x"11DF8E0",
    x"11DF562",
    x"11DF1E6",
    x"11DEE69",
    x"11DEAEE",
    x"11DE774",
    x"11DE3FB",
    x"11DE082",
    x"11DDD0A",
    x"11DD993",
    x"11DD61E",
    x"11DD2A8",
    x"11DCF34",
    x"11DCBC1",
    x"11DC84E",
    x"11DC4DD",
    x"11DC16C",
    x"11DBDFC",
    x"11DBA8D",
    x"11DB71F",
    x"11DB3B1",
    x"11DB045",
    x"11DACD9",
    x"11DA96E",
    x"11DA604",
    x"11DA29B",
    x"11D9F33",
    x"11D9BCC",
    x"11D9865",
    x"11D9500",
    x"11D919B",
    x"11D8E37",
    x"11D8AD4",
    x"11D8771",
    x"11D8410",
    x"11D80AF",
    x"11D7D50",
    x"11D79F1",
    x"11D7693",
    x"11D7335",
    x"11D6FD9",
    x"11D6C7D",
    x"11D6923",
    x"11D65C9",
    x"11D6270",
    x"11D5F18",
    x"11D5BC0",
    x"11D586A",
    x"11D5514",
    x"11D51BF",
    x"11D4E6B",
    x"11D4B18",
    x"11D47C6",
    x"11D4474",
    x"11D4123",
    x"11D3DD4",
    x"11D3A85",
    x"11D3736",
    x"11D33E9",
    x"11D309C",
    x"11D2D51",
    x"11D2A06",
    x"11D26BC",
    x"11D2372",
    x"11D202A",
    x"11D1CE2",
    x"11D199B",
    x"11D1655",
    x"11D1310",
    x"11D0FCC",
    x"11D0C88",
    x"11D0946",
    x"11D0604",
    x"11D02C3",
    x"11CFF82",
    x"11CFC43",
    x"11CF904",
    x"11CF5C6",
    x"11CF289",
    x"11CEF4D",
    x"11CEC12",
    x"11CE8D7",
    x"11CE59D",
    x"11CE264",
    x"11CDF2C",
    x"11CDBF5",
    x"11CD8BE",
    x"11CD588",
    x"11CD253",
    x"11CCF1F",
    x"11CCBEC",
    x"11CC8B9",
    x"11CC587",
    x"11CC256",
    x"11CBF26",
    x"11CBBF7",
    x"11CB8C8",
    x"11CB59A",
    x"11CB26D",
    x"11CAF41",
    x"11CAC16",
    x"11CA8EB",
    x"11CA5C1",
    x"11CA298",
    x"11C9F70",
    x"11C9C49",
    x"11C9922",
    x"11C95FC",
    x"11C92D7",
    x"11C8FB3",
    x"11C8C8F",
    x"11C896C",
    x"11C864A",
    x"11C8329",
    x"11C8009",
    x"11C7CE9",
    x"11C79CA",
    x"11C76AC",
    x"11C738F",
    x"11C7073",
    x"11C6D57",
    x"11C6A3C",
    x"11C6722",
    x"11C6408",
    x"11C60F0",
    x"11C5DD8",
    x"11C5AC1",
    x"11C57AA",
    x"11C5495",
    x"11C5180",
    x"11C4E6C",
    x"11C4B59",
    x"11C4846",
    x"11C4535",
    x"11C4224",
    x"11C3F14",
    x"11C3C04",
    x"11C38F6",
    x"11C35E8",
    x"11C32DB",
    x"11C2FCE",
    x"11C2CC3",
    x"11C29B8",
    x"11C26AE",
    x"11C23A5",
    x"11C209C",
    x"11C1D94",
    x"11C1A8D",
    x"11C1787",
    x"11C1482",
    x"11C117D",
    x"11C0E79",
    x"11C0B76",
    x"11C0873",
    x"11C0571",
    x"11C0270",
    x"11BFF70",
    x"11BFC71",
    x"11BF972",
    x"11BF674",
    x"11BF377",
    x"11BF07A",
    x"11BED7E",
    x"11BEA83",
    x"11BE789",
    x"11BE490",
    x"11BE197",
    x"11BDE9F",
    x"11BDBA8",
    x"11BD8B1",
    x"11BD5BB",
    x"11BD2C6",
    x"11BCFD2",
    x"11BCCDE",
    x"11BC9EB",
    x"11BC6F9",
    x"11BC408",
    x"11BC117",
    x"11BBE27",
    x"11BBB38",
    x"11BB84A",
    x"11BB55C",
    x"11BB26F",
    x"11BAF83",
    x"11BAC97",
    x"11BA9AD",
    x"11BA6C3",
    x"11BA3D9",
    x"11BA0F1",
    x"11B9E09",
    x"11B9B22",
    x"11B983B",
    x"11B9555",
    x"11B9271",
    x"11B8F8C",
    x"11B8CA9",
    x"11B89C6",
    x"11B86E4",
    x"11B8402",
    x"11B8122",
    x"11B7E42",
    x"11B7B63",
    x"11B7884",
    x"11B75A6",
    x"11B72C9",
    x"11B6FED",
    x"11B6D11",
    x"11B6A37",
    x"11B675C",
    x"11B6483",
    x"11B61AA",
    x"11B5ED2",
    x"11B5BFB",
    x"11B5924",
    x"11B564E",
    x"11B5379",
    x"11B50A4",
    x"11B4DD1",
    x"11B4AFD",
    x"11B482B",
    x"11B4559",
    x"11B4288",
    x"11B3FB8",
    x"11B3CE9",
    x"11B3A1A",
    x"11B374B",
    x"11B347E",
    x"11B31B1",
    x"11B2EE5",
    x"11B2C1A",
    x"11B294F",
    x"11B2685",
    x"11B23BC",
    x"11B20F3",
    x"11B1E2B",
    x"11B1B64",
    x"11B189E",
    x"11B15D8",
    x"11B1313",
    x"11B104E",
    x"11B0D8B",
    x"11B0AC8",
    x"11B0805",
    x"11B0544",
    x"11B0283",
    x"11AFFC2",
    x"11AFD03",
    x"11AFA44",
    x"11AF786",
    x"11AF4C8",
    x"11AF20B",
    x"11AEF4F",
    x"11AEC93",
    x"11AE9D9",
    x"11AE71F",
    x"11AE465",
    x"11AE1AC",
    x"11ADEF4",
    x"11ADC3D",
    x"11AD986",
    x"11AD6D0",
    x"11AD41B",
    x"11AD166",
    x"11ACEB2",
    x"11ACBFF",
    x"11AC94C",
    x"11AC69A",
    x"11AC3E9",
    x"11AC138",
    x"11ABE88",
    x"11ABBD9",
    x"11AB92A",
    x"11AB67C",
    x"11AB3CF",
    x"11AB122",
    x"11AAE76",
    x"11AABCB",
    x"11AA921",
    x"11AA677",
    x"11AA3CD",
    x"11AA125",
    x"11A9E7D",
    x"11A9BD5",
    x"11A992F",
    x"11A9689",
    x"11A93E4",
    x"11A913F",
    x"11A8E9B",
    x"11A8BF8",
    x"11A8955",
    x"11A86B3",
    x"11A8412",
    x"11A8171",
    x"11A7ED1",
    x"11A7C31",
    x"11A7993",
    x"11A76F5",
    x"11A7457",
    x"11A71BB",
    x"11A6F1E",
    x"11A6C83",
    x"11A69E8",
    x"11A674E",
    x"11A64B4",
    x"11A621C",
    x"11A5F83",
    x"11A5CEC",
    x"11A5A55",
    x"11A57BF",
    x"11A5529",
    x"11A5294",
    x"11A5000",
    x"11A4D6C",
    x"11A4AD9",
    x"11A4847",
    x"11A45B5",
    x"11A4324",
    x"11A4093",
    x"11A3E04",
    x"11A3B74",
    x"11A38E6",
    x"11A3658",
    x"11A33CB",
    x"11A313E",
    x"11A2EB2",
    x"11A2C27",
    x"11A299C",
    x"11A2712",
    x"11A2488",
    x"11A2200",
    x"11A1F77",
    x"11A1CF0",
    x"11A1A69",
    x"11A17E3",
    x"11A155D",
    x"11A12D8",
    x"11A1054",
    x"11A0DD0",
    x"11A0B4D",
    x"11A08CA",
    x"11A0648",
    x"11A03C7",
    x"11A0146",
    x"119FEC6",
    x"119FC47",
    x"119F9C8",
    x"119F74A",
    x"119F4CD",
    x"119F250",
    x"119EFD3",
    x"119ED58",
    x"119EADD",
    x"119E862",
    x"119E5E9",
    x"119E36F",
    x"119E0F7",
    x"119DE7F",
    x"119DC08",
    x"119D991",
    x"119D71B",
    x"119D4A5",
    x"119D230",
    x"119CFBC",
    x"119CD49",
    x"119CAD6",
    x"119C863",
    x"119C5F1",
    x"119C380",
    x"119C110",
    x"119BEA0",
    x"119BC30",
    x"119B9C2",
    x"119B753",
    x"119B4E6",
    x"119B279",
    x"119B00D",
    x"119ADA1",
    x"119AB36",
    x"119A8CB",
    x"119A661",
    x"119A3F8",
    x"119A190",
    x"1199F27",
    x"1199CC0",
    x"1199A59",
    x"11997F3",
    x"119958D",
    x"1199328",
    x"11990C3",
    x"1198E60",
    x"1198BFC",
    x"119899A",
    x"1198738",
    x"11984D6",
    x"1198275",
    x"1198015",
    x"1197DB5",
    x"1197B56",
    x"11978F7",
    x"1197699",
    x"119743C",
    x"11971DF",
    x"1196F83",
    x"1196D28",
    x"1196ACD",
    x"1196872",
    x"1196618",
    x"11963BF",
    x"1196166",
    x"1195F0E",
    x"1195CB7",
    x"1195A60",
    x"119580A",
    x"11955B4",
    x"119535F",
    x"119510A",
    x"1194EB6",
    x"1194C63",
    x"1194A10",
    x"11947BE",
    x"119456C",
    x"119431B",
    x"11940CB",
    x"1193E7B",
    x"1193C2C",
    x"11939DD",
    x"119378F",
    x"1193541",
    x"11932F4",
    x"11930A7",
    x"1192E5C",
    x"1192C10",
    x"11929C6",
    x"119277B",
    x"1192532",
    x"11922E9",
    x"11920A0",
    x"1191E59",
    x"1191C11",
    x"11919CA",
    x"1191784",
    x"119153F",
    x"11912FA",
    x"11910B5",
    x"1190E71",
    x"1190C2E",
    x"11909EB",
    x"11907A9",
    x"1190567",
    x"1190326",
    x"11900E6",
    x"118FEA6",
    x"118FC67",
    x"118FA28",
    x"118F7E9",
    x"118F5AC",
    x"118F36F",
    x"118F132",
    x"118EEF6",
    x"118ECBB",
    x"118EA80",
    x"118E845",
    x"118E60B",
    x"118E3D2",
    x"118E19A",
    x"118DF61",
    x"118DD2A",
    x"118DAF3",
    x"118D8BC",
    x"118D687",
    x"118D451",
    x"118D21C",
    x"118CFE8",
    x"118CDB4",
    x"118CB81",
    x"118C94F",
    x"118C71D",
    x"118C4EB",
    x"118C2BA",
    x"118C08A",
    x"118BE5A",
    x"118BC2B",
    x"118B9FC",
    x"118B7CE",
    x"118B5A0",
    x"118B373",
    x"118B146",
    x"118AF1A",
    x"118ACEF",
    x"118AAC4",
    x"118A899",
    x"118A66F",
    x"118A446",
    x"118A21D",
    x"1189FF5",
    x"1189DCD",
    x"1189BA6",
    x"118997F",
    x"1189759",
    x"1189534",
    x"118930F",
    x"11890EA",
    x"1188EC6",
    x"1188CA3",
    x"1188A80",
    x"118885E",
    x"118863C",
    x"118841A",
    x"11881FA",
    x"1187FD9",
    x"1187DBA",
    x"1187B9B",
    x"118797C",
    x"118775E",
    x"1187540",
    x"1187323",
    x"1187107",
    x"1186EEB",
    x"1186CCF",
    x"1186AB4",
    x"118689A",
    x"1186680",
    x"1186467",
    x"118624E",
    x"1186035",
    x"1185E1E",
    x"1185C06",
    x"11859F0",
    x"11857D9",
    x"11855C4",
    x"11853AF",
    x"118519A",
    x"1184F86",
    x"1184D72",
    x"1184B5F",
    x"118494C",
    x"118473A",
    x"1184529",
    x"1184318",
    x"1184107",
    x"1183EF7",
    x"1183CE8",
    x"1183AD9",
    x"11838CA",
    x"11836BC",
    x"11834AF",
    x"11832A2",
    x"1183096",
    x"1182E8A",
    x"1182C7E",
    x"1182A74",
    x"1182869",
    x"118265F",
    x"1182456",
    x"118224D",
    x"1182045",
    x"1181E3D",
    x"1181C36",
    x"1181A2F",
    x"1181829",
    x"1181623",
    x"118141E",
    x"1181219",
    x"1181015",
    x"1180E11",
    x"1180C0D",
    x"1180A0B",
    x"1180808",
    x"1180607",
    x"1180405",
    x"1180205",
    x"1180004",
    x"117FC0A",
    x"117F80B",
    x"117F40E",
    x"117F011",
    x"117EC16",
    x"117E81B",
    x"117E422",
    x"117E029",
    x"117DC32",
    x"117D83B",
    x"117D446",
    x"117D051",
    x"117CC5D",
    x"117C86B",
    x"117C479",
    x"117C089",
    x"117BC99",
    x"117B8AA",
    x"117B4BD",
    x"117B0D0",
    x"117ACE4",
    x"117A8F9",
    x"117A510",
    x"117A127",
    x"1179D3F",
    x"1179958",
    x"1179572",
    x"117918E",
    x"1178DAA",
    x"11789C7",
    x"11785E5",
    x"1178204",
    x"1177E24",
    x"1177A45",
    x"1177667",
    x"1177289",
    x"1176EAD",
    x"1176AD2",
    x"11766F8",
    x"117631F",
    x"1175F46",
    x"1175B6F",
    x"1175799",
    x"11753C3",
    x"1174FEF",
    x"1174C1B",
    x"1174849",
    x"1174477",
    x"11740A6",
    x"1173CD7",
    x"1173908",
    x"117353A",
    x"117316D",
    x"1172DA2",
    x"11729D7",
    x"117260D",
    x"1172244",
    x"1171E7B",
    x"1171AB4",
    x"11716EE",
    x"1171329",
    x"1170F65",
    x"1170BA1",
    x"11707DF",
    x"117041D",
    x"117005D",
    x"116FC9D",
    x"116F8DE",
    x"116F521",
    x"116F164",
    x"116EDA8",
    x"116E9ED",
    x"116E633",
    x"116E27A",
    x"116DEC2",
    x"116DB0B",
    x"116D754",
    x"116D39F",
    x"116CFEA",
    x"116CC37",
    x"116C884",
    x"116C4D3",
    x"116C122",
    x"116BD72",
    x"116B9C3",
    x"116B615",
    x"116B268",
    x"116AEBC",
    x"116AB11",
    x"116A766",
    x"116A3BD",
    x"116A015",
    x"1169C6D",
    x"11698C6",
    x"1169521",
    x"116917C",
    x"1168DD8",
    x"1168A35",
    x"1168693",
    x"11682F2",
    x"1167F51",
    x"1167BB2",
    x"1167813",
    x"1167476",
    x"11670D9",
    x"1166D3D",
    x"11669A3",
    x"1166609",
    x"1166270",
    x"1165ED7",
    x"1165B40",
    x"11657AA",
    x"1165414",
    x"1165080",
    x"1164CEC",
    x"1164959",
    x"11645C7",
    x"1164236",
    x"1163EA6",
    x"1163B17",
    x"1163789",
    x"11633FB",
    x"116306F",
    x"1162CE3",
    x"1162958",
    x"11625CE",
    x"1162245",
    x"1161EBD",
    x"1161B36",
    x"11617B0",
    x"116142A",
    x"11610A6",
    x"1160D22",
    x"116099F",
    x"116061D",
    x"116029C",
    x"115FF1C",
    x"115FB9C",
    x"115F81E",
    x"115F4A0",
    x"115F124",
    x"115EDA8",
    x"115EA2D",
    x"115E6B3",
    x"115E339",
    x"115DFC1",
    x"115DC4A",
    x"115D8D3",
    x"115D55D",
    x"115D1E8",
    x"115CE74",
    x"115CB01",
    x"115C78F",
    x"115C41D",
    x"115C0AD",
    x"115BD3D",
    x"115B9CE",
    x"115B660",
    x"115B2F3",
    x"115AF87",
    x"115AC1B",
    x"115A8B0",
    x"115A547",
    x"115A1DE",
    x"1159E76",
    x"1159B0F",
    x"11597A8",
    x"1159443",
    x"11590DE",
    x"1158D7A",
    x"1158A17",
    x"11586B5",
    x"1158354",
    x"1157FF4",
    x"1157C94",
    x"1157935",
    x"11575D7",
    x"115727A",
    x"1156F1E",
    x"1156BC3",
    x"1156868",
    x"115650F",
    x"11561B6",
    x"1155E5E",
    x"1155B07",
    x"11557B0",
    x"115545B",
    x"1155106",
    x"1154DB2",
    x"1154A5F",
    x"115470D",
    x"11543BC",
    x"115406B",
    x"1153D1B",
    x"11539CD",
    x"115367F",
    x"1153331",
    x"1152FE5",
    x"1152C99",
    x"115294F",
    x"1152605",
    x"11522BC",
    x"1151F73",
    x"1151C2C",
    x"11518E5",
    x"11515A0",
    x"115125B",
    x"1150F16",
    x"1150BD3",
    x"1150890",
    x"115054F",
    x"115020E",
    x"114FECE",
    x"114FB8E",
    x"114F850",
    x"114F512",
    x"114F1D5",
    x"114EE99",
    x"114EB5E",
    x"114E824",
    x"114E4EA",
    x"114E1B1",
    x"114DE79",
    x"114DB42",
    x"114D80B",
    x"114D4D6",
    x"114D1A1",
    x"114CE6D",
    x"114CB3A",
    x"114C807",
    x"114C4D6",
    x"114C1A5",
    x"114BE75",
    x"114BB46",
    x"0000000"
