library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity exponential_rom is
  port
  (
    clk       : in  std_logic;
    address   : in  std_logic_vector(15 downto 0);
    data_out  : out std_logic_vector(31 downto 0)
  );
end entity;

architecture rtl of exponential_rom is

  constant C_DATA_WIDTH  : integer := 32;
  constant C_ADDR_WIDTH  : integer := 16;

  constant RAM_DEPTH :integer := 2**C_ADDR_WIDTH;

  type RAM is array (integer range <>) of std_logic_vector (C_DATA_WIDTH-1 downto 0);
  signal mem : RAM (0 to RAM_DEPTH-1) :=
  (
    x"3F800000",
    x"3F7F9C14",
    x"3F7F384E",
    x"3F7ED4B0",
    x"3F7E7138",
    x"3F7E0DE7",
    x"3F7DAABD",
    x"3F7D47BA",
    x"3F7CE4DD",
    x"3F7C8227",
    x"3F7C1F97",
    x"3F7BBD2E",
    x"3F7B5AEB",
    x"3F7AF8CF",
    x"3F7A96D9",
    x"3F7A3509",
    x"3F79D360",
    x"3F7971DC",
    x"3F79107F",
    x"3F78AF47",
    x"3F784E36",
    x"3F77ED4A",
    x"3F778C84",
    x"3F772BE4",
    x"3F76CB6A",
    x"3F766B15",
    x"3F760AE6",
    x"3F75AADD",
    x"3F754AF9",
    x"3F74EB3A",
    x"3F748BA1",
    x"3F742C2D",
    x"3F73CCDE",
    x"3F736DB5",
    x"3F730EB1",
    x"3F72AFD1",
    x"3F725117",
    x"3F71F282",
    x"3F719412",
    x"3F7135C6",
    x"3F70D7A0",
    x"3F70799E",
    x"3F701BC1",
    x"3F6FBE08",
    x"3F6F6074",
    x"3F6F0305",
    x"3F6EA5BA",
    x"3F6E4893",
    x"3F6DEB91",
    x"3F6D8EB3",
    x"3F6D31FA",
    x"3F6CD564",
    x"3F6C78F3",
    x"3F6C1CA6",
    x"3F6BC07D",
    x"3F6B6477",
    x"3F6B0896",
    x"3F6AACD9",
    x"3F6A513F",
    x"3F69F5C9",
    x"3F699A77",
    x"3F693F48",
    x"3F68E43E",
    x"3F688956",
    x"3F682E92",
    x"3F67D3F2",
    x"3F677975",
    x"3F671F1B",
    x"3F66C4E4",
    x"3F666AD1",
    x"3F6610E1",
    x"3F65B714",
    x"3F655D6A",
    x"3F6503E3",
    x"3F64AA7F",
    x"3F64513E",
    x"3F63F81F",
    x"3F639F24",
    x"3F63464B",
    x"3F62ED95",
    x"3F629501",
    x"3F623C90",
    x"3F61E442",
    x"3F618C16",
    x"3F61340C",
    x"3F60DC25",
    x"3F608460",
    x"3F602CBE",
    x"3F5FD53D",
    x"3F5F7DDF",
    x"3F5F26A3",
    x"3F5ECF89",
    x"3F5E7891",
    x"3F5E21BB",
    x"3F5DCB07",
    x"3F5D7474",
    x"3F5D1E04",
    x"3F5CC7B5",
    x"3F5C7188",
    x"3F5C1B7C",
    x"3F5BC592",
    x"3F5B6FCA",
    x"3F5B1A23",
    x"3F5AC49D",
    x"3F5A6F39",
    x"3F5A19F6",
    x"3F59C4D5",
    x"3F596FD5",
    x"3F591AF5",
    x"3F58C637",
    x"3F58719B",
    x"3F581D1F",
    x"3F57C8C4",
    x"3F57748A",
    x"3F572071",
    x"3F56CC78",
    x"3F5678A1",
    x"3F5624EA",
    x"3F55D154",
    x"3F557DDF",
    x"3F552A8A",
    x"3F54D755",
    x"3F548441",
    x"3F54314E",
    x"3F53DE7B",
    x"3F538BC8",
    x"3F533936",
    x"3F52E6C4",
    x"3F529471",
    x"3F524240",
    x"3F51F02E",
    x"3F519E3C",
    x"3F514C6A",
    x"3F50FAB8",
    x"3F50A926",
    x"3F5057B4",
    x"3F500662",
    x"3F4FB52F",
    x"3F4F641C",
    x"3F4F1329",
    x"3F4EC255",
    x"3F4E71A1",
    x"3F4E210C",
    x"3F4DD097",
    x"3F4D8041",
    x"3F4D300B",
    x"3F4CDFF4",
    x"3F4C8FFC",
    x"3F4C4023",
    x"3F4BF06A",
    x"3F4BA0CF",
    x"3F4B5154",
    x"3F4B01F8",
    x"3F4AB2BB",
    x"3F4A639C",
    x"3F4A149D",
    x"3F49C5BC",
    x"3F4976FA",
    x"3F492857",
    x"3F48D9D3",
    x"3F488B6D",
    x"3F483D26",
    x"3F47EEFD",
    x"3F47A0F3",
    x"3F475307",
    x"3F47053A",
    x"3F46B78B",
    x"3F4669FB",
    x"3F461C88",
    x"3F45CF34",
    x"3F4581FF",
    x"3F4534E7",
    x"3F44E7ED",
    x"3F449B12",
    x"3F444E54",
    x"3F4401B4",
    x"3F43B533",
    x"3F4368CF",
    x"3F431C89",
    x"3F42D061",
    x"3F428456",
    x"3F423869",
    x"3F41EC9A",
    x"3F41A0E8",
    x"3F415554",
    x"3F4109DE",
    x"3F40BE84",
    x"3F407349",
    x"3F40282A",
    x"3F3FDD29",
    x"3F3F9246",
    x"3F3F477F",
    x"3F3EFCD6",
    x"3F3EB24A",
    x"3F3E67DA",
    x"3F3E1D88",
    x"3F3DD353",
    x"3F3D893B",
    x"3F3D3F40",
    x"3F3CF562",
    x"3F3CABA0",
    x"3F3C61FC",
    x"3F3C1874",
    x"3F3BCF09",
    x"3F3B85BA",
    x"3F3B3C88",
    x"3F3AF373",
    x"3F3AAA7A",
    x"3F3A619E",
    x"3F3A18DE",
    x"3F39D03A",
    x"3F3987B3",
    x"3F393F48",
    x"3F38F6FA",
    x"3F38AEC7",
    x"3F3866B1",
    x"3F381EB7",
    x"3F37D6D9",
    x"3F378F17",
    x"3F374771",
    x"3F36FFE7",
    x"3F36B879",
    x"3F367127",
    x"3F3629F1",
    x"3F35E2D6",
    x"3F359BD8",
    x"3F3554F5",
    x"3F350E2D",
    x"3F34C781",
    x"3F3480F1",
    x"3F343A7D",
    x"3F33F424",
    x"3F33ADE6",
    x"3F3367C4",
    x"3F3321BD",
    x"3F32DBD1",
    x"3F329601",
    x"3F32504C",
    x"3F320AB2",
    x"3F31C534",
    x"3F317FD0",
    x"3F313A88",
    x"3F30F55B",
    x"3F30B048",
    x"3F306B51",
    x"3F302674",
    x"3F2FE1B3",
    x"3F2F9D0C",
    x"3F2F5880",
    x"3F2F140F",
    x"3F2ECFB8",
    x"3F2E8B7D",
    x"3F2E475B",
    x"3F2E0355",
    x"3F2DBF69",
    x"3F2D7B97",
    x"3F2D37E0",
    x"3F2CF444",
    x"3F2CB0C1",
    x"3F2C6D59",
    x"3F2C2A0C",
    x"3F2BE6D9",
    x"3F2BA3C0",
    x"3F2B60C1",
    x"3F2B1DDC",
    x"3F2ADB11",
    x"3F2A9861",
    x"3F2A55CA",
    x"3F2A134E",
    x"3F29D0EB",
    x"3F298EA3",
    x"3F294C74",
    x"3F290A5F",
    x"3F28C864",
    x"3F288682",
    x"3F2844BB",
    x"3F28030C",
    x"3F27C178",
    x"3F277FFD",
    x"3F273E9C",
    x"3F26FD54",
    x"3F26BC26",
    x"3F267B11",
    x"3F263A16",
    x"3F25F934",
    x"3F25B86B",
    x"3F2577BC",
    x"3F253726",
    x"3F24F6A9",
    x"3F24B645",
    x"3F2475FA",
    x"3F2435C9",
    x"3F23F5B0",
    x"3F23B5B1",
    x"3F2375CA",
    x"3F2335FD",
    x"3F22F648",
    x"3F22B6AC",
    x"3F22772A",
    x"3F2237BF",
    x"3F21F86E",
    x"3F21B935",
    x"3F217A15",
    x"3F213B0E",
    x"3F20FC1F",
    x"3F20BD49",
    x"3F207E8B",
    x"3F203FE6",
    x"3F200159",
    x"3F1FC2E5",
    x"3F1F8489",
    x"3F1F4645",
    x"3F1F081A",
    x"3F1ECA07",
    x"3F1E8C0C",
    x"3F1E4E2A",
    x"3F1E105F",
    x"3F1DD2AD",
    x"3F1D9513",
    x"3F1D5790",
    x"3F1D1A26",
    x"3F1CDCD4",
    x"3F1C9F9A",
    x"3F1C6277",
    x"3F1C256D",
    x"3F1BE87A",
    x"3F1BAB9F",
    x"3F1B6EDC",
    x"3F1B3230",
    x"3F1AF59D",
    x"3F1AB921",
    x"3F1A7CBC",
    x"3F1A406F",
    x"3F1A043A",
    x"3F19C81C",
    x"3F198C15",
    x"3F195026",
    x"3F19144F",
    x"3F18D88E",
    x"3F189CE5",
    x"3F186154",
    x"3F1825D9",
    x"3F17EA76",
    x"3F17AF2A",
    x"3F1773F5",
    x"3F1738D8",
    x"3F16FDD1",
    x"3F16C2E1",
    x"3F168809",
    x"3F164D47",
    x"3F16129C",
    x"3F15D808",
    x"3F159D8C",
    x"3F156325",
    x"3F1528D6",
    x"3F14EE9D",
    x"3F14B47C",
    x"3F147A70",
    x"3F14407C",
    x"3F14069E",
    x"3F13CCD7",
    x"3F139326",
    x"3F13598C",
    x"3F132008",
    x"3F12E69B",
    x"3F12AD44",
    x"3F127403",
    x"3F123AD9",
    x"3F1201C5",
    x"3F11C8C8",
    x"3F118FE1",
    x"3F11570F",
    x"3F111E55",
    x"3F10E5B0",
    x"3F10AD21",
    x"3F1074A8",
    x"3F103C46",
    x"3F1003F9",
    x"3F0FCBC3",
    x"3F0F93A2",
    x"3F0F5B97",
    x"3F0F23A3",
    x"3F0EEBC4",
    x"3F0EB3FA",
    x"3F0E7C47",
    x"3F0E44A9",
    x"3F0E0D21",
    x"3F0DD5AF",
    x"3F0D9E52",
    x"3F0D670B",
    x"3F0D2FDA",
    x"3F0CF8BE",
    x"3F0CC1B8",
    x"3F0C8AC7",
    x"3F0C53EB",
    x"3F0C1D25",
    x"3F0BE674",
    x"3F0BAFD9",
    x"3F0B7953",
    x"3F0B42E2",
    x"3F0B0C87",
    x"3F0AD640",
    x"3F0AA00F",
    x"3F0A69F3",
    x"3F0A33EC",
    x"3F09FDFB",
    x"3F09C81E",
    x"3F099256",
    x"3F095CA4",
    x"3F092706",
    x"3F08F17D",
    x"3F08BC09",
    x"3F0886AA",
    x"3F085160",
    x"3F081C2B",
    x"3F07E70A",
    x"3F07B1FE",
    x"3F077D07",
    x"3F074825",
    x"3F071357",
    x"3F06DE9D",
    x"3F06A9F9",
    x"3F067569",
    x"3F0640ED",
    x"3F060C86",
    x"3F05D833",
    x"3F05A3F5",
    x"3F056FCB",
    x"3F053BB6",
    x"3F0507B4",
    x"3F04D3C8",
    x"3F049FEF",
    x"3F046C2B",
    x"3F04387A",
    x"3F0404DE",
    x"3F03D157",
    x"3F039DE3",
    x"3F036A83",
    x"3F033738",
    x"3F030400",
    x"3F02D0DD",
    x"3F029DCD",
    x"3F026AD1",
    x"3F0237E9",
    x"3F020516",
    x"3F01D255",
    x"3F019FA9",
    x"3F016D11",
    x"3F013A8C",
    x"3F01081B",
    x"3F00D5BE",
    x"3F00A374",
    x"3F00713E",
    x"3F003F1C",
    x"3F000D0D",
    x"3EFFB623",
    x"3EFF5253",
    x"3EFEEEAA",
    x"3EFE8B29",
    x"3EFE27CE",
    x"3EFDC499",
    x"3EFD618C",
    x"3EFCFEA5",
    x"3EFC9BE5",
    x"3EFC394B",
    x"3EFBD6D8",
    x"3EFB748B",
    x"3EFB1265",
    x"3EFAB065",
    x"3EFA4E8B",
    x"3EF9ECD8",
    x"3EF98B4A",
    x"3EF929E3",
    x"3EF8C8A2",
    x"3EF86786",
    x"3EF80691",
    x"3EF7A5C1",
    x"3EF74517",
    x"3EF6E493",
    x"3EF68435",
    x"3EF623FC",
    x"3EF5C3E8",
    x"3EF563FB",
    x"3EF50432",
    x"3EF4A48F",
    x"3EF44512",
    x"3EF3E5B9",
    x"3EF38686",
    x"3EF32778",
    x"3EF2C88F",
    x"3EF269CB",
    x"3EF20B2D",
    x"3EF1ACB3",
    x"3EF14E5E",
    x"3EF0F02E",
    x"3EF09222",
    x"3EF0343B",
    x"3EEFD679",
    x"3EEF78DC",
    x"3EEF1B63",
    x"3EEEBE0E",
    x"3EEE60DE",
    x"3EEE03D3",
    x"3EEDA6EB",
    x"3EED4A28",
    x"3EECED89",
    x"3EEC910F",
    x"3EEC34B8",
    x"3EEBD885",
    x"3EEB7C77",
    x"3EEB208C",
    x"3EEAC4C5",
    x"3EEA6922",
    x"3EEA0DA3",
    x"3EE9B248",
    x"3EE95710",
    x"3EE8FBFC",
    x"3EE8A10B",
    x"3EE8463E",
    x"3EE7EB94",
    x"3EE7910E",
    x"3EE736AB",
    x"3EE6DC6B",
    x"3EE6824F",
    x"3EE62855",
    x"3EE5CE7F",
    x"3EE574CC",
    x"3EE51B3C",
    x"3EE4C1CF",
    x"3EE46884",
    x"3EE40F5D",
    x"3EE3B658",
    x"3EE35D76",
    x"3EE304B7",
    x"3EE2AC1B",
    x"3EE253A1",
    x"3EE1FB49",
    x"3EE1A314",
    x"3EE14B02",
    x"3EE0F312",
    x"3EE09B44",
    x"3EE04399",
    x"3EDFEC0F",
    x"3EDF94A8",
    x"3EDF3D63",
    x"3EDEE640",
    x"3EDE8F3F",
    x"3EDE3860",
    x"3EDDE1A3",
    x"3EDD8B08",
    x"3EDD348E",
    x"3EDCDE37",
    x"3EDC8801",
    x"3EDC31ED",
    x"3EDBDBFA",
    x"3EDB8629",
    x"3EDB3079",
    x"3EDADAEB",
    x"3EDA857E",
    x"3EDA3032",
    x"3ED9DB08",
    x"3ED985FF",
    x"3ED93118",
    x"3ED8DC51",
    x"3ED887AB",
    x"3ED83327",
    x"3ED7DEC3",
    x"3ED78A81",
    x"3ED7365F",
    x"3ED6E25E",
    x"3ED68E7E",
    x"3ED63ABF",
    x"3ED5E720",
    x"3ED593A3",
    x"3ED54045",
    x"3ED4ED08",
    x"3ED499EC",
    x"3ED446F0",
    x"3ED3F414",
    x"3ED3A159",
    x"3ED34EBE",
    x"3ED2FC44",
    x"3ED2A9E9",
    x"3ED257AF",
    x"3ED20595",
    x"3ED1B39B",
    x"3ED161C0",
    x"3ED11006",
    x"3ED0BE6C",
    x"3ED06CF1",
    x"3ED01B97",
    x"3ECFCA5C",
    x"3ECF7941",
    x"3ECF2845",
    x"3ECED769",
    x"3ECE86AD",
    x"3ECE3610",
    x"3ECDE593",
    x"3ECD9535",
    x"3ECD44F6",
    x"3ECCF4D7",
    x"3ECCA4D7",
    x"3ECC54F6",
    x"3ECC0534",
    x"3ECBB592",
    x"3ECB660E",
    x"3ECB16AA",
    x"3ECAC765",
    x"3ECA783E",
    x"3ECA2937",
    x"3EC9DA4E",
    x"3EC98B84",
    x"3EC93CD9",
    x"3EC8EE4D",
    x"3EC89FDF",
    x"3EC85190",
    x"3EC8035F",
    x"3EC7B54D",
    x"3EC7675A",
    x"3EC71984",
    x"3EC6CBCE",
    x"3EC67E35",
    x"3EC630BB",
    x"3EC5E35F",
    x"3EC59621",
    x"3EC54902",
    x"3EC4FC00",
    x"3EC4AF1D",
    x"3EC46257",
    x"3EC415B0",
    x"3EC3C926",
    x"3EC37CBB",
    x"3EC3306D",
    x"3EC2E43D",
    x"3EC2982B",
    x"3EC24C36",
    x"3EC2005F",
    x"3EC1B4A6",
    x"3EC1690A",
    x"3EC11D8C",
    x"3EC0D22B",
    x"3EC086E7",
    x"3EC03BC1",
    x"3EBFF0B9",
    x"3EBFA5CD",
    x"3EBF5AFF",
    x"3EBF104E",
    x"3EBEC5BA",
    x"3EBE7B44",
    x"3EBE30EA",
    x"3EBDE6AE",
    x"3EBD9C8E",
    x"3EBD528B",
    x"3EBD08A5",
    x"3EBCBEDC",
    x"3EBC7530",
    x"3EBC2BA1",
    x"3EBBE22E",
    x"3EBB98D8",
    x"3EBB4F9F",
    x"3EBB0682",
    x"3EBABD82",
    x"3EBA749E",
    x"3EBA2BD7",
    x"3EB9E32C",
    x"3EB99A9D",
    x"3EB9522B",
    x"3EB909D5",
    x"3EB8C19B",
    x"3EB8797E",
    x"3EB8317C",
    x"3EB7E997",
    x"3EB7A1CE",
    x"3EB75A21",
    x"3EB7128F",
    x"3EB6CB1A",
    x"3EB683C1",
    x"3EB63C83",
    x"3EB5F561",
    x"3EB5AE5B",
    x"3EB56771",
    x"3EB520A2",
    x"3EB4D9F0",
    x"3EB49358",
    x"3EB44CDC",
    x"3EB4067C",
    x"3EB3C037",
    x"3EB37A0E",
    x"3EB33400",
    x"3EB2EE0D",
    x"3EB2A836",
    x"3EB2627A",
    x"3EB21CD9",
    x"3EB1D753",
    x"3EB191E9",
    x"3EB14C99",
    x"3EB10765",
    x"3EB0C24C",
    x"3EB07D4D",
    x"3EB0386A",
    x"3EAFF3A1",
    x"3EAFAEF3",
    x"3EAF6A60",
    x"3EAF25E8",
    x"3EAEE18B",
    x"3EAE9D48",
    x"3EAE5920",
    x"3EAE1512",
    x"3EADD11F",
    x"3EAD8D47",
    x"3EAD4989",
    x"3EAD05E5",
    x"3EACC25C",
    x"3EAC7EEE",
    x"3EAC3B99",
    x"3EABF85F",
    x"3EABB53F",
    x"3EAB7239",
    x"3EAB2F4E",
    x"3EAAEC7C",
    x"3EAAA9C5",
    x"3EAA6728",
    x"3EAA24A5",
    x"3EA9E23B",
    x"3EA99FEC",
    x"3EA95DB6",
    x"3EA91B9B",
    x"3EA8D999",
    x"3EA897B1",
    x"3EA855E2",
    x"3EA8142D",
    x"3EA7D292",
    x"3EA79111",
    x"3EA74FA9",
    x"3EA70E5B",
    x"3EA6CD26",
    x"3EA68C0A",
    x"3EA64B08",
    x"3EA60A20",
    x"3EA5C950",
    x"3EA5889A",
    x"3EA547FE",
    x"3EA5077A",
    x"3EA4C710",
    x"3EA486BF",
    x"3EA44687",
    x"3EA40668",
    x"3EA3C662",
    x"3EA38675",
    x"3EA346A0",
    x"3EA306E5",
    x"3EA2C743",
    x"3EA287BA",
    x"3EA24849",
    x"3EA208F1",
    x"3EA1C9B2",
    x"3EA18A8C",
    x"3EA14B7E",
    x"3EA10C89",
    x"3EA0CDAC",
    x"3EA08EE8",
    x"3EA0503C",
    x"3EA011A9",
    x"3E9FD32F",
    x"3E9F94CC",
    x"3E9F5682",
    x"3E9F1851",
    x"3E9EDA37",
    x"3E9E9C36",
    x"3E9E5E4D",
    x"3E9E207C",
    x"3E9DE2C4",
    x"3E9DA523",
    x"3E9D679B",
    x"3E9D2A2A",
    x"3E9CECD2",
    x"3E9CAF91",
    x"3E9C7269",
    x"3E9C3558",
    x"3E9BF85F",
    x"3E9BBB7E",
    x"3E9B7EB4",
    x"3E9B4203",
    x"3E9B0569",
    x"3E9AC8E7",
    x"3E9A8C7C",
    x"3E9A5029",
    x"3E9A13ED",
    x"3E99D7C9",
    x"3E999BBD",
    x"3E995FC8",
    x"3E9923EA",
    x"3E98E824",
    x"3E98AC74",
    x"3E9870DD",
    x"3E98355C",
    x"3E97F9F3",
    x"3E97BEA1",
    x"3E978366",
    x"3E974842",
    x"3E970D36",
    x"3E96D240",
    x"3E969761",
    x"3E965C9A",
    x"3E9621E9",
    x"3E95E74F",
    x"3E95ACCC",
    x"3E957260",
    x"3E95380B",
    x"3E94FDCC",
    x"3E94C3A5",
    x"3E948994",
    x"3E944F99",
    x"3E9415B5",
    x"3E93DBE8",
    x"3E93A232",
    x"3E936891",
    x"3E932F08",
    x"3E92F595",
    x"3E92BC38",
    x"3E9282F2",
    x"3E9249C2",
    x"3E9210A8",
    x"3E91D7A5",
    x"3E919EB8",
    x"3E9165E1",
    x"3E912D20",
    x"3E90F475",
    x"3E90BBE1",
    x"3E908363",
    x"3E904AFA",
    x"3E9012A8",
    x"3E8FDA6C",
    x"3E8FA245",
    x"3E8F6A35",
    x"3E8F323A",
    x"3E8EFA56",
    x"3E8EC287",
    x"3E8E8ACE",
    x"3E8E532A",
    x"3E8E1B9D",
    x"3E8DE425",
    x"3E8DACC2",
    x"3E8D7576",
    x"3E8D3E3F",
    x"3E8D071D",
    x"3E8CD011",
    x"3E8C991B",
    x"3E8C6239",
    x"3E8C2B6E",
    x"3E8BF4B8",
    x"3E8BBE17",
    x"3E8B878B",
    x"3E8B5115",
    x"3E8B1AB4",
    x"3E8AE468",
    x"3E8AAE31",
    x"3E8A7810",
    x"3E8A4203",
    x"3E8A0C0C",
    x"3E89D62A",
    x"3E89A05D",
    x"3E896AA5",
    x"3E893501",
    x"3E88FF73",
    x"3E88C9FA",
    x"3E889495",
    x"3E885F46",
    x"3E882A0B",
    x"3E87F4E5",
    x"3E87BFD4",
    x"3E878AD7",
    x"3E8755EF",
    x"3E87211C",
    x"3E86EC5D",
    x"3E86B7B3",
    x"3E86831E",
    x"3E864E9D",
    x"3E861A30",
    x"3E85E5D8",
    x"3E85B195",
    x"3E857D66",
    x"3E85494B",
    x"3E851544",
    x"3E84E152",
    x"3E84AD74",
    x"3E8479AB",
    x"3E8445F5",
    x"3E841254",
    x"3E83DEC7",
    x"3E83AB4E",
    x"3E8377E9",
    x"3E834498",
    x"3E83115B",
    x"3E82DE33",
    x"3E82AB1E",
    x"3E82781D",
    x"3E824530",
    x"3E821257",
    x"3E81DF92",
    x"3E81ACE0",
    x"3E817A43",
    x"3E8147B9",
    x"3E811543",
    x"3E80E2E0",
    x"3E80B091",
    x"3E807E56",
    x"3E804C2F",
    x"3E801A1B",
    x"3E7FD034",
    x"3E7F6C5B",
    x"3E7F08A8",
    x"3E7EA51C",
    x"3E7E41B7",
    x"3E7DDE78",
    x"3E7D7B61",
    x"3E7D1870",
    x"3E7CB5A6",
    x"3E7C5302",
    x"3E7BF085",
    x"3E7B8E2E",
    x"3E7B2BFE",
    x"3E7AC9F4",
    x"3E7A6810",
    x"3E7A0652",
    x"3E79A4BB",
    x"3E79434A",
    x"3E78E1FE",
    x"3E7880D9",
    x"3E781FDA",
    x"3E77BF00",
    x"3E775E4D",
    x"3E76FDBF",
    x"3E769D56",
    x"3E763D14",
    x"3E75DCF7",
    x"3E757CFF",
    x"3E751D2D",
    x"3E74BD80",
    x"3E745DF9",
    x"3E73FE97",
    x"3E739F5A",
    x"3E734042",
    x"3E72E150",
    x"3E728282",
    x"3E7223DA",
    x"3E71C556",
    x"3E7166F8",
    x"3E7108BE",
    x"3E70AAA9",
    x"3E704CB8",
    x"3E6FEEED",
    x"3E6F9146",
    x"3E6F33C3",
    x"3E6ED665",
    x"3E6E792C",
    x"3E6E1C17",
    x"3E6DBF26",
    x"3E6D6259",
    x"3E6D05B1",
    x"3E6CA92D",
    x"3E6C4CCD",
    x"3E6BF091",
    x"3E6B9479",
    x"3E6B3885",
    x"3E6ADCB5",
    x"3E6A8108",
    x"3E6A2580",
    x"3E69CA1B",
    x"3E696EDA",
    x"3E6913BC",
    x"3E68B8C2",
    x"3E685DEC",
    x"3E680339",
    x"3E67A8A9",
    x"3E674E3D",
    x"3E66F3F4",
    x"3E6699CF",
    x"3E663FCC",
    x"3E65E5ED",
    x"3E658C30",
    x"3E653297",
    x"3E64D921",
    x"3E647FCE",
    x"3E64269D",
    x"3E63CD8F",
    x"3E6374A4",
    x"3E631BDC",
    x"3E62C337",
    x"3E626AB4",
    x"3E621253",
    x"3E61BA15",
    x"3E6161FA",
    x"3E610A01",
    x"3E60B22A",
    x"3E605A76",
    x"3E6002E3",
    x"3E5FAB73",
    x"3E5F5425",
    x"3E5EFCFA",
    x"3E5EA5F0",
    x"3E5E4F08",
    x"3E5DF842",
    x"3E5DA19E",
    x"3E5D4B1C",
    x"3E5CF4BB",
    x"3E5C9E7C",
    x"3E5C485F",
    x"3E5BF264",
    x"3E5B9C8A",
    x"3E5B46D2",
    x"3E5AF13B",
    x"3E5A9BC5",
    x"3E5A4671",
    x"3E59F13E",
    x"3E599C2C",
    x"3E59473C",
    x"3E58F26D",
    x"3E589DBF",
    x"3E584932",
    x"3E57F4C5",
    x"3E57A07A",
    x"3E574C50",
    x"3E56F847",
    x"3E56A45E",
    x"3E565096",
    x"3E55FCEF",
    x"3E55A969",
    x"3E555603",
    x"3E5502BD",
    x"3E54AF99",
    x"3E545C94",
    x"3E5409B0",
    x"3E53B6ED",
    x"3E536449",
    x"3E5311C6",
    x"3E52BF63",
    x"3E526D21",
    x"3E521AFE",
    x"3E51C8FC",
    x"3E517719",
    x"3E512557",
    x"3E50D3B4",
    x"3E508231",
    x"3E5030CE",
    x"3E4FDF8B",
    x"3E4F8E68",
    x"3E4F3D64",
    x"3E4EEC80",
    x"3E4E9BBB",
    x"3E4E4B16",
    x"3E4DFA90",
    x"3E4DAA2A",
    x"3E4D59E3",
    x"3E4D09BC",
    x"3E4CB9B4",
    x"3E4C69CB",
    x"3E4C1A01",
    x"3E4BCA56",
    x"3E4B7ACB",
    x"3E4B2B5E",
    x"3E4ADC11",
    x"3E4A8CE3",
    x"3E4A3DD3",
    x"3E49EEE2",
    x"3E49A010",
    x"3E49515D",
    x"3E4902C9",
    x"3E48B453",
    x"3E4865FC",
    x"3E4817C3",
    x"3E47C9A9",
    x"3E477BAE",
    x"3E472DD1",
    x"3E46E012",
    x"3E469272",
    x"3E4644EF",
    x"3E45F78C",
    x"3E45AA46",
    x"3E455D1F",
    x"3E451015",
    x"3E44C32A",
    x"3E44765D",
    x"3E4429AE",
    x"3E43DD1C",
    x"3E4390A9",
    x"3E434453",
    x"3E42F81B",
    x"3E42AC01",
    x"3E426005",
    x"3E421426",
    x"3E41C865",
    x"3E417CC2",
    x"3E41313C",
    x"3E40E5D3",
    x"3E409A88",
    x"3E404F5B",
    x"3E40044A",
    x"3E3FB957",
    x"3E3F6E81",
    x"3E3F23C9",
    x"3E3ED92D",
    x"3E3E8EAF",
    x"3E3E444E",
    x"3E3DFA0A",
    x"3E3DAFE3",
    x"3E3D65D8",
    x"3E3D1BEB",
    x"3E3CD21B",
    x"3E3C8867",
    x"3E3C3ED0",
    x"3E3BF556",
    x"3E3BABF8",
    x"3E3B62B7",
    x"3E3B1993",
    x"3E3AD08B",
    x"3E3A87A0",
    x"3E3A3ED1",
    x"3E39F61F",
    x"3E39AD89",
    x"3E39650F",
    x"3E391CB2",
    x"3E38D471",
    x"3E388C4C",
    x"3E384443",
    x"3E37FC57",
    x"3E37B486",
    x"3E376CD2",
    x"3E372539",
    x"3E36DDBD",
    x"3E36965C",
    x"3E364F17",
    x"3E3607EE",
    x"3E35C0E1",
    x"3E3579F0",
    x"3E35331A",
    x"3E34EC60",
    x"3E34A5C1",
    x"3E345F3E",
    x"3E3418D7",
    x"3E33D28B",
    x"3E338C5A",
    x"3E334645",
    x"3E33004B",
    x"3E32BA6D",
    x"3E3274AA",
    x"3E322F02",
    x"3E31E975",
    x"3E31A403",
    x"3E315EAD",
    x"3E311971",
    x"3E30D451",
    x"3E308F4B",
    x"3E304A61",
    x"3E300591",
    x"3E2FC0DC",
    x"3E2F7C43",
    x"3E2F37C3",
    x"3E2EF35F",
    x"3E2EAF15",
    x"3E2E6AE6",
    x"3E2E26D2",
    x"3E2DE2D8",
    x"3E2D9EF8",
    x"3E2D5B34",
    x"3E2D1789",
    x"3E2CD3F9",
    x"3E2C9084",
    x"3E2C4D28",
    x"3E2C09E7",
    x"3E2BC6C1",
    x"3E2B83B4",
    x"3E2B40C2",
    x"3E2AFDE9",
    x"3E2ABB2B",
    x"3E2A7887",
    x"3E2A35FD",
    x"3E29F38D",
    x"3E29B137",
    x"3E296EFA",
    x"3E292CD8",
    x"3E28EACF",
    x"3E28A8E1",
    x"3E28670B",
    x"3E282550",
    x"3E27E3AE",
    x"3E27A226",
    x"3E2760B8",
    x"3E271F63",
    x"3E26DE27",
    x"3E269D05",
    x"3E265BFC",
    x"3E261B0D",
    x"3E25DA37",
    x"3E25997B",
    x"3E2558D7",
    x"3E25184D",
    x"3E24D7DC",
    x"3E249785",
    x"3E245746",
    x"3E241720",
    x"3E23D714",
    x"3E239720",
    x"3E235746",
    x"3E231784",
    x"3E22D7DB",
    x"3E22984C",
    x"3E2258D4",
    x"3E221976",
    x"3E21DA31",
    x"3E219B04",
    x"3E215BEF",
    x"3E211CF4",
    x"3E20DE11",
    x"3E209F46",
    x"3E206094",
    x"3E2021FB",
    x"3E1FE37A",
    x"3E1FA511",
    x"3E1F66C1",
    x"3E1F2889",
    x"3E1EEA69",
    x"3E1EAC62",
    x"3E1E6E72",
    x"3E1E309B",
    x"3E1DF2DC",
    x"3E1DB536",
    x"3E1D77A7",
    x"3E1D3A30",
    x"3E1CFCD1",
    x"3E1CBF8B",
    x"3E1C825C",
    x"3E1C4545",
    x"3E1C0846",
    x"3E1BCB5E",
    x"3E1B8E8F",
    x"3E1B51D7",
    x"3E1B1537",
    x"3E1AD8AE",
    x"3E1A9C3D",
    x"3E1A5FE4",
    x"3E1A23A3",
    x"3E19E778",
    x"3E19AB66",
    x"3E196F6A",
    x"3E193387",
    x"3E18F7BA",
    x"3E18BC05",
    x"3E188067",
    x"3E1844E1",
    x"3E180971",
    x"3E17CE19",
    x"3E1792D8",
    x"3E1757AF",
    x"3E171C9C",
    x"3E16E1A0",
    x"3E16A6BC",
    x"3E166BEE",
    x"3E163137",
    x"3E15F698",
    x"3E15BC0F",
    x"3E15819D",
    x"3E154741",
    x"3E150CFD",
    x"3E14D2CF",
    x"3E1498B8",
    x"3E145EB8",
    x"3E1424CE",
    x"3E13EAFB",
    x"3E13B13F",
    x"3E137799",
    x"3E133E09",
    x"3E130490",
    x"3E12CB2E",
    x"3E1291E1",
    x"3E1258AC",
    x"3E121F8C",
    x"3E11E683",
    x"3E11AD90",
    x"3E1174B3",
    x"3E113BED",
    x"3E11033D",
    x"3E10CAA2",
    x"3E10921E",
    x"3E1059B0",
    x"3E102158",
    x"3E0FE916",
    x"3E0FB0EA",
    x"3E0F78D4",
    x"3E0F40D4",
    x"3E0F08E9",
    x"3E0ED115",
    x"3E0E9956",
    x"3E0E61AD",
    x"3E0E2A1A",
    x"3E0DF29C",
    x"3E0DBB34",
    x"3E0D83E2",
    x"3E0D4CA5",
    x"3E0D157E",
    x"3E0CDE6C",
    x"3E0CA770",
    x"3E0C7089",
    x"3E0C39B8",
    x"3E0C02FC",
    x"3E0BCC56",
    x"3E0B95C5",
    x"3E0B5F49",
    x"3E0B28E2",
    x"3E0AF291",
    x"3E0ABC55",
    x"3E0A862E",
    x"3E0A501C",
    x"3E0A1A1F",
    x"3E09E437",
    x"3E09AE65",
    x"3E0978A7",
    x"3E0942FE",
    x"3E090D6B",
    x"3E08D7EC",
    x"3E08A282",
    x"3E086D2D",
    x"3E0837ED",
    x"3E0802C1",
    x"3E07CDAB",
    x"3E0798A9",
    x"3E0763BB",
    x"3E072EE3",
    x"3E06FA1F",
    x"3E06C56F",
    x"3E0690D4",
    x"3E065C4E",
    x"3E0627DC",
    x"3E05F37F",
    x"3E05BF36",
    x"3E058B02",
    x"3E0556E1",
    x"3E0522D6",
    x"3E04EEDE",
    x"3E04BAFB",
    x"3E04872C",
    x"3E045371",
    x"3E041FCB",
    x"3E03EC39",
    x"3E03B8BA",
    x"3E038550",
    x"3E0351FA",
    x"3E031EB8",
    x"3E02EB8A",
    x"3E02B870",
    x"3E02856A",
    x"3E025278",
    x"3E021F9A",
    x"3E01ECCF",
    x"3E01BA19",
    x"3E018776",
    x"3E0154E7",
    x"3E01226B",
    x"3E00F004",
    x"3E00BDB0",
    x"3E008B70",
    x"3E005943",
    x"3E00272A",
    x"3DFFEA49",
    x"3DFF8665",
    x"3DFF22A8",
    x"3DFEBF12",
    x"3DFE5BA3",
    x"3DFDF85A",
    x"3DFD9538",
    x"3DFD323E",
    x"3DFCCF69",
    x"3DFC6CBB",
    x"3DFC0A34",
    x"3DFBA7D3",
    x"3DFB4599",
    x"3DFAE385",
    x"3DFA8197",
    x"3DFA1FD0",
    x"3DF9BE2E",
    x"3DF95CB3",
    x"3DF8FB5E",
    x"3DF89A2F",
    x"3DF83926",
    x"3DF7D842",
    x"3DF77785",
    x"3DF716ED",
    x"3DF6B67B",
    x"3DF6562E",
    x"3DF5F607",
    x"3DF59606",
    x"3DF5362A",
    x"3DF4D674",
    x"3DF476E3",
    x"3DF41777",
    x"3DF3B830",
    x"3DF3590F",
    x"3DF2FA13",
    x"3DF29B3B",
    x"3DF23C89",
    x"3DF1DDFC",
    x"3DF17F94",
    x"3DF12150",
    x"3DF0C332",
    x"3DF06538",
    x"3DF00763",
    x"3DEFA9B2",
    x"3DEF4C26",
    x"3DEEEEBF",
    x"3DEE917C",
    x"3DEE345D",
    x"3DEDD763",
    x"3DED7A8D",
    x"3DED1DDB",
    x"3DECC14D",
    x"3DEC64E4",
    x"3DEC089E",
    x"3DEBAC7D",
    x"3DEB5080",
    x"3DEAF4A6",
    x"3DEA98F1",
    x"3DEA3D5F",
    x"3DE9E1F1",
    x"3DE986A6",
    x"3DE92B7F",
    x"3DE8D07C",
    x"3DE8759C",
    x"3DE81AE0",
    x"3DE7C047",
    x"3DE765D2",
    x"3DE70B80",
    x"3DE6B151",
    x"3DE65745",
    x"3DE5FD5D",
    x"3DE5A397",
    x"3DE549F5",
    x"3DE4F076",
    x"3DE49719",
    x"3DE43DE0",
    x"3DE3E4C9",
    x"3DE38BD5",
    x"3DE33303",
    x"3DE2DA55",
    x"3DE281C9",
    x"3DE2295F",
    x"3DE1D119",
    x"3DE178F4",
    x"3DE120F2",
    x"3DE0C912",
    x"3DE07155",
    x"3DE019BA",
    x"3DDFC241",
    x"3DDF6AEA",
    x"3DDF13B5",
    x"3DDEBCA3",
    x"3DDE65B2",
    x"3DDE0EE3",
    x"3DDDB836",
    x"3DDD61AB",
    x"3DDD0B42",
    x"3DDCB4FA",
    x"3DDC5ED5",
    x"3DDC08D0",
    x"3DDBB2EE",
    x"3DDB5D2C",
    x"3DDB078D",
    x"3DDAB20F",
    x"3DDA5CB2",
    x"3DDA0776",
    x"3DD9B25C",
    x"3DD95D63",
    x"3DD9088B",
    x"3DD8B3D4",
    x"3DD85F3E",
    x"3DD80ACA",
    x"3DD7B676",
    x"3DD76243",
    x"3DD70E31",
    x"3DD6BA40",
    x"3DD66670",
    x"3DD612C0",
    x"3DD5BF31",
    x"3DD56BC3",
    x"3DD51875",
    x"3DD4C547",
    x"3DD4723B",
    x"3DD41F4E",
    x"3DD3CC82",
    x"3DD379D6",
    x"3DD3274B",
    x"3DD2D4E0",
    x"3DD28295",
    x"3DD2306A",
    x"3DD1DE5F",
    x"3DD18C74",
    x"3DD13AA9",
    x"3DD0E8FE",
    x"3DD09773",
    x"3DD04608",
    x"3DCFF4BC",
    x"3DCFA390",
    x"3DCF5284",
    x"3DCF0198",
    x"3DCEB0CB",
    x"3DCE601E",
    x"3DCE0F90",
    x"3DCDBF22",
    x"3DCD6ED3",
    x"3DCD1EA3",
    x"3DCCCE93",
    x"3DCC7EA2",
    x"3DCC2ED0",
    x"3DCBDF1D",
    x"3DCB8F8A",
    x"3DCB4015",
    x"3DCAF0BF",
    x"3DCAA189",
    x"3DCA5271",
    x"3DCA0378",
    x"3DC9B49E",
    x"3DC965E3",
    x"3DC91747",
    x"3DC8C8C9",
    x"3DC87A6A",
    x"3DC82C29",
    x"3DC7DE07",
    x"3DC79004",
    x"3DC7421F",
    x"3DC6F458",
    x"3DC6A6B0",
    x"3DC65926",
    x"3DC60BBA",
    x"3DC5BE6D",
    x"3DC5713E",
    x"3DC5242C",
    x"3DC4D739",
    x"3DC48A64",
    x"3DC43DAD",
    x"3DC3F114",
    x"3DC3A499",
    x"3DC3583B",
    x"3DC30BFC",
    x"3DC2BFDA",
    x"3DC273D6",
    x"3DC227F0",
    x"3DC1DC27",
    x"3DC1907C",
    x"3DC144EE",
    x"3DC0F97E",
    x"3DC0AE2B",
    x"3DC062F6",
    x"3DC017DE",
    x"3DBFCCE3",
    x"3DBF8206",
    x"3DBF3745",
    x"3DBEECA2",
    x"3DBEA21C",
    x"3DBE57B4",
    x"3DBE0D68",
    x"3DBDC339",
    x"3DBD7927",
    x"3DBD2F33",
    x"3DBCE55B",
    x"3DBC9B9F",
    x"3DBC5201",
    x"3DBC087F",
    x"3DBBBF1A",
    x"3DBB75D2",
    x"3DBB2CA6",
    x"3DBAE397",
    x"3DBA9AA4",
    x"3DBA51CE",
    x"3DBA0914",
    x"3DB9C077",
    x"3DB977F6",
    x"3DB92F91",
    x"3DB8E749",
    x"3DB89F1D",
    x"3DB8570D",
    x"3DB80F19",
    x"3DB7C741",
    x"3DB77F85",
    x"3DB737E5",
    x"3DB6F061",
    x"3DB6A8F9",
    x"3DB661AD",
    x"3DB61A7D",
    x"3DB5D369",
    x"3DB58C70",
    x"3DB54593",
    x"3DB4FED1",
    x"3DB4B82C",
    x"3DB471A2",
    x"3DB42B33",
    x"3DB3E4E0",
    x"3DB39EA8",
    x"3DB3588C",
    x"3DB3128B",
    x"3DB2CCA5",
    x"3DB286DB",
    x"3DB2412C",
    x"3DB1FB98",
    x"3DB1B61F",
    x"3DB170C2",
    x"3DB12B7F",
    x"3DB0E658",
    x"3DB0A14B",
    x"3DB05C5A",
    x"3DB01783",
    x"3DAFD2C7",
    x"3DAF8E26",
    x"3DAF49A0",
    x"3DAF0535",
    x"3DAEC0E4",
    x"3DAE7CAE",
    x"3DAE3893",
    x"3DADF492",
    x"3DADB0AC",
    x"3DAD6CE0",
    x"3DAD292F",
    x"3DACE598",
    x"3DACA21B",
    x"3DAC5EB9",
    x"3DAC1B71",
    x"3DABD844",
    x"3DAB9530",
    x"3DAB5237",
    x"3DAB0F58",
    x"3DAACC93",
    x"3DAA89E8",
    x"3DAA4757",
    x"3DAA04E0",
    x"3DA9C284",
    x"3DA98040",
    x"3DA93E17",
    x"3DA8FC08",
    x"3DA8BA12",
    x"3DA87837",
    x"3DA83674",
    x"3DA7F4CC",
    x"3DA7B33D",
    x"3DA771C8",
    x"3DA7306C",
    x"3DA6EF2A",
    x"3DA6AE01",
    x"3DA66CF2",
    x"3DA62BFC",
    x"3DA5EB20",
    x"3DA5AA5D",
    x"3DA569B3",
    x"3DA52922",
    x"3DA4E8AB",
    x"3DA4A84C",
    x"3DA46807",
    x"3DA427DB",
    x"3DA3E7C8",
    x"3DA3A7CE",
    x"3DA367ED",
    x"3DA32825",
    x"3DA2E875",
    x"3DA2A8DF",
    x"3DA26961",
    x"3DA229FD",
    x"3DA1EAB1",
    x"3DA1AB7D",
    x"3DA16C63",
    x"3DA12D61",
    x"3DA0EE77",
    x"3DA0AFA6",
    x"3DA070EE",
    x"3DA0324E",
    x"3D9FF3C7",
    x"3D9FB558",
    x"3D9F7701",
    x"3D9F38C3",
    x"3D9EFA9D",
    x"3D9EBC8F",
    x"3D9E7E99",
    x"3D9E40BC",
    x"3D9E02F7",
    x"3D9DC54A",
    x"3D9D87B5",
    x"3D9D4A38",
    x"3D9D0CD3",
    x"3D9CCF86",
    x"3D9C9250",
    x"3D9C5533",
    x"3D9C182E",
    x"3D9BDB40",
    x"3D9B9E6B",
    x"3D9B61AD",
    x"3D9B2506",
    x"3D9AE878",
    x"3D9AAC01",
    x"3D9A6FA1",
    x"3D9A3359",
    x"3D99F729",
    x"3D99BB10",
    x"3D997F0F",
    x"3D994325",
    x"3D990752",
    x"3D98CB97",
    x"3D988FF3",
    x"3D985467",
    x"3D9818F1",
    x"3D97DD93",
    x"3D97A24C",
    x"3D97671C",
    x"3D972C04",
    x"3D96F102",
    x"3D96B617",
    x"3D967B44",
    x"3D964087",
    x"3D9605E1",
    x"3D95CB53",
    x"3D9590DB",
    x"3D955679",
    x"3D951C2F",
    x"3D94E1FB",
    x"3D94A7DE",
    x"3D946DD8",
    x"3D9433E9",
    x"3D93FA10",
    x"3D93C04D",
    x"3D9386A1",
    x"3D934D0C",
    x"3D93138D",
    x"3D92DA25",
    x"3D92A0D3",
    x"3D926797",
    x"3D922E72",
    x"3D91F563",
    x"3D91BC6A",
    x"3D918388",
    x"3D914ABB",
    x"3D911205",
    x"3D90D965",
    x"3D90A0DB",
    x"3D906868",
    x"3D90300A",
    x"3D8FF7C2",
    x"3D8FBF90",
    x"3D8F8774",
    x"3D8F4F6E",
    x"3D8F177E",
    x"3D8EDFA4",
    x"3D8EA7E0",
    x"3D8E7031",
    x"3D8E3898",
    x"3D8E0115",
    x"3D8DC9A7",
    x"3D8D924F",
    x"3D8D5B0D",
    x"3D8D23E0",
    x"3D8CECC9",
    x"3D8CB5C7",
    x"3D8C7EDB",
    x"3D8C4804",
    x"3D8C1142",
    x"3D8BDA96",
    x"3D8BA400",
    x"3D8B6D7E",
    x"3D8B3712",
    x"3D8B00BB",
    x"3D8ACA79",
    x"3D8A944D",
    x"3D8A5E36",
    x"3D8A2833",
    x"3D89F246",
    x"3D89BC6E",
    x"3D8986AB",
    x"3D8950FD",
    x"3D891B64",
    x"3D88E5DF",
    x"3D88B070",
    x"3D887B16",
    x"3D8845D0",
    x"3D88109F",
    x"3D87DB83",
    x"3D87A67B",
    x"3D877189",
    x"3D873CAB",
    x"3D8707E1",
    x"3D86D32D",
    x"3D869E8C",
    x"3D866A01",
    x"3D86358A",
    x"3D860127",
    x"3D85CCD9",
    x"3D85989F",
    x"3D856479",
    x"3D853068",
    x"3D84FC6C",
    x"3D84C883",
    x"3D8494AF",
    x"3D8460EF",
    x"3D842D43",
    x"3D83F9AC",
    x"3D83C628",
    x"3D8392B9",
    x"3D835F5D",
    x"3D832C16",
    x"3D82F8E3",
    x"3D82C5C4",
    x"3D8292B9",
    x"3D825FC1",
    x"3D822CDE",
    x"3D81FA0E",
    x"3D81C752",
    x"3D8194AA",
    x"3D816216",
    x"3D812F96",
    x"3D80FD29",
    x"3D80CAD0",
    x"3D80988B",
    x"3D806659",
    x"3D80343B",
    x"3D800230",
    x"3D7FA072",
    x"3D7F3CAB",
    x"3D7ED90A",
    x"3D7E7591",
    x"3D7E123E",
    x"3D7DAF13",
    x"3D7D4C0E",
    x"3D7CE92F",
    x"3D7C8677",
    x"3D7C23E6",
    x"3D7BC17B",
    x"3D7B5F37",
    x"3D7AFD19",
    x"3D7A9B21",
    x"3D7A3950",
    x"3D79D7A4",
    x"3D79761F",
    x"3D7914C0",
    x"3D78B387",
    x"3D785274",
    x"3D77F187",
    x"3D7790BF",
    x"3D77301E",
    x"3D76CFA2",
    x"3D766F4B",
    x"3D760F1B",
    x"3D75AF0F",
    x"3D754F2A",
    x"3D74EF6A",
    x"3D748FCF",
    x"3D743059",
    x"3D73D109",
    x"3D7371DE",
    x"3D7312D8",
    x"3D72B3F7",
    x"3D72553B",
    x"3D71F6A5",
    x"3D719833",
    x"3D7139E6",
    x"3D70DBBD",
    x"3D707DBA",
    x"3D701FDB",
    x"3D6FC221",
    x"3D6F648B",
    x"3D6F071A",
    x"3D6EA9CE",
    x"3D6E4CA6",
    x"3D6DEFA2",
    x"3D6D92C3",
    x"3D6D3607",
    x"3D6CD970",
    x"3D6C7CFD",
    x"3D6C20AF",
    x"3D6BC484",
    x"3D6B687D",
    x"3D6B0C9A",
    x"3D6AB0DB",
    x"3D6A5540",
    x"3D69F9C9",
    x"3D699E75",
    x"3D694345",
    x"3D68E838",
    x"3D688D4F",
    x"3D68328A",
    x"3D67D7E8",
    x"3D677D69",
    x"3D67230E",
    x"3D66C8D6",
    x"3D666EC1",
    x"3D6614CF",
    x"3D65BB01",
    x"3D656155",
    x"3D6507CD",
    x"3D64AE67",
    x"3D645524",
    x"3D63FC05",
    x"3D63A307",
    x"3D634A2D",
    x"3D62F175",
    x"3D6298E0",
    x"3D62406E",
    x"3D61E81E",
    x"3D618FF1",
    x"3D6137E6",
    x"3D60DFFD",
    x"3D608837",
    x"3D603093",
    x"3D5FD911",
    x"3D5F81B1",
    x"3D5F2A73",
    x"3D5ED358",
    x"3D5E7C5E",
    x"3D5E2587",
    x"3D5DCED1",
    x"3D5D783D",
    x"3D5D21CB",
    x"3D5CCB7B",
    x"3D5C754C",
    x"3D5C1F3F",
    x"3D5BC953",
    x"3D5B738A",
    x"3D5B1DE1",
    x"3D5AC85A",
    x"3D5A72F5",
    x"3D5A1DB0",
    x"3D59C88D",
    x"3D59738C",
    x"3D591EAB",
    x"3D58C9EC",
    x"3D58754D",
    x"3D5820D0",
    x"3D57CC74",
    x"3D577838",
    x"3D57241E",
    x"3D56D024",
    x"3D567C4B",
    x"3D562893",
    x"3D55D4FB",
    x"3D558185",
    x"3D552E2E",
    x"3D54DAF8",
    x"3D5487E3",
    x"3D5434EE",
    x"3D53E21A",
    x"3D538F66",
    x"3D533CD2",
    x"3D52EA5E",
    x"3D52980B",
    x"3D5245D7",
    x"3D51F3C4",
    x"3D51A1D1",
    x"3D514FFE",
    x"3D50FE4A",
    x"3D50ACB7",
    x"3D505B43",
    x"3D5009F0",
    x"3D4FB8BC",
    x"3D4F67A7",
    x"3D4F16B3",
    x"3D4EC5DE",
    x"3D4E7528",
    x"3D4E2492",
    x"3D4DD41B",
    x"3D4D83C4",
    x"3D4D338C",
    x"3D4CE374",
    x"3D4C937B",
    x"3D4C43A1",
    x"3D4BF3E6",
    x"3D4BA44A",
    x"3D4B54CE",
    x"3D4B0570",
    x"3D4AB631",
    x"3D4A6712",
    x"3D4A1811",
    x"3D49C92F",
    x"3D497A6C",
    x"3D492BC7",
    x"3D48DD41",
    x"3D488EDA",
    x"3D484092",
    x"3D47F268",
    x"3D47A45C",
    x"3D47566F",
    x"3D4708A1",
    x"3D46BAF1",
    x"3D466D5F",
    x"3D461FEB",
    x"3D45D296",
    x"3D45855F",
    x"3D453846",
    x"3D44EB4B",
    x"3D449E6E",
    x"3D4451AF",
    x"3D44050E",
    x"3D43B88B",
    x"3D436C26",
    x"3D431FDE",
    x"3D42D3B5",
    x"3D4287A9",
    x"3D423BBB",
    x"3D41EFEA",
    x"3D41A437",
    x"3D4158A2",
    x"3D410D2A",
    x"3D40C1D0",
    x"3D407693",
    x"3D402B73",
    x"3D3FE071",
    x"3D3F958C",
    x"3D3F4AC4",
    x"3D3F0019",
    x"3D3EB58C",
    x"3D3E6B1B",
    x"3D3E20C8",
    x"3D3DD692",
    x"3D3D8C78",
    x"3D3D427C",
    x"3D3CF89C",
    x"3D3CAEDA",
    x"3D3C6534",
    x"3D3C1BAB",
    x"3D3BD23E",
    x"3D3B88EE",
    x"3D3B3FBB",
    x"3D3AF6A5",
    x"3D3AADAB",
    x"3D3A64CD",
    x"3D3A1C0C",
    x"3D39D367",
    x"3D398ADF",
    x"3D394272",
    x"3D38FA23",
    x"3D38B1EF",
    x"3D3869D8",
    x"3D3821DC",
    x"3D37D9FD",
    x"3D37923A",
    x"3D374A93",
    x"3D370308",
    x"3D36BB99",
    x"3D367445",
    x"3D362D0E",
    x"3D35E5F2",
    x"3D359EF2",
    x"3D35580E",
    x"3D351145",
    x"3D34CA98",
    x"3D348407",
    x"3D343D91",
    x"3D33F737",
    x"3D33B0F8",
    x"3D336AD5",
    x"3D3324CC",
    x"3D32DEE0",
    x"3D32990E",
    x"3D325358",
    x"3D320DBD",
    x"3D31C83D",
    x"3D3182D9",
    x"3D313D8F",
    x"3D30F861",
    x"3D30B34D",
    x"3D306E55",
    x"3D302977",
    x"3D2FE4B4",
    x"3D2FA00C",
    x"3D2F5B7F",
    x"3D2F170D",
    x"3D2ED2B5",
    x"3D2E8E78",
    x"3D2E4A56",
    x"3D2E064E",
    x"3D2DC261",
    x"3D2D7E8E",
    x"3D2D3AD6",
    x"3D2CF738",
    x"3D2CB3B5",
    x"3D2C704C",
    x"3D2C2CFD",
    x"3D2BE9C9",
    x"3D2BA6AE",
    x"3D2B63AE",
    x"3D2B20C9",
    x"3D2ADDFD",
    x"3D2A9B4B",
    x"3D2A58B3",
    x"3D2A1636",
    x"3D29D3D2",
    x"3D299188",
    x"3D294F58",
    x"3D290D42",
    x"3D28CB46",
    x"3D288963",
    x"3D28479B",
    x"3D2805EB",
    x"3D27C456",
    x"3D2782DA",
    x"3D274178",
    x"3D27002F",
    x"3D26BF00",
    x"3D267DEA",
    x"3D263CED",
    x"3D25FC0A",
    x"3D25BB40",
    x"3D257A90",
    x"3D2539F9",
    x"3D24F97A",
    x"3D24B916",
    x"3D2478CA",
    x"3D243897",
    x"3D23F87E",
    x"3D23B87D",
    x"3D237896",
    x"3D2338C7",
    x"3D22F911",
    x"3D22B974",
    x"3D2279F0",
    x"3D223A85",
    x"3D21FB33",
    x"3D21BBF9",
    x"3D217CD8",
    x"3D213DCF",
    x"3D20FEDF",
    x"3D20C008",
    x"3D208149",
    x"3D2042A3",
    x"3D200415",
    x"3D1FC5A0",
    x"3D1F8743",
    x"3D1F48FE",
    x"3D1F0AD2",
    x"3D1ECCBE",
    x"3D1E8EC2",
    x"3D1E50DE",
    x"3D1E1313",
    x"3D1DD55F",
    x"3D1D97C4",
    x"3D1D5A41",
    x"3D1D1CD5",
    x"3D1CDF82",
    x"3D1CA247",
    x"3D1C6523",
    x"3D1C2818",
    x"3D1BEB24",
    x"3D1BAE48",
    x"3D1B7184",
    x"3D1B34D7",
    x"3D1AF843",
    x"3D1ABBC5",
    x"3D1A7F60",
    x"3D1A4312",
    x"3D1A06DB",
    x"3D19CABC",
    x"3D198EB5",
    x"3D1952C5",
    x"3D1916EC",
    x"3D18DB2B",
    x"3D189F81",
    x"3D1863EE",
    x"3D182873",
    x"3D17ED0F",
    x"3D17B1C2",
    x"3D17768C",
    x"3D173B6D",
    x"3D170065",
    x"3D16C575",
    x"3D168A9B",
    x"3D164FD9",
    x"3D16152D",
    x"3D15DA98",
    x"3D15A01A",
    x"3D1565B3",
    x"3D152B63",
    x"3D14F129",
    x"3D14B706",
    x"3D147CFA",
    x"3D144305",
    x"3D140926",
    x"3D13CF5D",
    x"3D1395AC",
    x"3D135C10",
    x"3D13228C",
    x"3D12E91D",
    x"3D12AFC6",
    x"3D127684",
    x"3D123D59",
    x"3D120444",
    x"3D11CB46",
    x"3D11925D",
    x"3D11598B",
    x"3D1120CF",
    x"3D10E82A",
    x"3D10AF9A",
    x"3D107720",
    x"3D103EBD",
    x"3D10066F",
    x"3D0FCE38",
    x"3D0F9616",
    x"3D0F5E0B",
    x"3D0F2615",
    x"3D0EEE35",
    x"3D0EB66B",
    x"3D0E7EB6",
    x"3D0E4718",
    x"3D0E0F8F",
    x"3D0DD81B",
    x"3D0DA0BE",
    x"3D0D6976",
    x"3D0D3243",
    x"3D0CFB27",
    x"3D0CC41F",
    x"3D0C8D2D",
    x"3D0C5651",
    x"3D0C1F8A",
    x"3D0BE8D8",
    x"3D0BB23C",
    x"3D0B7BB5",
    x"3D0B4543",
    x"3D0B0EE7",
    x"3D0AD8A0",
    x"3D0AA26E",
    x"3D0A6C51",
    x"3D0A3649",
    x"3D0A0056",
    x"3D09CA79",
    x"3D0994B0",
    x"3D095EFD",
    x"3D09295E",
    x"3D08F3D4",
    x"3D08BE5F",
    x"3D088900",
    x"3D0853B4",
    x"3D081E7E",
    x"3D07E95D",
    x"3D07B450",
    x"3D077F58",
    x"3D074A74",
    x"3D0715A6",
    x"3D06E0EB",
    x"3D06AC46",
    x"3D0677B5",
    x"3D064338",
    x"3D060ED0",
    x"3D05DA7D",
    x"3D05A63E",
    x"3D057213",
    x"3D053DFC",
    x"3D0509FA",
    x"3D04D60D",
    x"3D04A233",
    x"3D046E6E",
    x"3D043ABD",
    x"3D040720",
    x"3D03D397",
    x"3D03A023",
    x"3D036CC2",
    x"3D033976",
    x"3D03063D",
    x"3D02D319",
    x"3D02A008",
    x"3D026D0C",
    x"3D023A23",
    x"3D02074E",
    x"3D01D48D",
    x"3D01A1E0",
    x"3D016F47",
    x"3D013CC1",
    x"3D010A4F",
    x"3D00D7F1",
    x"3D00A5A7",
    x"3D007370",
    x"3D00414D",
    x"3D000F3D",
    x"3CFFBA81",
    x"3CFF56B0",
    x"3CFEF306",
    x"3CFE8F82",
    x"3CFE2C25",
    x"3CFDC8F0",
    x"3CFD65E0",
    x"3CFD02F8",
    x"3CFCA036",
    x"3CFC3D9B",
    x"3CFBDB26",
    x"3CFB78D8",
    x"3CFB16AF",
    x"3CFAB4AE",
    x"3CFA52D2",
    x"3CF9F11D",
    x"3CF98F8E",
    x"3CF92E25",
    x"3CF8CCE2",
    x"3CF86BC5",
    x"3CF80ACE",
    x"3CF7A9FC",
    x"3CF74951",
    x"3CF6E8CB",
    x"3CF6886B",
    x"3CF62830",
    x"3CF5C81C",
    x"3CF5682C",
    x"3CF50862",
    x"3CF4A8BE",
    x"3CF4493E",
    x"3CF3E9E4",
    x"3CF38AB0",
    x"3CF32BA0",
    x"3CF2CCB5",
    x"3CF26DF0",
    x"3CF20F50",
    x"3CF1B0D4",
    x"3CF1527D",
    x"3CF0F44C",
    x"3CF0963E",
    x"3CF03856",
    x"3CEFDA92",
    x"3CEF7CF3",
    x"3CEF1F79",
    x"3CEEC223",
    x"3CEE64F1",
    x"3CEE07E4",
    x"3CEDAAFB",
    x"3CED4E36",
    x"3CECF196",
    x"3CEC951A",
    x"3CEC38C1",
    x"3CEBDC8D",
    x"3CEB807D",
    x"3CEB2491",
    x"3CEAC8C8",
    x"3CEA6D24",
    x"3CEA11A3",
    x"3CE9B646",
    x"3CE95B0D",
    x"3CE8FFF7",
    x"3CE8A505",
    x"3CE84A36",
    x"3CE7EF8B",
    x"3CE79503",
    x"3CE73A9E",
    x"3CE6E05D",
    x"3CE6863F",
    x"3CE62C44",
    x"3CE5D26C",
    x"3CE578B8",
    x"3CE51F26",
    x"3CE4C5B7",
    x"3CE46C6C",
    x"3CE41343",
    x"3CE3BA3C",
    x"3CE36159",
    x"3CE30898",
    x"3CE2AFFA",
    x"3CE2577F",
    x"3CE1FF26",
    x"3CE1A6F0",
    x"3CE14EDC",
    x"3CE0F6EA",
    x"3CE09F1B",
    x"3CE0476E",
    x"3CDFEFE3",
    x"3CDF987A",
    x"3CDF4134",
    x"3CDEEA0F",
    x"3CDE930D",
    x"3CDE3C2C",
    x"3CDDE56E",
    x"3CDD8ED1",
    x"3CDD3856",
    x"3CDCE1FD",
    x"3CDC8BC6",
    x"3CDC35B0",
    x"3CDBDFBC",
    x"3CDB89E9",
    x"3CDB3438",
    x"3CDADEA8",
    x"3CDA893A",
    x"3CDA33ED",
    x"3CD9DEC1",
    x"3CD989B7",
    x"3CD934CE",
    x"3CD8E006",
    x"3CD88B5F",
    x"3CD836D9",
    x"3CD7E274",
    x"3CD78E30",
    x"3CD73A0D",
    x"3CD6E60A",
    x"3CD69229",
    x"3CD63E68",
    x"3CD5EAC8",
    x"3CD59749",
    x"3CD543EA",
    x"3CD4F0AC",
    x"3CD49D8E",
    x"3CD44A91",
    x"3CD3F7B4",
    x"3CD3A4F7",
    x"3CD3525B",
    x"3CD2FFDF",
    x"3CD2AD83",
    x"3CD25B47",
    x"3CD2092C",
    x"3CD1B730",
    x"3CD16554",
    x"3CD11399",
    x"3CD0C1FD",
    x"3CD07081",
    x"3CD01F25",
    x"3CCFCDE9",
    x"3CCF7CCC",
    x"3CCF2BCF",
    x"3CCEDAF2",
    x"3CCE8A34",
    x"3CCE3996",
    x"3CCDE917",
    x"3CCD98B8",
    x"3CCD4878",
    x"3CCCF857",
    x"3CCCA856",
    x"3CCC5874",
    x"3CCC08B1",
    x"3CCBB90D",
    x"3CCB6988",
    x"3CCB1A23",
    x"3CCACADC",
    x"3CCA7BB4",
    x"3CCA2CAB",
    x"3CC9DDC1",
    x"3CC98EF6",
    x"3CC94049",
    x"3CC8F1BC",
    x"3CC8A34D",
    x"3CC854FC",
    x"3CC806CA",
    x"3CC7B8B7",
    x"3CC76AC2",
    x"3CC71CEB",
    x"3CC6CF33",
    x"3CC68199",
    x"3CC6341E",
    x"3CC5E6C1",
    x"3CC59982",
    x"3CC54C61",
    x"3CC4FF5E",
    x"3CC4B279",
    x"3CC465B3",
    x"3CC4190A",
    x"3CC3CC7F",
    x"3CC38012",
    x"3CC333C3",
    x"3CC2E792",
    x"3CC29B7E",
    x"3CC24F88",
    x"3CC203B0",
    x"3CC1B7F5",
    x"3CC16C58",
    x"3CC120D9",
    x"3CC0D576",
    x"3CC08A32",
    x"3CC03F0A",
    x"3CBFF400",
    x"3CBFA914",
    x"3CBF5E44",
    x"3CBF1392",
    x"3CBEC8FD",
    x"3CBE7E85",
    x"3CBE342A",
    x"3CBDE9EC",
    x"3CBD9FCB",
    x"3CBD55C7",
    x"3CBD0BE0",
    x"3CBCC216",
    x"3CBC7869",
    x"3CBC2ED8",
    x"3CBBE564",
    x"3CBB9C0D",
    x"3CBB52D2",
    x"3CBB09B4",
    x"3CBAC0B3",
    x"3CBA77CE",
    x"3CBA2F05",
    x"3CB9E659",
    x"3CB99DC9",
    x"3CB95556",
    x"3CB90CFE",
    x"3CB8C4C3",
    x"3CB87CA5",
    x"3CB834A2",
    x"3CB7ECBB",
    x"3CB7A4F1",
    x"3CB75D43",
    x"3CB715B0",
    x"3CB6CE3A",
    x"3CB686DF",
    x"3CB63FA0",
    x"3CB5F87D",
    x"3CB5B176",
    x"3CB56A8B",
    x"3CB523BB",
    x"3CB4DD07",
    x"3CB4966E",
    x"3CB44FF1",
    x"3CB40990",
    x"3CB3C34A",
    x"3CB37D1F",
    x"3CB33710",
    x"3CB2F11C",
    x"3CB2AB44",
    x"3CB26586",
    x"3CB21FE4",
    x"3CB1DA5D",
    x"3CB194F2",
    x"3CB14FA1",
    x"3CB10A6B",
    x"3CB0C551",
    x"3CB08051",
    x"3CB03B6D",
    x"3CAFF6A3",
    x"3CAFB1F4",
    x"3CAF6D60",
    x"3CAF28E6",
    x"3CAEE488",
    x"3CAEA044",
    x"3CAE5C1B",
    x"3CAE180C",
    x"3CADD418",
    x"3CAD903E",
    x"3CAD4C7F",
    x"3CAD08DA",
    x"3CACC550",
    x"3CAC81E0",
    x"3CAC3E8B",
    x"3CABFB4F",
    x"3CABB82E",
    x"3CAB7527",
    x"3CAB323B",
    x"3CAAEF68",
    x"3CAAACB0",
    x"3CAA6A11",
    x"3CAA278D",
    x"3CA9E522",
    x"3CA9A2D2",
    x"3CA9609B",
    x"3CA91E7E",
    x"3CA8DC7B",
    x"3CA89A92",
    x"3CA858C3",
    x"3CA8170D",
    x"3CA7D571",
    x"3CA793EE",
    x"3CA75285",
    x"3CA71135",
    x"3CA6CFFF",
    x"3CA68EE3",
    x"3CA64DE0",
    x"3CA60CF6",
    x"3CA5CC26",
    x"3CA58B6F",
    x"3CA54AD1",
    x"3CA50A4C",
    x"3CA4C9E1",
    x"3CA4898E",
    x"3CA44955",
    x"3CA40935",
    x"3CA3C92E",
    x"3CA38940",
    x"3CA3496B",
    x"3CA309AF",
    x"3CA2CA0B",
    x"3CA28A81",
    x"3CA24B0F",
    x"3CA20BB6",
    x"3CA1CC76",
    x"3CA18D4E",
    x"3CA14E3F",
    x"3CA10F49",
    x"3CA0D06B",
    x"3CA091A6",
    x"3CA052FA",
    x"3CA01465",
    x"3C9FD5EA",
    x"3C9F9786",
    x"3C9F593B",
    x"3C9F1B09",
    x"3C9EDCEE",
    x"3C9E9EEC",
    x"3C9E6102",
    x"3C9E2330",
    x"3C9DE576",
    x"3C9DA7D5",
    x"3C9D6A4B",
    x"3C9D2CDA",
    x"3C9CEF80",
    x"3C9CB23F",
    x"3C9C7515",
    x"3C9C3803",
    x"3C9BFB09",
    x"3C9BBE27",
    x"3C9B815D",
    x"3C9B44AA",
    x"3C9B080F",
    x"3C9ACB8C",
    x"3C9A8F20",
    x"3C9A52CC",
    x"3C9A168F",
    x"3C99DA6A",
    x"3C999E5D",
    x"3C996267",
    x"3C992688",
    x"3C98EAC0",
    x"3C98AF10",
    x"3C987378",
    x"3C9837F6",
    x"3C97FC8C",
    x"3C97C139",
    x"3C9785FD",
    x"3C974AD8",
    x"3C970FCA",
    x"3C96D4D4",
    x"3C9699F4",
    x"3C965F2C",
    x"3C96247A",
    x"3C95E9DF",
    x"3C95AF5B",
    x"3C9574EE",
    x"3C953A98",
    x"3C950058",
    x"3C94C62F",
    x"3C948C1D",
    x"3C945222",
    x"3C94183D",
    x"3C93DE6F",
    x"3C93A4B7",
    x"3C936B16",
    x"3C93318C",
    x"3C92F818",
    x"3C92BEBA",
    x"3C928573",
    x"3C924C42",
    x"3C921327",
    x"3C91DA23",
    x"3C91A135",
    x"3C91685D",
    x"3C912F9B",
    x"3C90F6EF",
    x"3C90BE5A",
    x"3C9085DB",
    x"3C904D72",
    x"3C90151E",
    x"3C8FDCE1",
    x"3C8FA4BA",
    x"3C8F6CA8",
    x"3C8F34AD",
    x"3C8EFCC7",
    x"3C8EC4F7",
    x"3C8E8D3D",
    x"3C8E5599",
    x"3C8E1E0A",
    x"3C8DE691",
    x"3C8DAF2E",
    x"3C8D77E1",
    x"3C8D40A9",
    x"3C8D0986",
    x"3C8CD279",
    x"3C8C9B82",
    x"3C8C64A0",
    x"3C8C2DD3",
    x"3C8BF71C",
    x"3C8BC07A",
    x"3C8B89ED",
    x"3C8B5376",
    x"3C8B1D14",
    x"3C8AE6C7",
    x"3C8AB090",
    x"3C8A7A6D",
    x"3C8A4460",
    x"3C8A0E68",
    x"3C89D885",
    x"3C89A2B7",
    x"3C896CFE",
    x"3C89375A",
    x"3C8901CB",
    x"3C88CC50",
    x"3C8896EB",
    x"3C88619A",
    x"3C882C5F",
    x"3C87F738",
    x"3C87C226",
    x"3C878D28",
    x"3C87583F",
    x"3C87236B",
    x"3C86EEAC",
    x"3C86BA01",
    x"3C86856A",
    x"3C8650E8",
    x"3C861C7B",
    x"3C85E822",
    x"3C85B3DE",
    x"3C857FAE",
    x"3C854B92",
    x"3C85178B",
    x"3C84E397",
    x"3C84AFB9",
    x"3C847BEE",
    x"3C844838",
    x"3C841496",
    x"3C83E108",
    x"3C83AD8E",
    x"3C837A28",
    x"3C8346D7",
    x"3C831399",
    x"3C82E06F",
    x"3C82AD59",
    x"3C827A58",
    x"3C82476A",
    x"3C821490",
    x"3C81E1CA",
    x"3C81AF18",
    x"3C817C79",
    x"3C8149EE",
    x"3C811777",
    x"3C80E514",
    x"3C80B2C4",
    x"3C808088",
    x"3C804E60",
    x"3C801C4B",
    x"3C7FD493",
    x"3C7F70B8",
    x"3C7F0D03",
    x"3C7EA976",
    x"3C7E460F",
    x"3C7DE2CF",
    x"3C7D7FB6",
    x"3C7D1CC3",
    x"3C7CB9F7",
    x"3C7C5752",
    x"3C7BF4D3",
    x"3C7B927B",
    x"3C7B3049",
    x"3C7ACE3D",
    x"3C7A6C57",
    x"3C7A0A98",
    x"3C79A8FF",
    x"3C79478C",
    x"3C78E63F",
    x"3C788518",
    x"3C782417",
    x"3C77C33C",
    x"3C776287",
    x"3C7701F7",
    x"3C76A18D",
    x"3C764149",
    x"3C75E12A",
    x"3C758131",
    x"3C75215D",
    x"3C74C1AF",
    x"3C746226",
    x"3C7402C2",
    x"3C73A384",
    x"3C73446A",
    x"3C72E576",
    x"3C7286A7",
    x"3C7227FD",
    x"3C71C978",
    x"3C716B18",
    x"3C710CDC",
    x"3C70AEC6",
    x"3C7050D4",
    x"3C6FF306",
    x"3C6F955E",
    x"3C6F37DA",
    x"3C6EDA7A",
    x"3C6E7D3F",
    x"3C6E2028",
    x"3C6DC336",
    x"3C6D6668",
    x"3C6D09BE",
    x"3C6CAD38",
    x"3C6C50D6",
    x"3C6BF499",
    x"3C6B987F",
    x"3C6B3C8A",
    x"3C6AE0B8",
    x"3C6A850A",
    x"3C6A2980",
    x"3C69CE1A",
    x"3C6972D7",
    x"3C6917B8",
    x"3C68BCBC",
    x"3C6861E4",
    x"3C680730",
    x"3C67AC9F",
    x"3C675231",
    x"3C66F7E7",
    x"3C669DBF",
    x"3C6643BB",
    x"3C65E9DA",
    x"3C65901D",
    x"3C653682",
    x"3C64DD0A",
    x"3C6483B5",
    x"3C642A83",
    x"3C63D174",
    x"3C637887",
    x"3C631FBE",
    x"3C62C717",
    x"3C626E92",
    x"3C621630",
    x"3C61BDF1",
    x"3C6165D4",
    x"3C610DD9",
    x"3C60B601",
    x"3C605E4B",
    x"3C6006B7",
    x"3C5FAF46",
    x"3C5F57F6",
    x"3C5F00C9",
    x"3C5EA9BE",
    x"3C5E52D4",
    x"3C5DFC0D",
    x"3C5DA567",
    x"3C5D4EE4",
    x"3C5CF882",
    x"3C5CA242",
    x"3C5C4C23",
    x"3C5BF626",
    x"3C5BA04B",
    x"3C5B4A91",
    x"3C5AF4F8",
    x"3C5A9F81",
    x"3C5A4A2C",
    x"3C59F4F8",
    x"3C599FE4",
    x"3C594AF3",
    x"3C58F622",
    x"3C58A172",
    x"3C584CE4",
    x"3C57F876",
    x"3C57A42A",
    x"3C574FFE",
    x"3C56FBF3",
    x"3C56A809",
    x"3C565440",
    x"3C560097",
    x"3C55AD0F",
    x"3C5559A8",
    x"3C550661",
    x"3C54B33B",
    x"3C546035",
    x"3C540D50",
    x"3C53BA8B",
    x"3C5367E6",
    x"3C531562",
    x"3C52C2FD",
    x"3C5270B9",
    x"3C521E95",
    x"3C51CC91",
    x"3C517AAD",
    x"3C5128E9",
    x"3C50D745",
    x"3C5085C1",
    x"3C50345D",
    x"3C4FE318",
    x"3C4F91F4",
    x"3C4F40EE",
    x"3C4EF009",
    x"3C4E9F43",
    x"3C4E4E9C",
    x"3C4DFE15",
    x"3C4DADAE",
    x"3C4D5D66",
    x"3C4D0D3D",
    x"3C4CBD33",
    x"3C4C6D49",
    x"3C4C1D7E",
    x"3C4BCDD2",
    x"3C4B7E45",
    x"3C4B2ED7",
    x"3C4ADF88",
    x"3C4A9059",
    x"3C4A4148",
    x"3C49F256",
    x"3C49A382",
    x"3C4954CE",
    x"3C490638",
    x"3C48B7C1",
    x"3C486969",
    x"3C481B2F",
    x"3C47CD13",
    x"3C477F16",
    x"3C473138",
    x"3C46E378",
    x"3C4695D6",
    x"3C464853",
    x"3C45FAEE",
    x"3C45ADA7",
    x"3C45607E",
    x"3C451373",
    x"3C44C687",
    x"3C4479B8",
    x"3C442D08",
    x"3C43E075",
    x"3C439400",
    x"3C4347A9",
    x"3C42FB70",
    x"3C42AF55",
    x"3C426357",
    x"3C421777",
    x"3C41CBB5",
    x"3C418010",
    x"3C413489",
    x"3C40E91F",
    x"3C409DD3",
    x"3C4052A4",
    x"3C400792",
    x"3C3FBC9E",
    x"3C3F71C7",
    x"3C3F270D",
    x"3C3EDC70",
    x"3C3E91F1",
    x"3C3E478E",
    x"3C3DFD49",
    x"3C3DB320",
    x"3C3D6915",
    x"3C3D1F26",
    x"3C3CD555",
    x"3C3C8BA0",
    x"3C3C4207",
    x"3C3BF88C",
    x"3C3BAF2D",
    x"3C3B65EB",
    x"3C3B1CC6",
    x"3C3AD3BD",
    x"3C3A8AD0",
    x"3C3A4200",
    x"3C39F94D",
    x"3C39B0B5",
    x"3C39683B",
    x"3C391FDC",
    x"3C38D79A",
    x"3C388F73",
    x"3C38476A",
    x"3C37FF7C",
    x"3C37B7AA",
    x"3C376FF4",
    x"3C37285A",
    x"3C36E0DD",
    x"3C36997B",
    x"3C365235",
    x"3C360B0B",
    x"3C35C3FC",
    x"3C357D09",
    x"3C353632",
    x"3C34EF77",
    x"3C34A8D7",
    x"3C346253",
    x"3C341BEA",
    x"3C33D59D",
    x"3C338F6C",
    x"3C334955",
    x"3C33035A",
    x"3C32BD7B",
    x"3C3277B6",
    x"3C32320D",
    x"3C31EC7F",
    x"3C31A70C",
    x"3C3161B5",
    x"3C311C78",
    x"3C30D756",
    x"3C309250",
    x"3C304D64",
    x"3C300893",
    x"3C2FC3DD",
    x"3C2F7F42",
    x"3C2F3AC2",
    x"3C2EF65C",
    x"3C2EB211",
    x"3C2E6DE1",
    x"3C2E29CC",
    x"3C2DE5D0",
    x"3C2DA1F0",
    x"3C2D5E2A",
    x"3C2D1A7E",
    x"3C2CD6ED",
    x"3C2C9376",
    x"3C2C501A",
    x"3C2C0CD8",
    x"3C2BC9B0",
    x"3C2B86A2",
    x"3C2B43AF",
    x"3C2B00D5",
    x"3C2ABE16",
    x"3C2A7B71",
    x"3C2A38E6",
    x"3C29F674",
    x"3C29B41D",
    x"3C2971E0",
    x"3C292FBC",
    x"3C28EDB2",
    x"3C28ABC2",
    x"3C2869EC",
    x"3C282830",
    x"3C27E68D",
    x"3C27A504",
    x"3C276394",
    x"3C27223E",
    x"3C26E101",
    x"3C269FDE",
    x"3C265ED4",
    x"3C261DE4",
    x"3C25DD0D",
    x"3C259C4F",
    x"3C255BAB",
    x"3C251B1F",
    x"3C24DAAD",
    x"3C249A55",
    x"3C245A15",
    x"3C2419EE",
    x"3C23D9E1",
    x"3C2399EC",
    x"3C235A10",
    x"3C231A4E",
    x"3C22DAA4",
    x"3C229B13",
    x"3C225B9B",
    x"3C221C3B",
    x"3C21DCF5",
    x"3C219DC7",
    x"3C215EB1",
    x"3C211FB5",
    x"3C20E0D1",
    x"3C20A205",
    x"3C206352",
    x"3C2024B7",
    x"3C1FE635",
    x"3C1FA7CB",
    x"3C1F697A",
    x"3C1F2B41",
    x"3C1EED20",
    x"3C1EAF18",
    x"3C1E7128",
    x"3C1E334F",
    x"3C1DF58F",
    x"3C1DB7E8",
    x"3C1D7A58",
    x"3C1D3CE0",
    x"3C1CFF80",
    x"3C1CC238",
    x"3C1C8508",
    x"3C1C47F0",
    x"3C1C0AF0",
    x"3C1BCE08",
    x"3C1B9137",
    x"3C1B547E",
    x"3C1B17DD",
    x"3C1ADB54",
    x"3C1A9EE2",
    x"3C1A6288",
    x"3C1A2645",
    x"3C19EA1A",
    x"3C19AE06",
    x"3C19720A",
    x"3C193625",
    x"3C18FA57",
    x"3C18BEA1",
    x"3C188302",
    x"3C18477B",
    x"3C180C0B",
    x"3C17D0B1",
    x"3C179570",
    x"3C175A45",
    x"3C171F31",
    x"3C16E434",
    x"3C16A94F",
    x"3C166E80",
    x"3C1633C8",
    x"3C15F928",
    x"3C15BE9E",
    x"3C15842B",
    x"3C1549CE",
    x"3C150F89",
    x"3C14D55A",
    x"3C149B42",
    x"3C146141",
    x"3C142756",
    x"3C13ED82",
    x"3C13B3C5",
    x"3C137A1E",
    x"3C13408D",
    x"3C130713",
    x"3C12CDB0",
    x"3C129463",
    x"3C125B2C",
    x"3C12220B",
    x"3C11E901",
    x"3C11B00D",
    x"3C117730",
    x"3C113E68",
    x"3C1105B7",
    x"3C10CD1C",
    x"3C109497",
    x"3C105C28",
    x"3C1023CF",
    x"3C0FEB8C",
    x"3C0FB35F",
    x"3C0F7B48",
    x"3C0F4346",
    x"3C0F0B5B",
    x"3C0ED385",
    x"3C0E9BC6",
    x"3C0E641C",
    x"3C0E2C87",
    x"3C0DF509",
    x"3C0DBDA0",
    x"3C0D864D",
    x"3C0D4F0F",
    x"3C0D17E7",
    x"3C0CE0D4",
    x"3C0CA9D7",
    x"3C0C72F0",
    x"3C0C3C1E",
    x"3C0C0561",
    x"3C0BCEB9",
    x"3C0B9827",
    x"3C0B61AA",
    x"3C0B2B43",
    x"3C0AF4F1",
    x"3C0ABEB4",
    x"3C0A888C",
    x"3C0A5279",
    x"3C0A1C7B",
    x"3C09E693",
    x"3C09B0BF",
    x"3C097B00",
    x"3C094557",
    x"3C090FC2",
    x"3C08DA43",
    x"3C08A4D8",
    x"3C086F82",
    x"3C083A41",
    x"3C080514",
    x"3C07CFFD",
    x"3C079AFA",
    x"3C07660C",
    x"3C073132",
    x"3C06FC6D",
    x"3C06C7BD",
    x"3C069321",
    x"3C065E9A",
    x"3C062A27",
    x"3C05F5C9",
    x"3C05C17F",
    x"3C058D4A",
    x"3C055929",
    x"3C05251C",
    x"3C04F124",
    x"3C04BD40",
    x"3C048970",
    x"3C0455B4",
    x"3C04220D",
    x"3C03EE7A",
    x"3C03BAFB",
    x"3C038790",
    x"3C035439",
    x"3C0320F6",
    x"3C02EDC7",
    x"3C02BAAC",
    x"3C0287A5",
    x"3C0254B2",
    x"3C0221D3",
    x"3C01EF08",
    x"3C01BC50",
    x"3C0189AC",
    x"3C01571D",
    x"3C0124A0",
    x"3C00F238",
    x"3C00BFE3",
    x"3C008DA2",
    x"3C005B74",
    x"3C00295B",
    x"3BFFEEA8",
    x"3BFF8AC3",
    x"3BFF2704",
    x"3BFEC36C",
    x"3BFE5FFB",
    x"3BFDFCB1",
    x"3BFD998E",
    x"3BFD3691",
    x"3BFCD3BB",
    x"3BFC710C",
    x"3BFC0E83",
    x"3BFBAC20",
    x"3BFB49E4",
    x"3BFAE7CF",
    x"3BFA85DF",
    x"3BFA2416",
    x"3BF9C273",
    x"3BF960F6",
    x"3BF8FF9F",
    x"3BF89E6E",
    x"3BF83D63",
    x"3BF7DC7E",
    x"3BF77BBF",
    x"3BF71B26",
    x"3BF6BAB2",
    x"3BF65A64",
    x"3BF5FA3B",
    x"3BF59A38",
    x"3BF53A5B",
    x"3BF4DAA3",
    x"3BF47B10",
    x"3BF41BA3",
    x"3BF3BC5A",
    x"3BF35D37",
    x"3BF2FE3A",
    x"3BF29F61",
    x"3BF240AD",
    x"3BF1E21E",
    x"3BF183B4",
    x"3BF1256F",
    x"3BF0C74F",
    x"3BF06954",
    x"3BF00B7D",
    x"3BEFADCB",
    x"3BEF503D",
    x"3BEEF2D4",
    x"3BEE958F",
    x"3BEE386F",
    x"3BEDDB73",
    x"3BED7E9C",
    x"3BED21E8",
    x"3BECC559",
    x"3BEC68EE",
    x"3BEC0CA7",
    x"3BEBB084",
    x"3BEB5485",
    x"3BEAF8AA",
    x"3BEA9CF3",
    x"3BEA415F",
    x"3BE9E5F0",
    x"3BE98AA4",
    x"3BE92F7B",
    x"3BE8D477",
    x"3BE87995",
    x"3BE81ED8",
    x"3BE7C43D",
    x"3BE769C6",
    x"3BE70F73",
    x"3BE6B542",
    x"3BE65B35",
    x"3BE6014B",
    x"3BE5A784",
    x"3BE54DE0",
    x"3BE4F45F",
    x"3BE49B01",
    x"3BE441C6",
    x"3BE3E8AE",
    x"3BE38FB8",
    x"3BE336E5",
    x"3BE2DE35",
    x"3BE285A8",
    x"3BE22D3D",
    x"3BE1D4F4",
    x"3BE17CCE",
    x"3BE124CB",
    x"3BE0CCEA",
    x"3BE0752B",
    x"3BE01D8E",
    x"3BDFC614",
    x"3BDF6EBB",
    x"3BDF1785",
    x"3BDEC071",
    x"3BDE697F",
    x"3BDE12AF",
    x"3BDDBC00",
    x"3BDD6574",
    x"3BDD0F09",
    x"3BDCB8C0",
    x"3BDC6299",
    x"3BDC0C93",
    x"3BDBB6AF",
    x"3BDB60EC",
    x"3BDB0B4B",
    x"3BDAB5CB",
    x"3BDA606D",
    x"3BDA0B30",
    x"3BD9B614",
    x"3BD9611A",
    x"3BD90C40",
    x"3BD8B788",
    x"3BD862F1",
    x"3BD80E7B",
    x"3BD7BA26",
    x"3BD765F1",
    x"3BD711DE",
    x"3BD6BDEB",
    x"3BD66A1A",
    x"3BD61668",
    x"3BD5C2D8",
    x"3BD56F68",
    x"3BD51C19",
    x"3BD4C8EA",
    x"3BD475DC",
    x"3BD422EE",
    x"3BD3D021",
    x"3BD37D74",
    x"3BD32AE7",
    x"3BD2D87A",
    x"3BD2862D",
    x"3BD23401",
    x"3BD1E1F5",
    x"3BD19009",
    x"3BD13E3C",
    x"3BD0EC90",
    x"3BD09B03",
    x"3BD04997",
    x"3BCFF84A",
    x"3BCFA71D",
    x"3BCF560F",
    x"3BCF0522",
    x"3BCEB453",
    x"3BCE63A5",
    x"3BCE1316",
    x"3BCDC2A6",
    x"3BCD7255",
    x"3BCD2224",
    x"3BCCD213",
    x"3BCC8220",
    x"3BCC324D",
    x"3BCBE299",
    x"3BCB9304",
    x"3BCB438E",
    x"3BCAF437",
    x"3BCAA4FF",
    x"3BCA55E6",
    x"3BCA06EC",
    x"3BC9B811",
    x"3BC96954",
    x"3BC91AB7",
    x"3BC8CC37",
    x"3BC87DD7",
    x"3BC82F95",
    x"3BC7E172",
    x"3BC7936D",
    x"3BC74587",
    x"3BC6F7BF",
    x"3BC6AA15",
    x"3BC65C8A",
    x"3BC60F1D",
    x"3BC5C1CE",
    x"3BC5749D",
    x"3BC5278B",
    x"3BC4DA96",
    x"3BC48DC0",
    x"3BC44108",
    x"3BC3F46D",
    x"3BC3A7F1",
    x"3BC35B92",
    x"3BC30F51",
    x"3BC2C32E",
    x"3BC27729",
    x"3BC22B41",
    x"3BC1DF77",
    x"3BC193CA",
    x"3BC1483B",
    x"3BC0FCCA",
    x"3BC0B176",
    x"3BC0663F",
    x"3BC01B26",
    x"3BBFD02A",
    x"3BBF854B",
    x"3BBF3A8A",
    x"3BBEEFE6",
    x"3BBEA55E",
    x"3BBE5AF4",
    x"3BBE10A7",
    x"3BBDC677",
    x"3BBD7C64",
    x"3BBD326E",
    x"3BBCE895",
    x"3BBC9ED8",
    x"3BBC5539",
    x"3BBC0BB6",
    x"3BBBC250",
    x"3BBB7906",
    x"3BBB2FD9",
    x"3BBAE6C9",
    x"3BBA9DD5",
    x"3BBA54FD",
    x"3BBA0C42",
    x"3BB9C3A4",
    x"3BB97B21",
    x"3BB932BB",
    x"3BB8EA72",
    x"3BB8A244",
    x"3BB85A33",
    x"3BB8123E",
    x"3BB7CA65",
    x"3BB782A8",
    x"3BB73B07",
    x"3BB6F382",
    x"3BB6AC18",
    x"3BB664CB",
    x"3BB61D9A",
    x"3BB5D684",
    x"3BB58F8A",
    x"3BB548AC",
    x"3BB501E9",
    x"3BB4BB42",
    x"3BB474B7",
    x"3BB42E47",
    x"3BB3E7F3",
    x"3BB3A1BA",
    x"3BB35B9C",
    x"3BB3159A",
    x"3BB2CFB4",
    x"3BB289E8",
    x"3BB24438",
    x"3BB1FEA3",
    x"3BB1B929",
    x"3BB173CA",
    x"3BB12E86",
    x"3BB0E95E",
    x"3BB0A450",
    x"3BB05F5D",
    x"3BB01A85",
    x"3BAFD5C9",
    x"3BAF9126",
    x"3BAF4C9F",
    x"3BAF0833",
    x"3BAEC3E1",
    x"3BAE7FAA",
    x"3BAE3B8D",
    x"3BADF78B",
    x"3BADB3A4",
    x"3BAD6FD7",
    x"3BAD2C24",
    x"3BACE88C",
    x"3BACA50E",
    x"3BAC61AB",
    x"3BAC1E62",
    x"3BABDB33",
    x"3BAB981F",
    x"3BAB5525",
    x"3BAB1244",
    x"3BAACF7E",
    x"3BAA8CD2",
    x"3BAA4A40",
    x"3BAA07C8",
    x"3BA9C56A",
    x"3BA98326",
    x"3BA940FC",
    x"3BA8FEEB",
    x"3BA8BCF5",
    x"3BA87B18",
    x"3BA83954",
    x"3BA7F7AB",
    x"3BA7B61B",
    x"3BA774A4",
    x"3BA73348",
    x"3BA6F204",
    x"3BA6B0DB",
    x"3BA66FCA",
    x"3BA62ED3",
    x"3BA5EDF6",
    x"3BA5AD31",
    x"3BA56C86",
    x"3BA52BF5",
    x"3BA4EB7C",
    x"3BA4AB1D",
    x"3BA46AD6",
    x"3BA42AA9",
    x"3BA3EA95",
    x"3BA3AA9A",
    x"3BA36AB8",
    x"3BA32AEE",
    x"3BA2EB3E",
    x"3BA2ABA7",
    x"3BA26C28",
    x"3BA22CC2",
    x"3BA1ED75",
    x"3BA1AE41",
    x"3BA16F25",
    x"3BA13022",
    x"3BA0F137",
    x"3BA0B265",
    x"3BA073AC",
    x"3BA0350B",
    x"3B9FF682",
    x"3B9FB812",
    x"3B9F79BB",
    x"3B9F3B7B",
    x"3B9EFD54",
    x"3B9EBF45",
    x"3B9E814F",
    x"3B9E4370",
    x"3B9E05AA",
    x"3B9DC7FC",
    x"3B9D8A66",
    x"3B9D4CE8",
    x"3B9D0F82",
    x"3B9CD234",
    x"3B9C94FD",
    x"3B9C57DF",
    x"3B9C1AD9",
    x"3B9BDDEA",
    x"3B9BA113",
    x"3B9B6454",
    x"3B9B27AD",
    x"3B9AEB1D",
    x"3B9AAEA5",
    x"3B9A7245",
    x"3B9A35FC",
    x"3B99F9CB",
    x"3B99BDB1",
    x"3B9981AE",
    x"3B9945C3",
    x"3B9909F0",
    x"3B98CE34",
    x"3B98928F",
    x"3B985701",
    x"3B981B8B",
    x"3B97E02C",
    x"3B97A4E4",
    x"3B9769B3",
    x"3B972E99",
    x"3B96F396",
    x"3B96B8AB",
    x"3B967DD6",
    x"3B964318",
    x"3B960872",
    x"3B95CDE2",
    x"3B959369",
    x"3B955907",
    x"3B951EBB",
    x"3B94E487",
    x"3B94AA69",
    x"3B947062",
    x"3B943671",
    x"3B93FC97",
    x"3B93C2D4",
    x"3B938927",
    x"3B934F90",
    x"3B931611",
    x"3B92DCA7",
    x"3B92A354",
    x"3B926A18",
    x"3B9230F1",
    x"3B91F7E1",
    x"3B91BEE8",
    x"3B918604",
    x"3B914D37",
    x"3B911480",
    x"3B90DBDF",
    x"3B90A354",
    x"3B906ADF",
    x"3B903281",
    x"3B8FFA38",
    x"3B8FC205",
    x"3B8F89E8",
    x"3B8F51E1",
    x"3B8F19F0",
    x"3B8EE215",
    x"3B8EAA50",
    x"3B8E72A0",
    x"3B8E3B06",
    x"3B8E0382",
    x"3B8DCC13",
    x"3B8D94BA",
    x"3B8D5D77",
    x"3B8D2649",
    x"3B8CEF31",
    x"3B8CB82E",
    x"3B8C8141",
    x"3B8C4A69",
    x"3B8C13A7",
    x"3B8BDCFA",
    x"3B8BA662",
    x"3B8B6FE0",
    x"3B8B3973",
    x"3B8B031B",
    x"3B8ACCD9",
    x"3B8A96AB",
    x"3B8A6093",
    x"3B8A2A90",
    x"3B89F4A2",
    x"3B89BEC9",
    x"3B898905",
    x"3B895356",
    x"3B891DBB",
    x"3B88E836",
    x"3B88B2C6",
    x"3B887D6B",
    x"3B884824",
    x"3B8812F2",
    x"3B87DDD5",
    x"3B87A8CD",
    x"3B8773D9",
    x"3B873EFA",
    x"3B870A30",
    x"3B86D57A",
    x"3B86A0D9",
    x"3B866C4D",
    x"3B8637D5",
    x"3B860371",
    x"3B85CF22",
    x"3B859AE7",
    x"3B8566C1",
    x"3B8532AF",
    x"3B84FEB1",
    x"3B84CAC8",
    x"3B8496F3",
    x"3B846332",
    x"3B842F85",
    x"3B83FBED",
    x"3B83C869",
    x"3B8394F8",
    x"3B83619C",
    x"3B832E54",
    x"3B82FB20",
    x"3B82C800",
    x"3B8294F4",
    x"3B8261FC",
    x"3B822F17",
    x"3B81FC47",
    x"3B81C98A",
    x"3B8196E1",
    x"3B81644C",
    x"3B8131CB",
    x"3B80FF5D",
    x"3B80CD03",
    x"3B809ABD",
    x"3B80688A",
    x"3B80366B",
    x"3B800460",
    x"3B7FA4D0",
    x"3B7F4107",
    x"3B7EDD65",
    x"3B7E79EA",
    x"3B7E1696",
    x"3B7DB368",
    x"3B7D5062",
    x"3B7CED82",
    x"3B7C8AC8",
    x"3B7C2835",
    x"3B7BC5C9",
    x"3B7B6383",
    x"3B7B0163",
    x"3B7A9F6A",
    x"3B7A3D96",
    x"3B79DBE9",
    x"3B797A63",
    x"3B791902",
    x"3B78B7C7",
    x"3B7856B2",
    x"3B77F5C3",
    x"3B7794FA",
    x"3B773457",
    x"3B76D3D9",
    x"3B767381",
    x"3B76134F",
    x"3B75B342",
    x"3B75535B",
    x"3B74F399",
    x"3B7493FD",
    x"3B743485",
    x"3B73D534",
    x"3B737607",
    x"3B7316FF",
    x"3B72B81D",
    x"3B72595F",
    x"3B71FAC7",
    x"3B719C54",
    x"3B713E05",
    x"3B70DFDB",
    x"3B7081D6",
    x"3B7023F6",
    x"3B6FC63A",
    x"3B6F68A3",
    x"3B6F0B30",
    x"3B6EADE2",
    x"3B6E50B8",
    x"3B6DF3B3",
    x"3B6D96D2",
    x"3B6D3A15",
    x"3B6CDD7C",
    x"3B6C8108",
    x"3B6C24B8",
    x"3B6BC88B",
    x"3B6B6C83",
    x"3B6B109E",
    x"3B6AB4DE",
    x"3B6A5941",
    x"3B69FDC8",
    x"3B69A273",
    x"3B694741",
    x"3B68EC33",
    x"3B689149",
    x"3B683682",
    x"3B67DBDE",
    x"3B67815E",
    x"3B672701",
    x"3B66CCC7",
    x"3B6672B1",
    x"3B6618BE",
    x"3B65BEEE",
    x"3B656541",
    x"3B650BB7",
    x"3B64B24F",
    x"3B64590B",
    x"3B63FFEA",
    x"3B63A6EB",
    x"3B634E0F",
    x"3B62F556",
    x"3B629CC0",
    x"3B62444C",
    x"3B61EBFA",
    x"3B6193CB",
    x"3B613BBF",
    x"3B60E3D5",
    x"3B608C0D",
    x"3B603467",
    x"3B5FDCE4",
    x"3B5F8583",
    x"3B5F2E44",
    x"3B5ED727",
    x"3B5E802B",
    x"3B5E2952",
    x"3B5DD29B",
    x"3B5D7C06",
    x"3B5D2592",
    x"3B5CCF40",
    x"3B5C7910",
    x"3B5C2302",
    x"3B5BCD15",
    x"3B5B774A",
    x"3B5B21A0",
    x"3B5ACC17",
    x"3B5A76B0",
    x"3B5A216B",
    x"3B59CC46",
    x"3B597743",
    x"3B592261",
    x"3B58CDA0",
    x"3B587900",
    x"3B582482",
    x"3B57D024",
    x"3B577BE7",
    x"3B5727CB",
    x"3B56D3D0",
    x"3B567FF5",
    x"3B562C3C",
    x"3B55D8A3",
    x"3B55852B",
    x"3B5531D3",
    x"3B54DE9C",
    x"3B548B85",
    x"3B54388F",
    x"3B53E5B9",
    x"3B539303",
    x"3B53406E",
    x"3B52EDF9",
    x"3B529BA4",
    x"3B52496F",
    x"3B51F75B",
    x"3B51A566",
    x"3B515391",
    x"3B5101DD",
    x"3B50B048",
    x"3B505ED3",
    x"3B500D7E",
    x"3B4FBC48",
    x"3B4F6B33",
    x"3B4F1A3D",
    x"3B4EC966",
    x"3B4E78AF",
    x"3B4E2818",
    x"3B4DD7A0",
    x"3B4D8747",
    x"3B4D370E",
    x"3B4CE6F4",
    x"3B4C96FA",
    x"3B4C471E",
    x"3B4BF762",
    x"3B4BA7C5",
    x"3B4B5847",
    x"3B4B08E8",
    x"3B4AB9A8",
    x"3B4A6A87",
    x"3B4A1B85",
    x"3B49CCA2",
    x"3B497DDD",
    x"3B492F37",
    x"3B48E0B0",
    x"3B489248",
    x"3B4843FE",
    x"3B47F5D2",
    x"3B47A7C6",
    x"3B4759D7",
    x"3B470C07",
    x"3B46BE56",
    x"3B4670C3",
    x"3B46234E",
    x"3B45D5F7",
    x"3B4588BF",
    x"3B453BA4",
    x"3B44EEA8",
    x"3B44A1CA",
    x"3B44550A",
    x"3B440867",
    x"3B43BBE3",
    x"3B436F7D",
    x"3B432334",
    x"3B42D709",
    x"3B428AFC",
    x"3B423F0D",
    x"3B41F33B",
    x"3B41A786",
    x"3B415BF0",
    x"3B411077",
    x"3B40C51B",
    x"3B4079DD",
    x"3B402EBC",
    x"3B3FE3B8",
    x"3B3F98D2",
    x"3B3F4E09",
    x"3B3F035D",
    x"3B3EB8CE",
    x"3B3E6E5C",
    x"3B3E2408",
    x"3B3DD9D0",
    x"3B3D8FB6",
    x"3B3D45B8",
    x"3B3CFBD7",
    x"3B3CB213",
    x"3B3C686C",
    x"3B3C1EE2",
    x"3B3BD574",
    x"3B3B8C23",
    x"3B3B42EE",
    x"3B3AF9D7",
    x"3B3AB0DB",
    x"3B3A67FC",
    x"3B3A1F3A",
    x"3B39D694",
    x"3B398E0A",
    x"3B39459D",
    x"3B38FD4C",
    x"3B38B517",
    x"3B386CFE",
    x"3B382502",
    x"3B37DD21",
    x"3B37955D",
    x"3B374DB5",
    x"3B370628",
    x"3B36BEB8",
    x"3B367763",
    x"3B36302B",
    x"3B35E90E",
    x"3B35A20D",
    x"3B355B27",
    x"3B35145D",
    x"3B34CDAF",
    x"3B34871D",
    x"3B3440A6",
    x"3B33FA4A",
    x"3B33B40A",
    x"3B336DE5",
    x"3B3327DC",
    x"3B32E1EE",
    x"3B329C1C",
    x"3B325664",
    x"3B3210C8",
    x"3B31CB47",
    x"3B3185E1",
    x"3B314097",
    x"3B30FB67",
    x"3B30B652",
    x"3B307158",
    x"3B302C7A",
    x"3B2FE7B6",
    x"3B2FA30D",
    x"3B2F5E7E",
    x"3B2F1A0B",
    x"3B2ED5B2",
    x"3B2E9174",
    x"3B2E4D50",
    x"3B2E0947",
    x"3B2DC559",
    x"3B2D8185",
    x"3B2D3DCC",
    x"3B2CFA2D",
    x"3B2CB6A8",
    x"3B2C733E",
    x"3B2C2FEE",
    x"3B2BECB9",
    x"3B2BA99D",
    x"3B2B669C",
    x"3B2B23B5",
    x"3B2AE0E8",
    x"3B2A9E35",
    x"3B2A5B9D",
    x"3B2A191E",
    x"3B29D6B9",
    x"3B29946E",
    x"3B29523D",
    x"3B291026",
    x"3B28CE28",
    x"3B288C45",
    x"3B284A7B",
    x"3B2808CB",
    x"3B27C734",
    x"3B2785B7",
    x"3B274453",
    x"3B270309",
    x"3B26C1D9",
    x"3B2680C2",
    x"3B263FC4",
    x"3B25FEE0",
    x"3B25BE15",
    x"3B257D64",
    x"3B253CCB",
    x"3B24FC4C",
    x"3B24BBE6",
    x"3B247B99",
    x"3B243B66",
    x"3B23FB4B",
    x"3B23BB49",
    x"3B237B61",
    x"3B233B91",
    x"3B22FBDA",
    x"3B22BC3C",
    x"3B227CB7",
    x"3B223D4B",
    x"3B21FDF7",
    x"3B21BEBC",
    x"3B217F9A",
    x"3B214091",
    x"3B2101A0",
    x"3B20C2C7",
    x"3B208407",
    x"3B204560",
    x"3B2006D1",
    x"3B1FC85B",
    x"3B1F89FD",
    x"3B1F4BB7",
    x"3B1F0D8A",
    x"3B1ECF74",
    x"3B1E9177",
    x"3B1E5393",
    x"3B1E15C6",
    x"3B1DD812",
    x"3B1D9A75",
    x"3B1D5CF1",
    x"3B1D1F85",
    x"3B1CE230",
    x"3B1CA4F4",
    x"3B1C67CF",
    x"3B1C2AC3",
    x"3B1BEDCE",
    x"3B1BB0F1",
    x"3B1B742C",
    x"3B1B377E",
    x"3B1AFAE8",
    x"3B1ABE6A",
    x"3B1A8204",
    x"3B1A45B5",
    x"3B1A097D",
    x"3B19CD5D",
    x"3B199155",
    x"3B195564",
    x"3B19198A",
    x"3B18DDC8",
    x"3B18A21D",
    x"3B186689",
    x"3B182B0D",
    x"3B17EFA7",
    x"3B17B459",
    x"3B177923",
    x"3B173E03",
    x"3B1702FA",
    x"3B16C808",
    x"3B168D2E",
    x"3B16526A",
    x"3B1617BD",
    x"3B15DD28",
    x"3B15A2A9",
    x"3B156840",
    x"3B152DEF",
    x"3B14F3B5",
    x"3B14B991",
    x"3B147F84",
    x"3B14458D",
    x"3B140BAD",
    x"3B13D1E4",
    x"3B139831",
    x"3B135E95",
    x"3B13250F",
    x"3B12EBA0",
    x"3B12B247",
    x"3B127905",
    x"3B123FD9",
    x"3B1206C3",
    x"3B11CDC3",
    x"3B1194DA",
    x"3B115C07",
    x"3B11234A",
    x"3B10EAA4",
    x"3B10B213",
    x"3B107998",
    x"3B104134",
    x"3B1008E5",
    x"3B0FD0AD",
    x"3B0F988A",
    x"3B0F607E",
    x"3B0F2887",
    x"3B0EF0A6",
    x"3B0EB8DB",
    x"3B0E8126",
    x"3B0E4986",
    x"3B0E11FC",
    x"3B0DDA88",
    x"3B0DA329",
    x"3B0D6BE1",
    x"3B0D34AD",
    x"3B0CFD8F",
    x"3B0CC687",
    x"3B0C8F94",
    x"3B0C58B7",
    x"3B0C21EF",
    x"3B0BEB3C",
    x"3B0BB49F",
    x"3B0B7E17",
    x"3B0B47A5",
    x"3B0B1147",
    x"3B0ADAFF",
    x"3B0AA4CC",
    x"3B0A6EAE",
    x"3B0A38A6",
    x"3B0A02B2",
    x"3B09CCD4",
    x"3B09970A",
    x"3B096156",
    x"3B092BB6",
    x"3B08F62B",
    x"3B08C0B6",
    x"3B088B55",
    x"3B085609",
    x"3B0820D2",
    x"3B07EBAF",
    x"3B07B6A1",
    x"3B0781A8",
    x"3B074CC4",
    x"3B0717F4",
    x"3B06E339",
    x"3B06AE93",
    x"3B067A01",
    x"3B064584",
    x"3B06111B",
    x"3B05DCC6",
    x"3B05A886",
    x"3B05745B",
    x"3B054043",
    x"3B050C40",
    x"3B04D852",
    x"3B04A477",
    x"3B0470B1",
    x"3B043CFF",
    x"3B040962",
    x"3B03D5D8",
    x"3B03A262",
    x"3B036F01",
    x"3B033BB4",
    x"3B03087A",
    x"3B02D555",
    x"3B02A244",
    x"3B026F46",
    x"3B023C5D",
    x"3B020987",
    x"3B01D6C5",
    x"3B01A417",
    x"3B01717D",
    x"3B013EF7",
    x"3B010C84",
    x"3B00DA25",
    x"3B00A7DA",
    x"3B0075A2",
    x"3B00437E",
    x"3B00116D",
    x"3AFFBEE0",
    x"3AFF5B0D",
    x"3AFEF761",
    x"3AFE93DC",
    x"3AFE307D",
    x"3AFDCD46",
    x"3AFD6A35",
    x"3AFD074B",
    x"3AFCA487",
    x"3AFC41EA",
    x"3AFBDF74",
    x"3AFB7D24",
    x"3AFB1AFA",
    x"3AFAB8F7",
    x"3AFA5719",
    x"3AF9F562",
    x"3AF993D2",
    x"3AF93267",
    x"3AF8D122",
    x"3AF87004",
    x"3AF80F0B",
    x"3AF7AE38",
    x"3AF74D8B",
    x"3AF6ED03",
    x"3AF68CA1",
    x"3AF62C65",
    x"3AF5CC4F",
    x"3AF56C5E",
    x"3AF50C92",
    x"3AF4ACEC",
    x"3AF44D6B",
    x"3AF3EE0F",
    x"3AF38ED9",
    x"3AF32FC8",
    x"3AF2D0DC",
    x"3AF27215",
    x"3AF21372",
    x"3AF1B4F5",
    x"3AF1569D",
    x"3AF0F86A",
    x"3AF09A5B",
    x"3AF03C71",
    x"3AEFDEAC",
    x"3AEF810B",
    x"3AEF238F",
    x"3AEEC637",
    x"3AEE6904",
    x"3AEE0BF5",
    x"3AEDAF0B",
    x"3AED5244",
    x"3AECF5A2",
    x"3AEC9924",
    x"3AEC3CCB",
    x"3AEBE095",
    x"3AEB8483",
    x"3AEB2895",
    x"3AEACCCB",
    x"3AEA7125",
    x"3AEA15A3",
    x"3AE9BA44",
    x"3AE95F0A",
    x"3AE903F2",
    x"3AE8A8FE",
    x"3AE84E2E",
    x"3AE7F381",
    x"3AE798F8",
    x"3AE73E92",
    x"3AE6E44F",
    x"3AE68A2F",
    x"3AE63033",
    x"3AE5D65A",
    x"3AE57CA4",
    x"3AE52310",
    x"3AE4C9A0",
    x"3AE47053",
    x"3AE41728",
    x"3AE3BE21",
    x"3AE3653C",
    x"3AE30C7A",
    x"3AE2B3DA",
    x"3AE25B5D",
    x"3AE20303",
    x"3AE1AACB",
    x"3AE152B5",
    x"3AE0FAC2",
    x"3AE0A2F1",
    x"3AE04B43",
    x"3ADFF3B6",
    x"3ADF9C4C",
    x"3ADF4504",
    x"3ADEEDDE",
    x"3ADE96DA",
    x"3ADE3FF9",
    x"3ADDE939",
    x"3ADD929A",
    x"3ADD3C1E",
    x"3ADCE5C3",
    x"3ADC8F8A",
    x"3ADC3973",
    x"3ADBE37E",
    x"3ADB8DA9",
    x"3ADB37F7",
    x"3ADAE266",
    x"3ADA8CF6",
    x"3ADA37A8",
    x"3AD9E27A",
    x"3AD98D6F",
    x"3AD93884",
    x"3AD8E3BA",
    x"3AD88F12",
    x"3AD83A8B",
    x"3AD7E624",
    x"3AD791DF",
    x"3AD73DBA",
    x"3AD6E9B7",
    x"3AD695D4",
    x"3AD64212",
    x"3AD5EE70",
    x"3AD59AEF",
    x"3AD5478F",
    x"3AD4F44F",
    x"3AD4A130",
    x"3AD44E31",
    x"3AD3FB53",
    x"3AD3A895",
    x"3AD355F7",
    x"3AD3037A",
    x"3AD2B11D",
    x"3AD25EDF",
    x"3AD20CC2",
    x"3AD1BAC5",
    x"3AD168E8",
    x"3AD1172B",
    x"3AD0C58E",
    x"3AD07411",
    x"3AD022B4",
    x"3ACFD176",
    x"3ACF8058",
    x"3ACF2F5A",
    x"3ACEDE7B",
    x"3ACE8DBC",
    x"3ACE3D1C",
    x"3ACDEC9C",
    x"3ACD9C3B",
    x"3ACD4BFA",
    x"3ACCFBD8",
    x"3ACCABD5",
    x"3ACC5BF2",
    x"3ACC0C2D",
    x"3ACBBC88",
    x"3ACB6D02",
    x"3ACB1D9B",
    x"3ACACE53",
    x"3ACA7F2A",
    x"3ACA3020",
    x"3AC9E134",
    x"3AC99268",
    x"3AC943BA",
    x"3AC8F52B",
    x"3AC8A6BA",
    x"3AC85868",
    x"3AC80A35",
    x"3AC7BC20",
    x"3AC76E2A",
    x"3AC72052",
    x"3AC6D299",
    x"3AC684FE",
    x"3AC63781",
    x"3AC5EA22",
    x"3AC59CE2",
    x"3AC54FC0",
    x"3AC502BC",
    x"3AC4B5D6",
    x"3AC4690E",
    x"3AC41C64",
    x"3AC3CFD8",
    x"3AC38369",
    x"3AC33719",
    x"3AC2EAE6",
    x"3AC29ED1",
    x"3AC252DA",
    x"3AC20701",
    x"3AC1BB45",
    x"3AC16FA6",
    x"3AC12425",
    x"3AC0D8C2",
    x"3AC08D7C",
    x"3AC04253",
    x"3ABFF748",
    x"3ABFAC5A",
    x"3ABF618A",
    x"3ABF16D6",
    x"3ABECC40",
    x"3ABE81C6",
    x"3ABE376A",
    x"3ABDED2B",
    x"3ABDA309",
    x"3ABD5904",
    x"3ABD0F1B",
    x"3ABCC550",
    x"3ABC7BA1",
    x"3ABC320F",
    x"3ABBE89A",
    x"3ABB9F42",
    x"3ABB5606",
    x"3ABB0CE6",
    x"3ABAC3E4",
    x"3ABA7AFD",
    x"3ABA3233",
    x"3AB9E986",
    x"3AB9A0F5",
    x"3AB95880",
    x"3AB91028",
    x"3AB8C7EC",
    x"3AB87FCC",
    x"3AB837C8",
    x"3AB7EFE0",
    x"3AB7A814",
    x"3AB76065",
    x"3AB718D1",
    x"3AB6D159",
    x"3AB689FE",
    x"3AB642BE",
    x"3AB5FB99",
    x"3AB5B491",
    x"3AB56DA4",
    x"3AB526D3",
    x"3AB4E01E",
    x"3AB49984",
    x"3AB45306",
    x"3AB40CA3",
    x"3AB3C65C",
    x"3AB38030",
    x"3AB33A20",
    x"3AB2F42B",
    x"3AB2AE51",
    x"3AB26893",
    x"3AB222EF",
    x"3AB1DD67",
    x"3AB197FA",
    x"3AB152A9",
    x"3AB10D72",
    x"3AB0C856",
    x"3AB08355",
    x"3AB03E70",
    x"3AAFF9A5",
    x"3AAFB4F4",
    x"3AAF705F",
    x"3AAF2BE5",
    x"3AAEE785",
    x"3AAEA340",
    x"3AAE5F15",
    x"3AAE1B05",
    x"3AADD710",
    x"3AAD9335",
    x"3AAD4F75",
    x"3AAD0BCF",
    x"3AACC844",
    x"3AAC84D3",
    x"3AAC417C",
    x"3AABFE40",
    x"3AABBB1E",
    x"3AAB7816",
    x"3AAB3528",
    x"3AAAF254",
    x"3AAAAF9A",
    x"3AAA6CFB",
    x"3AAA2A75",
    x"3AA9E80A",
    x"3AA9A5B8",
    x"3AA96380",
    x"3AA92162",
    x"3AA8DF5E",
    x"3AA89D74",
    x"3AA85BA3",
    x"3AA819EC",
    x"3AA7D84F",
    x"3AA796CB",
    x"3AA75561",
    x"3AA71410",
    x"3AA6D2D9",
    x"3AA691BC",
    x"3AA650B7",
    x"3AA60FCD",
    x"3AA5CEFB",
    x"3AA58E43",
    x"3AA54DA4",
    x"3AA50D1E",
    x"3AA4CCB2",
    x"3AA48C5E",
    x"3AA44C24",
    x"3AA40C03",
    x"3AA3CBFB",
    x"3AA38C0B",
    x"3AA34C35",
    x"3AA30C78",
    x"3AA2CCD3",
    x"3AA28D48",
    x"3AA24DD5",
    x"3AA20E7B",
    x"3AA1CF3A",
    x"3AA19011",
    x"3AA15101",
    x"3AA1120A",
    x"3AA0D32B",
    x"3AA09465",
    x"3AA055B7",
    x"3AA01722",
    x"3A9FD8A5",
    x"3A9F9A40",
    x"3A9F5BF4",
    x"3A9F1DC1",
    x"3A9EDFA5",
    x"3A9EA1A2",
    x"3A9E63B7",
    x"3A9E25E4",
    x"3A9DE829",
    x"3A9DAA87",
    x"3A9D6CFC",
    x"3A9D2F89",
    x"3A9CF22F",
    x"3A9CB4EC",
    x"3A9C77C1",
    x"3A9C3AAF",
    x"3A9BFDB4",
    x"3A9BC0D0",
    x"3A9B8405",
    x"3A9B4751",
    x"3A9B0AB5",
    x"3A9ACE31",
    x"3A9A91C4",
    x"3A9A556F",
    x"3A9A1931",
    x"3A99DD0B",
    x"3A99A0FD",
    x"3A996506",
    x"3A992926",
    x"3A98ED5D",
    x"3A98B1AC",
    x"3A987613",
    x"3A983A90",
    x"3A97FF25",
    x"3A97C3D1",
    x"3A978894",
    x"3A974D6E",
    x"3A97125F",
    x"3A96D768",
    x"3A969C87",
    x"3A9661BD",
    x"3A96270B",
    x"3A95EC6F",
    x"3A95B1EA",
    x"3A95777C",
    x"3A953D25",
    x"3A9502E4",
    x"3A94C8BA",
    x"3A948EA7",
    x"3A9454AB",
    x"3A941AC5",
    x"3A93E0F6",
    x"3A93A73D",
    x"3A936D9B",
    x"3A933410",
    x"3A92FA9B",
    x"3A92C13C",
    x"3A9287F4",
    x"3A924EC2",
    x"3A9215A6",
    x"3A91DCA1",
    x"3A91A3B2",
    x"3A916AD9",
    x"3A913216",
    x"3A90F96A",
    x"3A90C0D3",
    x"3A908853",
    x"3A904FE9",
    x"3A901795",
    x"3A8FDF56",
    x"3A8FA72E",
    x"3A8F6F1C",
    x"3A8F371F",
    x"3A8EFF39",
    x"3A8EC768",
    x"3A8E8FAD",
    x"3A8E5808",
    x"3A8E2078",
    x"3A8DE8FE",
    x"3A8DB19A",
    x"3A8D7A4B",
    x"3A8D4312",
    x"3A8D0BEF",
    x"3A8CD4E1",
    x"3A8C9DE9",
    x"3A8C6706",
    x"3A8C3038",
    x"3A8BF980",
    x"3A8BC2DD",
    x"3A8B8C50",
    x"3A8B55D8",
    x"3A8B1F75",
    x"3A8AE927",
    x"3A8AB2EF",
    x"3A8A7CCB",
    x"3A8A46BD",
    x"3A8A10C4",
    x"3A89DAE0",
    x"3A89A511",
    x"3A896F57",
    x"3A8939B2",
    x"3A890422",
    x"3A88CEA7",
    x"3A889940",
    x"3A8863EF",
    x"3A882EB2",
    x"3A87F98B",
    x"3A87C477",
    x"3A878F79",
    x"3A875A8F",
    x"3A8725BA",
    x"3A86F0FA",
    x"3A86BC4E",
    x"3A8687B7",
    x"3A865334",
    x"3A861EC6",
    x"3A85EA6C",
    x"3A85B627",
    x"3A8581F6",
    x"3A854DD9",
    x"3A8519D1",
    x"3A84E5DD",
    x"3A84B1FD",
    x"3A847E32",
    x"3A844A7B",
    x"3A8416D8",
    x"3A83E349",
    x"3A83AFCE",
    x"3A837C67",
    x"3A834915",
    x"3A8315D6",
    x"3A82E2AC",
    x"3A82AF95",
    x"3A827C93",
    x"3A8249A4",
    x"3A8216C9",
    x"3A81E402",
    x"3A81B14F",
    x"3A817EAF",
    x"3A814C24",
    x"3A8119AC",
    x"3A80E748",
    x"3A80B4F7",
    x"3A8082BA",
    x"3A805091",
    x"3A801E7B",
    x"3A7FD8F3",
    x"3A7F7515",
    x"3A7F115F",
    x"3A7EADD0",
    x"3A7E4A67",
    x"3A7DE726",
    x"3A7D840B",
    x"3A7D2117",
    x"3A7CBE49",
    x"3A7C5BA2",
    x"3A7BF921",
    x"3A7B96C7",
    x"3A7B3493",
    x"3A7AD286",
    x"3A7A709F",
    x"3A7A0EDE",
    x"3A79AD43",
    x"3A794BCF",
    x"3A78EA80",
    x"3A788957",
    x"3A782855",
    x"3A77C778",
    x"3A7766C1",
    x"3A770630",
    x"3A76A5C4",
    x"3A76457E",
    x"3A75E55E",
    x"3A758563",
    x"3A75258E",
    x"3A74C5DE",
    x"3A746653",
    x"3A7406EE",
    x"3A73A7AD",
    x"3A734893",
    x"3A72E99D",
    x"3A728ACC",
    x"3A722C20",
    x"3A71CD9A",
    x"3A716F38",
    x"3A7110FB",
    x"3A70B2E2",
    x"3A7054EF",
    x"3A6FF720",
    x"3A6F9976",
    x"3A6F3BF0",
    x"3A6EDE8F",
    x"3A6E8152",
    x"3A6E243A",
    x"3A6DC746",
    x"3A6D6A76",
    x"3A6D0DCB",
    x"3A6CB143",
    x"3A6C54E0",
    x"3A6BF8A1",
    x"3A6B9C86",
    x"3A6B408F",
    x"3A6AE4BB",
    x"3A6A890C",
    x"3A6A2D80",
    x"3A69D218",
    x"3A6976D4",
    x"3A691BB4",
    x"3A68C0B7",
    x"3A6865DD",
    x"3A680B27",
    x"3A67B094",
    x"3A675625",
    x"3A66FBD9",
    x"3A66A1B0",
    x"3A6647AB",
    x"3A65EDC8",
    x"3A659409",
    x"3A653A6D",
    x"3A64E0F3",
    x"3A64879D",
    x"3A642E69",
    x"3A63D559",
    x"3A637C6B",
    x"3A63239F",
    x"3A62CAF7",
    x"3A627271",
    x"3A621A0D",
    x"3A61C1CC",
    x"3A6169AE",
    x"3A6111B2",
    x"3A60B9D8",
    x"3A606221",
    x"3A600A8B",
    x"3A5FB318",
    x"3A5F5BC7",
    x"3A5F0499",
    x"3A5EAD8C",
    x"3A5E56A1",
    x"3A5DFFD8",
    x"3A5DA931",
    x"3A5D52AC",
    x"3A5CFC49",
    x"3A5CA607",
    x"3A5C4FE7",
    x"3A5BF9E8",
    x"3A5BA40C",
    x"3A5B4E50",
    x"3A5AF8B6",
    x"3A5AA33E",
    x"3A5A4DE7",
    x"3A59F8B1",
    x"3A59A39C",
    x"3A594EA9",
    x"3A58F9D7",
    x"3A58A526",
    x"3A585096",
    x"3A57FC27",
    x"3A57A7D9",
    x"3A5753AC",
    x"3A56FFA0",
    x"3A56ABB4",
    x"3A5657E9",
    x"3A56043F",
    x"3A55B0B6",
    x"3A555D4D",
    x"3A550A05",
    x"3A54B6DD",
    x"3A5463D6",
    x"3A5410EF",
    x"3A53BE29",
    x"3A536B83",
    x"3A5318FD",
    x"3A52C697",
    x"3A527452",
    x"3A52222C",
    x"3A51D027",
    x"3A517E42",
    x"3A512C7C",
    x"3A50DAD7",
    x"3A508951",
    x"3A5037EC",
    x"3A4FE6A6",
    x"3A4F9580",
    x"3A4F4479",
    x"3A4EF392",
    x"3A4EA2CB",
    x"3A4E5223",
    x"3A4E019A",
    x"3A4DB132",
    x"3A4D60E8",
    x"3A4D10BE",
    x"3A4CC0B3",
    x"3A4C70C7",
    x"3A4C20FB",
    x"3A4BD14E",
    x"3A4B81BF",
    x"3A4B3250",
    x"3A4AE300",
    x"3A4A93CF",
    x"3A4A44BC",
    x"3A49F5C9",
    x"3A49A6F4",
    x"3A49583F",
    x"3A4909A7",
    x"3A48BB2F",
    x"3A486CD5",
    x"3A481E9A",
    x"3A47D07D",
    x"3A47827F",
    x"3A47349F",
    x"3A46E6DE",
    x"3A46993B",
    x"3A464BB6",
    x"3A45FE50",
    x"3A45B108",
    x"3A4563DD",
    x"3A4516D2",
    x"3A44C9E4",
    x"3A447D14",
    x"3A443062",
    x"3A43E3CE",
    x"3A439758",
    x"3A434B00",
    x"3A42FEC5",
    x"3A42B2A9",
    x"3A4266AA",
    x"3A421AC8",
    x"3A41CF05",
    x"3A41835F",
    x"3A4137D6",
    x"3A40EC6B",
    x"3A40A11D",
    x"3A4055ED",
    x"3A400ADA",
    x"3A3FBFE5",
    x"3A3F750C",
    x"3A3F2A51",
    x"3A3EDFB3",
    x"3A3E9532",
    x"3A3E4ACF",
    x"3A3E0088",
    x"3A3DB65E",
    x"3A3D6C51",
    x"3A3D2262",
    x"3A3CD88F",
    x"3A3C8ED8",
    x"3A3C453F",
    x"3A3BFBC2",
    x"3A3BB262",
    x"3A3B691F",
    x"3A3B1FF8",
    x"3A3AD6EE",
    x"3A3A8E00",
    x"3A3A452F",
    x"3A39FC7A",
    x"3A39B3E2",
    x"3A396B66",
    x"3A392306",
    x"3A38DAC2",
    x"3A38929B",
    x"3A384A90",
    x"3A3802A1",
    x"3A37BACE",
    x"3A377317",
    x"3A372B7C",
    x"3A36E3FD",
    x"3A369C9A",
    x"3A365552",
    x"3A360E27",
    x"3A35C717",
    x"3A358023",
    x"3A35394B",
    x"3A34F28F",
    x"3A34ABEE",
    x"3A346568",
    x"3A341EFE",
    x"3A33D8B0",
    x"3A33927D",
    x"3A334C66",
    x"3A330669",
    x"3A32C089",
    x"3A327AC3",
    x"3A323519",
    x"3A31EF89",
    x"3A31AA15",
    x"3A3164BD",
    x"3A311F7F",
    x"3A30DA5C",
    x"3A309554",
    x"3A305067",
    x"3A300B95",
    x"3A2FC6DE",
    x"3A2F8242",
    x"3A2F3DC0",
    x"3A2EF95A",
    x"3A2EB50E",
    x"3A2E70DC",
    x"3A2E2CC5",
    x"3A2DE8C9",
    x"3A2DA4E8",
    x"3A2D6120",
    x"3A2D1D74",
    x"3A2CD9E1",
    x"3A2C9669",
    x"3A2C530C",
    x"3A2C0FC9",
    x"3A2BCC9F",
    x"3A2B8991",
    x"3A2B469C",
    x"3A2B03C1",
    x"3A2AC101",
    x"3A2A7E5B",
    x"3A2A3BCE",
    x"3A29F95C",
    x"3A29B703",
    x"3A2974C5",
    x"3A2932A0",
    x"3A28F095",
    x"3A28AEA4",
    x"3A286CCD",
    x"3A282B0F",
    x"3A27E96B",
    x"3A27A7E1",
    x"3A276670",
    x"3A272519",
    x"3A26E3DB",
    x"3A26A2B7",
    x"3A2661AC",
    x"3A2620BB",
    x"3A25DFE2",
    x"3A259F24",
    x"3A255E7E",
    x"3A251DF2",
    x"3A24DD7F",
    x"3A249D25",
    x"3A245CE4",
    x"3A241CBC",
    x"3A23DCAD",
    x"3A239CB8",
    x"3A235CDB",
    x"3A231D17",
    x"3A22DD6C",
    x"3A229DDA",
    x"3A225E61",
    x"3A221F00",
    x"3A21DFB9",
    x"3A21A08A",
    x"3A216173",
    x"3A212275",
    x"3A20E390",
    x"3A20A4C4",
    x"3A206610",
    x"3A202774",
    x"3A1FE8F1",
    x"3A1FAA86",
    x"3A1F6C33",
    x"3A1F2DF9",
    x"3A1EEFD8",
    x"3A1EB1CE",
    x"3A1E73DD",
    x"3A1E3603",
    x"3A1DF842",
    x"3A1DBA99",
    x"3A1D7D09",
    x"3A1D3F90",
    x"3A1D022F",
    x"3A1CC4E6",
    x"3A1C87B5",
    x"3A1C4A9C",
    x"3A1C0D9B",
    x"3A1BD0B1",
    x"3A1B93E0",
    x"3A1B5726",
    x"3A1B1A84",
    x"3A1ADDF9",
    x"3A1AA186",
    x"3A1A652B",
    x"3A1A28E7",
    x"3A19ECBB",
    x"3A19B0A6",
    x"3A1974A9",
    x"3A1938C3",
    x"3A18FCF5",
    x"3A18C13D",
    x"3A18859E",
    x"3A184A15",
    x"3A180EA4",
    x"3A17D34A",
    x"3A179807",
    x"3A175CDB",
    x"3A1721C6",
    x"3A16E6C8",
    x"3A16ABE2",
    x"3A167112",
    x"3A163659",
    x"3A15FBB8",
    x"3A15C12D",
    x"3A1586B9",
    x"3A154C5C",
    x"3A151215",
    x"3A14D7E5",
    x"3A149DCC",
    x"3A1463CA",
    x"3A1429DE",
    x"3A13F009",
    x"3A13B64B",
    x"3A137CA3",
    x"3A134311",
    x"3A130997",
    x"3A12D032",
    x"3A1296E4",
    x"3A125DAC",
    x"3A12248B",
    x"3A11EB80",
    x"3A11B28B",
    x"3A1179AC",
    x"3A1140E4",
    x"3A110831",
    x"3A10CF95",
    x"3A10970F",
    x"3A105E9F",
    x"3A102645",
    x"3A0FEE01",
    x"3A0FB5D3",
    x"3A0F7DBB",
    x"3A0F45B9",
    x"3A0F0DCD",
    x"3A0ED5F6",
    x"3A0E9E36",
    x"3A0E668B",
    x"3A0E2EF5",
    x"3A0DF776",
    x"3A0DC00C",
    x"3A0D88B8",
    x"3A0D5179",
    x"3A0D1A50",
    x"3A0CE33D",
    x"3A0CAC3F",
    x"3A0C7556",
    x"3A0C3E83",
    x"3A0C07C5",
    x"3A0BD11D",
    x"3A0B9A8A",
    x"3A0B640C",
    x"3A0B2DA4",
    x"3A0AF750",
    x"3A0AC112",
    x"3A0A8AEA",
    x"3A0A54D6",
    x"3A0A1ED7",
    x"3A09E8EE",
    x"3A09B319",
    x"3A097D5A",
    x"3A0947AF",
    x"3A09121A",
    x"3A08DC99",
    x"3A08A72E",
    x"3A0871D7",
    x"3A083C95",
    x"3A080767",
    x"3A07D24F",
    x"3A079D4B",
    x"3A07685C",
    x"3A073381",
    x"3A06FEBC",
    x"3A06CA0A",
    x"3A06956E",
    x"3A0660E6",
    x"3A062C72",
    x"3A05F813",
    x"3A05C3C8",
    x"3A058F92",
    x"3A055B70",
    x"3A052763",
    x"3A04F369",
    x"3A04BF84",
    x"3A048BB4",
    x"3A0457F7",
    x"3A04244F",
    x"3A03F0BB",
    x"3A03BD3B",
    x"3A0389CF",
    x"3A035677",
    x"3A032333",
    x"3A02F004",
    x"3A02BCE8",
    x"3A0289E0",
    x"3A0256EC",
    x"3A02240C",
    x"3A01F140",
    x"3A01BE88",
    x"3A018BE3",
    x"3A015952",
    x"3A0126D5",
    x"3A00F46C",
    x"3A00C216",
    x"3A008FD4",
    x"3A005DA6",
    x"3A002B8B",
    x"39FFF308",
    x"39FF8F21",
    x"39FF2B60",
    x"39FEC7C7",
    x"39FE6454",
    x"39FE0108",
    x"39FD9DE3",
    x"39FD3AE5",
    x"39FCD80D",
    x"39FC755C",
    x"39FC12D1",
    x"39FBB06D",
    x"39FB4E30",
    x"39FAEC18",
    x"39FA8A27",
    x"39FA285C",
    x"39F9C6B8",
    x"39F96539",
    x"39F903E1",
    x"39F8A2AE",
    x"39F841A1",
    x"39F7E0BB",
    x"39F77FFA",
    x"39F71F5F",
    x"39F6BEE9",
    x"39F65E9A",
    x"39F5FE6F",
    x"39F59E6B",
    x"39F53E8C",
    x"39F4DED2",
    x"39F47F3D",
    x"39F41FCE",
    x"39F3C085",
    x"39F36160",
    x"39F30261",
    x"39F2A386",
    x"39F244D1",
    x"39F1E640",
    x"39F187D5",
    x"39F1298E",
    x"39F0CB6C",
    x"39F06D6F",
    x"39F00F97",
    x"39EFB1E3",
    x"39EF5454",
    x"39EEF6E9",
    x"39EE99A3",
    x"39EE3C81",
    x"39EDDF84",
    x"39ED82AA",
    x"39ED25F6",
    x"39ECC965",
    x"39EC6CF8",
    x"39EC10B0",
    x"39EBB48B",
    x"39EB588B",
    x"39EAFCAE",
    x"39EAA0F5",
    x"39EA4560",
    x"39E9E9EF",
    x"39E98EA1",
    x"39E93377",
    x"39E8D871",
    x"39E87D8E",
    x"39E822CF",
    x"39E7C833",
    x"39E76DBB",
    x"39E71365",
    x"39E6B933",
    x"39E65F25",
    x"39E60539",
    x"39E5AB71",
    x"39E551CB",
    x"39E4F849",
    x"39E49EE9",
    x"39E445AD",
    x"39E3EC93",
    x"39E3939C",
    x"39E33AC7",
    x"39E2E216",
    x"39E28987",
    x"39E2311A",
    x"39E1D8D0",
    x"39E180A9",
    x"39E128A4",
    x"39E0D0C1",
    x"39E07901",
    x"39E02163",
    x"39DFC9E7",
    x"39DF728D",
    x"39DF1B55",
    x"39DEC43F",
    x"39DE6D4C",
    x"39DE167A",
    x"39DDBFCA",
    x"39DD693C",
    x"39DD12D0",
    x"39DCBC85",
    x"39DC665D",
    x"39DC1055",
    x"39DBBA70",
    x"39DB64AC",
    x"39DB0F09",
    x"39DAB988",
    x"39DA6428",
    x"39DA0EEA",
    x"39D9B9CD",
    x"39D964D1",
    x"39D90FF6",
    x"39D8BB3C",
    x"39D866A4",
    x"39D8122C",
    x"39D7BDD5",
    x"39D769A0",
    x"39D7158B",
    x"39D6C197",
    x"39D66DC4",
    x"39D61A11",
    x"39D5C67F",
    x"39D5730E",
    x"39D51FBD",
    x"39D4CC8D",
    x"39D4797D",
    x"39D4268E",
    x"39D3D3BF",
    x"39D38111",
    x"39D32E82",
    x"39D2DC14",
    x"39D289C6",
    x"39D23799",
    x"39D1E58B",
    x"39D1939D",
    x"39D141D0",
    x"39D0F022",
    x"39D09E94",
    x"39D04D26",
    x"39CFFBD8",
    x"39CFAAA9",
    x"39CF599A",
    x"39CF08AB",
    x"39CEB7DC",
    x"39CE672C",
    x"39CE169B",
    x"39CDC62A",
    x"39CD75D8",
    x"39CD25A6",
    x"39CCD593",
    x"39CC859F",
    x"39CC35CA",
    x"39CBE615",
    x"39CB967F",
    x"39CB4707",
    x"39CAF7AF",
    x"39CAA876",
    x"39CA595B",
    x"39CA0A60",
    x"39C9BB83",
    x"39C96CC5",
    x"39C91E26",
    x"39C8CFA6",
    x"39C88144",
    x"39C83301",
    x"39C7E4DC",
    x"39C796D6",
    x"39C748EE",
    x"39C6FB25",
    x"39C6AD7A",
    x"39C65FEE",
    x"39C6127F",
    x"39C5C52F",
    x"39C577FD",
    x"39C52AE9",
    x"39C4DDF4",
    x"39C4911C",
    x"39C44462",
    x"39C3F7C6",
    x"39C3AB49",
    x"39C35EE9",
    x"39C312A6",
    x"39C2C682",
    x"39C27A7B",
    x"39C22E92",
    x"39C1E2C7",
    x"39C19719",
    x"39C14B89",
    x"39C10016",
    x"39C0B4C1",
    x"39C06989",
    x"39C01E6E",
    x"39BFD371",
    x"39BF8891",
    x"39BF3DCE",
    x"39BEF329",
    x"39BEA8A0",
    x"39BE5E35",
    x"39BE13E7",
    x"39BDC9B6",
    x"39BD7FA1",
    x"39BD35AA",
    x"39BCEBCF",
    x"39BCA212",
    x"39BC5871",
    x"39BC0EEC",
    x"39BBC585",
    x"39BB7C3A",
    x"39BB330C",
    x"39BAE9FA",
    x"39BAA105",
    x"39BA582C",
    x"39BA0F70",
    x"39B9C6D0",
    x"39B97E4D",
    x"39B935E6",
    x"39B8ED9B",
    x"39B8A56C",
    x"39B85D59",
    x"39B81563",
    x"39B7CD89",
    x"39B785CA",
    x"39B73E28",
    x"39B6F6A2",
    x"39B6AF38",
    x"39B667E9",
    x"39B620B6",
    x"39B5D99F",
    x"39B592A4",
    x"39B54BC5",
    x"39B50501",
    x"39B4BE59",
    x"39B477CC",
    x"39B4315B",
    x"39B3EB06",
    x"39B3A4CC",
    x"39B35EAD",
    x"39B318AA",
    x"39B2D2C2",
    x"39B28CF5",
    x"39B24744",
    x"39B201AD",
    x"39B1BC32",
    x"39B176D2",
    x"39B1318D",
    x"39B0EC64",
    x"39B0A755",
    x"39B06261",
    x"39B01D88",
    x"39AFD8CA",
    x"39AF9426",
    x"39AF4F9E",
    x"39AF0B30",
    x"39AEC6DD",
    x"39AE82A5",
    x"39AE3E87",
    x"39ADFA84",
    x"39ADB69B",
    x"39AD72CD",
    x"39AD2F1A",
    x"39ACEB81",
    x"39ACA802",
    x"39AC649D",
    x"39AC2153",
    x"39ABDE23",
    x"39AB9B0E",
    x"39AB5812",
    x"39AB1531",
    x"39AAD26A",
    x"39AA8FBC",
    x"39AA4D29",
    x"39AA0AB0",
    x"39A9C851",
    x"39A9860C",
    x"39A943E0",
    x"39A901CF",
    x"39A8BFD7",
    x"39A87DF9",
    x"39A83C34",
    x"39A7FA8A",
    x"39A7B8F9",
    x"39A77781",
    x"39A73623",
    x"39A6F4DF",
    x"39A6B3B4",
    x"39A672A2",
    x"39A631AA",
    x"39A5F0CC",
    x"39A5B006",
    x"39A56F5A",
    x"39A52EC7",
    x"39A4EE4D",
    x"39A4ADED",
    x"39A46DA6",
    x"39A42D77",
    x"39A3ED62",
    x"39A3AD66",
    x"39A36D83",
    x"39A32DB8",
    x"39A2EE07",
    x"39A2AE6E",
    x"39A26EEF",
    x"39A22F88",
    x"39A1F039",
    x"39A1B104",
    x"39A171E7",
    x"39A132E3",
    x"39A0F3F7",
    x"39A0B524",
    x"39A0766A",
    x"39A037C8",
    x"399FF93E",
    x"399FBACD",
    x"399F7C74",
    x"399F3E34",
    x"399F000C",
    x"399EC1FC",
    x"399E8404",
    x"399E4625",
    x"399E085D",
    x"399DCAAE",
    x"399D8D17",
    x"399D4F98",
    x"399D1231",
    x"399CD4E2",
    x"399C97AA",
    x"399C5A8B",
    x"399C1D84",
    x"399BE094",
    x"399BA3BC",
    x"399B66FC",
    x"399B2A54",
    x"399AEDC3",
    x"399AB14A",
    x"399A74E8",
    x"399A389F",
    x"3999FC6C",
    x"3999C051",
    x"3999844E",
    x"39994862",
    x"39990C8D",
    x"3998D0D0",
    x"3998952A",
    x"3998599C",
    x"39981E24",
    x"3997E2C4",
    x"3997A77B",
    x"39976C49",
    x"3997312E",
    x"3996F62B",
    x"3996BB3E",
    x"39968068",
    x"399645AA",
    x"39960B02",
    x"3995D071",
    x"399595F7",
    x"39955B94",
    x"39952148",
    x"3994E712",
    x"3994ACF3",
    x"399472EB",
    x"399438F9",
    x"3993FF1E",
    x"3993C55A",
    x"39938BAC",
    x"39935215",
    x"39931894",
    x"3992DF2A",
    x"3992A5D6",
    x"39926C98",
    x"39923371",
    x"3991FA60",
    x"3991C165",
    x"39918881",
    x"39914FB3",
    x"399116FA",
    x"3990DE59",
    x"3990A5CD",
    x"39906D57",
    x"399034F7",
    x"398FFCAE",
    x"398FC47A",
    x"398F8C5C",
    x"398F5454",
    x"398F1C62",
    x"398EE486",
    x"398EACC0",
    x"398E750F",
    x"398E3D74",
    x"398E05EF",
    x"398DCE80",
    x"398D9726",
    x"398D5FE1",
    x"398D28B3",
    x"398CF19A",
    x"398CBA96",
    x"398C83A8",
    x"398C4CCF",
    x"398C160C",
    x"398BDF5E",
    x"398BA8C5",
    x"398B7242",
    x"398B3BD4",
    x"398B057B",
    x"398ACF38",
    x"398A9909",
    x"398A62F0",
    x"398A2CEC",
    x"3989F6FD",
    x"3989C123",
    x"39898B5E",
    x"398955AE",
    x"39892013",
    x"3988EA8D",
    x"3988B51C",
    x"39887FC0",
    x"39884A78",
    x"39881546",
    x"3987E028",
    x"3987AB1E",
    x"3987762A",
    x"3987414A",
    x"39870C7F",
    x"3986D7C8",
    x"3986A326",
    x"39866E99",
    x"39863A20",
    x"398605BB",
    x"3985D16B",
    x"39859D30",
    x"39856909",
    x"398534F6",
    x"398500F7",
    x"3984CD0D",
    x"39849937",
    x"39846575",
    x"398431C8",
    x"3983FE2E",
    x"3983CAA9",
    x"39839738",
    x"398363DB",
    x"39833092",
    x"3982FD5D",
    x"3982CA3C",
    x"3982972F",
    x"39826436",
    x"39823151",
    x"3981FE7F",
    x"3981CBC2",
    x"39819918",
    x"39816682",
    x"39813400",
    x"39810192",
    x"3980CF37",
    x"39809CF0",
    x"39806ABC",
    x"3980389C",
    x"39800690",
    x"397FA92E",
    x"397F4564",
    x"397EE1C0",
    x"397E7E43",
    x"397E1AED",
    x"397DB7BE",
    x"397D54B6",
    x"397CF1D4",
    x"397C8F19",
    x"397C2C84",
    x"397BCA16",
    x"397B67CE",
    x"397B05AD",
    x"397AA3B2",
    x"397A41DD",
    x"3979E02E",
    x"39797EA6",
    x"39791D44",
    x"3978BC07",
    x"39785AF1",
    x"3977FA00",
    x"39779935",
    x"39773890",
    x"3976D811",
    x"397677B7",
    x"39761784",
    x"3975B775",
    x"3975578C",
    x"3974F7C9",
    x"3974982B",
    x"397438B2",
    x"3973D95E",
    x"39737A30",
    x"39731B27",
    x"3972BC43",
    x"39725D84",
    x"3971FEEA",
    x"3971A075",
    x"39714224",
    x"3970E3F9",
    x"397085F2",
    x"39702810",
    x"396FCA53",
    x"396F6CBA",
    x"396F0F46",
    x"396EB1F6",
    x"396E54CB",
    x"396DF7C4",
    x"396D9AE1",
    x"396D3E23",
    x"396CE189",
    x"396C8513",
    x"396C28C1",
    x"396BCC93",
    x"396B7089",
    x"396B14A3",
    x"396AB8E1",
    x"396A5D42",
    x"396A01C8",
    x"3969A671",
    x"39694B3E",
    x"3968F02E",
    x"39689542",
    x"39683A7A",
    x"3967DFD4",
    x"39678553",
    x"39672AF4",
    x"3966D0B9",
    x"396676A1",
    x"39661CAC",
    x"3965C2DB",
    x"3965692C",
    x"39650FA1",
    x"3964B638",
    x"39645CF2",
    x"396403CF",
    x"3963AACF",
    x"396351F2",
    x"3962F937",
    x"3962A09F",
    x"3962482A",
    x"3961EFD7",
    x"396197A6",
    x"39613F98",
    x"3960E7AD",
    x"39608FE3",
    x"3960383C",
    x"395FE0B7",
    x"395F8955",
    x"395F3214",
    x"395EDAF5",
    x"395E83F9",
    x"395E2D1E",
    x"395DD666",
    x"395D7FCF",
    x"395D295A",
    x"395CD306",
    x"395C7CD5",
    x"395C26C5",
    x"395BD0D7",
    x"395B7B0A",
    x"395B255E",
    x"395ACFD5",
    x"395A7A6C",
    x"395A2525",
    x"3959CFFF",
    x"39597AFA",
    x"39592617",
    x"3958D155",
    x"39587CB3",
    x"39582833",
    x"3957D3D4",
    x"39577F96",
    x"39572B78",
    x"3956D77C",
    x"395683A0",
    x"39562FE5",
    x"3955DC4A",
    x"395588D1",
    x"39553578",
    x"3954E23F",
    x"39548F27",
    x"39543C2F",
    x"3953E958",
    x"395396A1",
    x"3953440A",
    x"3952F194",
    x"39529F3D",
    x"39524D07",
    x"3951FAF1",
    x"3951A8FB",
    x"39515725",
    x"3951056F",
    x"3950B3D9",
    x"39506262",
    x"3950110C",
    x"394FBFD5",
    x"394F6EBE",
    x"394F1DC7",
    x"394ECCEF",
    x"394E7C36",
    x"394E2B9E",
    x"394DDB24",
    x"394D8ACA",
    x"394D3A90",
    x"394CEA75",
    x"394C9A79",
    x"394C4A9C",
    x"394BFADE",
    x"394BAB40",
    x"394B5BC1",
    x"394B0C60",
    x"394ABD1F",
    x"394A6DFD",
    x"394A1EF9",
    x"3949D014",
    x"3949814E",
    x"394932A7",
    x"3948E41F",
    x"394895B5",
    x"3948476A",
    x"3947F93D",
    x"3947AB2F",
    x"39475D3F",
    x"39470F6E",
    x"3946C1BB",
    x"39467427",
    x"394626B1",
    x"3945D959",
    x"39458C1F",
    x"39453F03",
    x"3944F206",
    x"3944A526",
    x"39445865",
    x"39440BC1",
    x"3943BF3B",
    x"394372D4",
    x"3943268A",
    x"3942DA5D",
    x"39428E4F",
    x"3942425E",
    x"3941F68B",
    x"3941AAD6",
    x"39415F3E",
    x"394113C3",
    x"3940C866",
    x"39407D27",
    x"39403204",
    x"393FE700",
    x"393F9C18",
    x"393F514E",
    x"393F06A0",
    x"393EBC10",
    x"393E719D",
    x"393E2748",
    x"393DDD0F",
    x"393D92F3",
    x"393D48F4",
    x"393CFF12",
    x"393CB54D",
    x"393C6BA4",
    x"393C2219",
    x"393BD8AA",
    x"393B8F57",
    x"393B4622",
    x"393AFD08",
    x"393AB40C",
    x"393A6B2C",
    x"393A2268",
    x"3939D9C1",
    x"39399136",
    x"393948C7",
    x"39390075",
    x"3938B83F",
    x"39387025",
    x"39382827",
    x"3937E046",
    x"39379880",
    x"393750D7",
    x"39370949",
    x"3936C1D7",
    x"39367A82",
    x"39363348",
    x"3935EC2A",
    x"3935A527",
    x"39355E40",
    x"39351775",
    x"3934D0C6",
    x"39348A32",
    x"393443BA",
    x"3933FD5D",
    x"3933B71C",
    x"393370F6",
    x"39332AEC",
    x"3932E4FD",
    x"39329F29",
    x"39325970",
    x"393213D3",
    x"3931CE51",
    x"393188EA",
    x"3931439E",
    x"3930FE6D",
    x"3930B957",
    x"3930745C",
    x"39302F7C",
    x"392FEAB7",
    x"392FA60D",
    x"392F617D",
    x"392F1D09",
    x"392ED8AF",
    x"392E946F",
    x"392E504B",
    x"392E0C41",
    x"392DC851",
    x"392D847C",
    x"392D40C2",
    x"392CFD22",
    x"392CB99C",
    x"392C7631",
    x"392C32E0",
    x"392BEFA9",
    x"392BAC8C",
    x"392B698A",
    x"392B26A2",
    x"392AE3D4",
    x"392AA120",
    x"392A5E86",
    x"392A1C06",
    x"3929D9A0",
    x"39299754",
    x"39295522",
    x"39291309",
    x"3928D10B",
    x"39288F26",
    x"39284D5B",
    x"39280BAA",
    x"3927CA12",
    x"39278894",
    x"3927472F",
    x"392705E4",
    x"3926C4B3",
    x"3926839A",
    x"3926429C",
    x"392601B6",
    x"3925C0EA",
    x"39258038",
    x"39253F9E",
    x"3924FF1E",
    x"3924BEB7",
    x"39247E69",
    x"39243E34",
    x"3923FE18",
    x"3923BE16",
    x"39237E2C",
    x"39233E5B",
    x"3922FEA3",
    x"3922BF04",
    x"39227F7E",
    x"39224010",
    x"392200BC",
    x"3921C180",
    x"3921825D",
    x"39214352",
    x"39210460",
    x"3920C587",
    x"392086C6",
    x"3920481D",
    x"3920098D",
    x"391FCB16",
    x"391F8CB7",
    x"391F4E70",
    x"391F1041",
    x"391ED22B",
    x"391E942D",
    x"391E5647",
    x"391E187A",
    x"391DDAC4",
    x"391D9D27",
    x"391D5FA1",
    x"391D2234",
    x"391CE4DF",
    x"391CA7A1",
    x"391C6A7C",
    x"391C2D6E",
    x"391BF078",
    x"391BB39A",
    x"391B76D4",
    x"391B3A25",
    x"391AFD8E",
    x"391AC10F",
    x"391A84A8",
    x"391A4858",
    x"391A0C1F",
    x"3919CFFE",
    x"391993F5",
    x"39195802",
    x"39191C28",
    x"3918E064",
    x"3918A4B8",
    x"39186924",
    x"39182DA6",
    x"3917F240",
    x"3917B6F1",
    x"39177BB9",
    x"39174098",
    x"3917058F",
    x"3916CA9C",
    x"39168FC0",
    x"391654FC",
    x"39161A4E",
    x"3915DFB7",
    x"3915A537",
    x"39156ACE",
    x"3915307C",
    x"3914F640",
    x"3914BC1B",
    x"3914820D",
    x"39144816",
    x"39140E35",
    x"3913D46B",
    x"39139AB7",
    x"3913611A",
    x"39132793",
    x"3912EE23",
    x"3912B4C9",
    x"39127B86",
    x"39124258",
    x"39120942",
    x"3911D041",
    x"39119757",
    x"39115E83",
    x"391125C5",
    x"3910ED1D",
    x"3910B48C",
    x"39107C10",
    x"391043AB",
    x"39100B5C",
    x"390FD322",
    x"390F9AFF",
    x"390F62F1",
    x"390F2AF9",
    x"390EF317",
    x"390EBB4B",
    x"390E8395",
    x"390E4BF5",
    x"390E146A",
    x"390DDCF5",
    x"390DA595",
    x"390D6E4B",
    x"390D3717",
    x"390CFFF8",
    x"390CC8EF",
    x"390C91FB",
    x"390C5B1D",
    x"390C2454",
    x"390BEDA0",
    x"390BB702",
    x"390B8079",
    x"390B4A06",
    x"390B13A8",
    x"390ADD5F",
    x"390AA72B",
    x"390A710C",
    x"390A3B02",
    x"390A050E",
    x"3909CF2E",
    x"39099964",
    x"390963AF",
    x"39092E0E",
    x"3908F883",
    x"3908C30C",
    x"39088DAA",
    x"3908585D",
    x"39082325",
    x"3907EE02",
    x"3907B8F3",
    x"390783F9",
    x"39074F14",
    x"39071A43",
    x"3906E588",
    x"3906B0E0",
    x"39067C4D",
    x"390647CF",
    x"39061365",
    x"3905DF10",
    x"3905AACF",
    x"390576A2",
    x"3905428A",
    x"39050E86",
    x"3904DA97",
    x"3904A6BC",
    x"390472F5",
    x"39043F42",
    x"39040BA3",
    x"3903D819",
    x"3903A4A2",
    x"39037140",
    x"39033DF2",
    x"39030AB8",
    x"3902D791",
    x"3902A47F",
    x"39027181",
    x"39023E97",
    x"39020BC0",
    x"3901D8FD",
    x"3901A64F",
    x"390173B3",
    x"3901412C",
    x"39010EB9",
    x"3900DC59",
    x"3900AA0C",
    x"390077D4",
    x"390045AF",
    x"3900139D",
    x"38FFC33F",
    x"38FF5F6A",
    x"38FEFBBC",
    x"38FE9835",
    x"38FE34D5",
    x"38FDD19C",
    x"38FD6E8A",
    x"38FD0B9E",
    x"38FCA8D8",
    x"38FC463A",
    x"38FBE3C2",
    x"38FB8170",
    x"38FB1F44",
    x"38FABD3F",
    x"38FA5B61",
    x"38F9F9A8",
    x"38F99815",
    x"38F936A9",
    x"38F8D563",
    x"38F87442",
    x"38F81348",
    x"38F7B273",
    x"38F751C4",
    x"38F6F13B",
    x"38F690D8",
    x"38F6309A",
    x"38F5D082",
    x"38F5708F",
    x"38F510C2",
    x"38F4B11A",
    x"38F45198",
    x"38F3F23A",
    x"38F39302",
    x"38F333F0",
    x"38F2D502",
    x"38F27639",
    x"38F21795",
    x"38F1B917",
    x"38F15ABD",
    x"38F0FC88",
    x"38F09E78",
    x"38F0408C",
    x"38EFE2C5",
    x"38EF8523",
    x"38EF27A5",
    x"38EECA4C",
    x"38EE6D17",
    x"38EE1007",
    x"38EDB31A",
    x"38ED5653",
    x"38ECF9AF",
    x"38EC9D30",
    x"38EC40D4",
    x"38EBE49D",
    x"38EB888A",
    x"38EB2C9A",
    x"38EAD0CF",
    x"38EA7527",
    x"38EA19A3",
    x"38E9BE43",
    x"38E96306",
    x"38E907EE",
    x"38E8ACF8",
    x"38E85226",
    x"38E7F778",
    x"38E79CED",
    x"38E74285",
    x"38E6E841",
    x"38E68E20",
    x"38E63422",
    x"38E5DA47",
    x"38E5808F",
    x"38E526FB",
    x"38E4CD89",
    x"38E4743A",
    x"38E41B0E",
    x"38E3C205",
    x"38E3691F",
    x"38E3105B",
    x"38E2B7BA",
    x"38E25F3B",
    x"38E206DF",
    x"38E1AEA6",
    x"38E1568F",
    x"38E0FE9A",
    x"38E0A6C8",
    x"38E04F18",
    x"38DFF78A",
    x"38DFA01F",
    x"38DF48D5",
    x"38DEF1AE",
    x"38DE9AA8",
    x"38DE43C5",
    x"38DDED03",
    x"38DD9664",
    x"38DD3FE6",
    x"38DCE98A",
    x"38DC934F",
    x"38DC3D37",
    x"38DBE73F",
    x"38DB916A",
    x"38DB3BB6",
    x"38DAE623",
    x"38DA90B2",
    x"38DA3B62",
    x"38D9E634",
    x"38D99126",
    x"38D93C3A",
    x"38D8E76F",
    x"38D892C5",
    x"38D83E3D",
    x"38D7E9D5",
    x"38D7958E",
    x"38D74168",
    x"38D6ED63",
    x"38D6997E",
    x"38D645BB",
    x"38D5F218",
    x"38D59E96",
    x"38D54B34",
    x"38D4F7F3",
    x"38D4A4D2",
    x"38D451D2",
    x"38D3FEF2",
    x"38D3AC33",
    x"38D35994",
    x"38D30715",
    x"38D2B4B6",
    x"38D26278",
    x"38D21059",
    x"38D1BE5B",
    x"38D16C7D",
    x"38D11ABE",
    x"38D0C920",
    x"38D077A1",
    x"38D02642",
    x"38CFD503",
    x"38CF83E4",
    x"38CF32E4",
    x"38CEE204",
    x"38CE9143",
    x"38CE40A2",
    x"38CDF021",
    x"38CD9FBF",
    x"38CD4F7C",
    x"38CCFF59",
    x"38CCAF55",
    x"38CC5F70",
    x"38CC0FAA",
    x"38CBC004",
    x"38CB707C",
    x"38CB2114",
    x"38CAD1CA",
    x"38CA82A0",
    x"38CA3394",
    x"38C9E4A7",
    x"38C995D9",
    x"38C9472A",
    x"38C8F89A",
    x"38C8AA28",
    x"38C85BD5",
    x"38C80DA0",
    x"38C7BF8A",
    x"38C77193",
    x"38C723B9",
    x"38C6D5FF",
    x"38C68862",
    x"38C63AE4",
    x"38C5ED84",
    x"38C5A043",
    x"38C5531F",
    x"38C5061A",
    x"38C4B932",
    x"38C46C69",
    x"38C41FBE",
    x"38C3D330",
    x"38C386C1",
    x"38C33A6F",
    x"38C2EE3B",
    x"38C2A225",
    x"38C2562C",
    x"38C20A51",
    x"38C1BE94",
    x"38C172F4",
    x"38C12772",
    x"38C0DC0E",
    x"38C090C6",
    x"38C0459C",
    x"38BFFA90",
    x"38BFAFA1",
    x"38BF64CF",
    x"38BF1A1A",
    x"38BECF82",
    x"38BE8508",
    x"38BE3AAA",
    x"38BDF06A",
    x"38BDA647",
    x"38BD5C40",
    x"38BD1256",
    x"38BCC88A",
    x"38BC7EDA",
    x"38BC3547",
    x"38BBEBD0",
    x"38BBA276",
    x"38BB5939",
    x"38BB1019",
    x"38BAC715",
    x"38BA7E2D",
    x"38BA3562",
    x"38B9ECB3",
    x"38B9A421",
    x"38B95BAB",
    x"38B91351",
    x"38B8CB14",
    x"38B882F3",
    x"38B83AEE",
    x"38B7F305",
    x"38B7AB38",
    x"38B76387",
    x"38B71BF2",
    x"38B6D479",
    x"38B68D1C",
    x"38B645DB",
    x"38B5FEB5",
    x"38B5B7AC",
    x"38B570BE",
    x"38B529EC",
    x"38B4E335",
    x"38B49C9A",
    x"38B4561B",
    x"38B40FB7",
    x"38B3C96F",
    x"38B38342",
    x"38B33D30",
    x"38B2F73A",
    x"38B2B15F",
    x"38B26B9F",
    x"38B225FB",
    x"38B1E071",
    x"38B19B03",
    x"38B155B0",
    x"38B11078",
    x"38B0CB5B",
    x"38B0865A",
    x"38B04173",
    x"38AFFCA6",
    x"38AFB7F5",
    x"38AF735F",
    x"38AF2EE3",
    x"38AEEA82",
    x"38AEA63C",
    x"38AE6210",
    x"38AE1DFF",
    x"38ADDA09",
    x"38AD962D",
    x"38AD526B",
    x"38AD0EC4",
    x"38ACCB38",
    x"38AC87C6",
    x"38AC446E",
    x"38AC0130",
    x"38ABBE0D",
    x"38AB7B04",
    x"38AB3815",
    x"38AAF540",
    x"38AAB285",
    x"38AA6FE4",
    x"38AA2D5E",
    x"38A9EAF1",
    x"38A9A89E",
    x"38A96665",
    x"38A92446",
    x"38A8E241",
    x"38A8A055",
    x"38A85E83",
    x"38A81CCB",
    x"38A7DB2D",
    x"38A799A8",
    x"38A7583D",
    x"38A716EB",
    x"38A6D5B3",
    x"38A69494",
    x"38A6538F",
    x"38A612A3",
    x"38A5D1D0",
    x"38A59117",
    x"38A55077",
    x"38A50FF0",
    x"38A4CF83",
    x"38A48F2E",
    x"38A44EF3",
    x"38A40ED0",
    x"38A3CEC7",
    x"38A38ED7",
    x"38A34EFF",
    x"38A30F41",
    x"38A2CF9C",
    x"38A2900F",
    x"38A2509B",
    x"38A21140",
    x"38A1D1FD",
    x"38A192D4",
    x"38A153C3",
    x"38A114CA",
    x"38A0D5EB",
    x"38A09723",
    x"38A05874",
    x"38A019DE",
    x"389FDB60",
    x"389F9CFB",
    x"389F5EAE",
    x"389F2079",
    x"389EE25C",
    x"389EA458",
    x"389E666C",
    x"389E2898",
    x"389DEADC",
    x"389DAD38",
    x"389D6FAD",
    x"389D3239",
    x"389CF4DD",
    x"389CB79A",
    x"389C7A6E",
    x"389C3D5A",
    x"389C005E",
    x"389BC37A",
    x"389B86AD",
    x"389B49F9",
    x"389B0D5C",
    x"389AD0D6",
    x"389A9468",
    x"389A5812",
    x"389A1BD4",
    x"3899DFAC",
    x"3899A39D",
    x"389967A5",
    x"38992BC4",
    x"3898EFFA",
    x"3898B448",
    x"389878AE",
    x"38983D2A",
    x"389801BE",
    x"3897C669",
    x"38978B2B",
    x"38975004",
    x"389714F4",
    x"3896D9FC",
    x"38969F1A",
    x"3896644F",
    x"3896299B",
    x"3895EEFF",
    x"3895B479",
    x"38957A0A",
    x"38953FB1",
    x"38950570",
    x"3894CB45",
    x"38949131",
    x"38945734",
    x"38941D4D",
    x"3893E37D",
    x"3893A9C3",
    x"38937020",
    x"38933694",
    x"3892FD1E",
    x"3892C3BE",
    x"38928A75",
    x"38925142",
    x"38921825",
    x"3891DF1F",
    x"3891A62F",
    x"38916D55",
    x"38913491",
    x"3890FBE4",
    x"3890C34D",
    x"38908ACB",
    x"38905260",
    x"38901A0B",
    x"388FE1CC",
    x"388FA9A3",
    x"388F718F",
    x"388F3992",
    x"388F01AA",
    x"388EC9D8",
    x"388E921D",
    x"388E5A76",
    x"388E22E6",
    x"388DEB6B",
    x"388DB406",
    x"388D7CB6",
    x"388D457C",
    x"388D0E58",
    x"388CD749",
    x"388CA050",
    x"388C696C",
    x"388C329E",
    x"388BFBE4",
    x"388BC541",
    x"388B8EB2",
    x"388B5839",
    x"388B21D5",
    x"388AEB87",
    x"388AB54D",
    x"388A7F29",
    x"388A491A",
    x"388A1320",
    x"3889DD3B",
    x"3889A76B",
    x"388971B0",
    x"38893C0A",
    x"38890679",
    x"3888D0FD",
    x"38889B96",
    x"38886644",
    x"38883106",
    x"3887FBDD",
    x"3887C6C9",
    x"388791CA",
    x"38875CDF",
    x"38872809",
    x"3886F348",
    x"3886BE9B",
    x"38868A03",
    x"38865580",
    x"38862110",
    x"3885ECB6",
    x"3885B86F",
    x"3885843E",
    x"38855020",
    x"38851C17",
    x"3884E822",
    x"3884B442",
    x"38848075",
    x"38844CBD",
    x"38841919",
    x"3883E58A",
    x"3883B20E",
    x"38837EA7",
    x"38834B53",
    x"38831814",
    x"3882E4E8",
    x"3882B1D1",
    x"38827ECD",
    x"38824BDE",
    x"38821902",
    x"3881E63A",
    x"3881B386",
    x"388180E6",
    x"38814E5A",
    x"38811BE1",
    x"3880E97C",
    x"3880B72A",
    x"388084ED",
    x"388052C2",
    x"388020AC",
    x"387FDD52",
    x"387F7973",
    x"387F15BB",
    x"387EB22A",
    x"387E4EC0",
    x"387DEB7C",
    x"387D8860",
    x"387D256A",
    x"387CC29B",
    x"387C5FF2",
    x"387BFD70",
    x"387B9B14",
    x"387B38DE",
    x"387AD6CF",
    x"387A74E7",
    x"387A1324",
    x"3879B188",
    x"38795011",
    x"3878EEC1",
    x"38788D97",
    x"38782C92",
    x"3877CBB4",
    x"38776AFB",
    x"38770A68",
    x"3876A9FB",
    x"387649B3",
    x"3875E991",
    x"38758995",
    x"387529BE",
    x"3874CA0C",
    x"38746A80",
    x"38740B19",
    x"3873ABD7",
    x"38734CBB",
    x"3872EDC3",
    x"38728EF1",
    x"38723044",
    x"3871D1BB",
    x"38717358",
    x"38711519",
    x"3870B6FF",
    x"3870590A",
    x"386FFB3A",
    x"386F9D8E",
    x"386F4007",
    x"386EE2A4",
    x"386E8566",
    x"386E284C",
    x"386DCB56",
    x"386D6E85",
    x"386D11D8",
    x"386CB54F",
    x"386C58EA",
    x"386BFCA9",
    x"386BA08D",
    x"386B4494",
    x"386AE8BF",
    x"386A8D0E",
    x"386A3181",
    x"3869D617",
    x"38697AD2",
    x"38691FAF",
    x"3868C4B1",
    x"386869D6",
    x"38680F1E",
    x"3867B48A",
    x"38675A19",
    x"3866FFCB",
    x"3866A5A1",
    x"38664B9A",
    x"3865F1B6",
    x"386597F5",
    x"38653E57",
    x"3864E4DC",
    x"38648B85",
    x"3864324F",
    x"3863D93D",
    x"3863804E",
    x"38632781",
    x"3862CED7",
    x"3862764F",
    x"38621DEA",
    x"3861C5A8",
    x"38616D88",
    x"3861158A",
    x"3860BDAF",
    x"386065F6",
    x"38600E5F",
    x"385FB6EB",
    x"385F5F99",
    x"385F0868",
    x"385EB15A",
    x"385E5A6E",
    x"385E03A3",
    x"385DACFB",
    x"385D5674",
    x"385D000F",
    x"385CA9CC",
    x"385C53AB",
    x"385BFDAB",
    x"385BA7CC",
    x"385B5210",
    x"385AFC74",
    x"385AA6FA",
    x"385A51A2",
    x"3859FC6B",
    x"3859A755",
    x"38595260",
    x"3858FD8C",
    x"3858A8DA",
    x"38585448",
    x"3857FFD8",
    x"3857AB88",
    x"3857575A",
    x"3857034C",
    x"3856AF5F",
    x"38565B93",
    x"385607E8",
    x"3855B45D",
    x"385560F3",
    x"38550DA9",
    x"3854BA80",
    x"38546777",
    x"3854148F",
    x"3853C1C7",
    x"38536F20",
    x"38531C98",
    x"3852CA31",
    x"385277EB",
    x"385225C4",
    x"3851D3BD",
    x"385181D6",
    x"38513010",
    x"3850DE69",
    x"38508CE2",
    x"38503B7B",
    x"384FEA33",
    x"384F990C",
    x"384F4804",
    x"384EF71B",
    x"384EA653",
    x"384E55A9",
    x"384E0520",
    x"384DB4B5",
    x"384D646B",
    x"384D143F",
    x"384CC433",
    x"384C7446",
    x"384C2478",
    x"384BD4C9",
    x"384B853A",
    x"384B35C9",
    x"384AE678",
    x"384A9745",
    x"384A4831",
    x"3849F93D",
    x"3849AA67",
    x"38495BAF",
    x"38490D17",
    x"3848BE9D",
    x"38487042",
    x"38482205",
    x"3847D3E7",
    x"384785E8",
    x"38473807",
    x"3846EA44",
    x"38469CA0",
    x"38464F1A",
    x"384601B2",
    x"3845B468",
    x"3845673D",
    x"38451A30",
    x"3844CD41",
    x"3844806F",
    x"384433BC",
    x"3843E727",
    x"38439AB0",
    x"38434E56",
    x"3843021A",
    x"3842B5FC",
    x"384269FC",
    x"38421E1A",
    x"3841D255",
    x"384186AD",
    x"38413B23",
    x"3840EFB7",
    x"3840A468",
    x"38405937",
    x"38400E22",
    x"383FC32C",
    x"383F7852",
    x"383F2D95",
    x"383EE2F6",
    x"383E9874",
    x"383E4E0F",
    x"383E03C7",
    x"383DB99C",
    x"383D6F8E",
    x"383D259D",
    x"383CDBC9",
    x"383C9211",
    x"383C4877",
    x"383BFEF9",
    x"383BB597",
    x"383B6C53",
    x"383B232B",
    x"383ADA1F",
    x"383A9130",
    x"383A485E",
    x"3839FFA8",
    x"3839B70E",
    x"38396E91",
    x"38392630",
    x"3838DDEB",
    x"383895C2",
    x"38384DB6",
    x"383805C6",
    x"3837BDF1",
    x"38377639",
    x"38372E9D",
    x"3836E71D",
    x"38369FB8",
    x"38365870",
    x"38361143",
    x"3835CA32",
    x"3835833D",
    x"38353C64",
    x"3834F5A6",
    x"3834AF04",
    x"3834687D",
    x"38342212",
    x"3833DBC3",
    x"3833958F",
    x"38334F76",
    x"38330979",
    x"3832C397",
    x"38327DD0",
    x"38323824",
    x"3831F294",
    x"3831AD1F",
    x"383167C5",
    x"38312286",
    x"3830DD62",
    x"38309859",
    x"3830536B",
    x"38300E97",
    x"382FC9DF",
    x"382F8542",
    x"382F40BF",
    x"382EFC57",
    x"382EB80A",
    x"382E73D7",
    x"382E2FBF",
    x"382DEBC2",
    x"382DA7DF",
    x"382D6417",
    x"382D2069",
    x"382CDCD6",
    x"382C995C",
    x"382C55FE",
    x"382C12B9",
    x"382BCF8F",
    x"382B8C7F",
    x"382B4989",
    x"382B06AE",
    x"382AC3EC",
    x"382A8145",
    x"382A3EB7",
    x"3829FC44",
    x"3829B9EA",
    x"382977AA",
    x"38293584",
    x"3828F378",
    x"3828B186",
    x"38286FAE",
    x"38282DEF",
    x"3827EC4A",
    x"3827AABE",
    x"3827694C",
    x"382727F4",
    x"3826E6B5",
    x"3826A590",
    x"38266484",
    x"38262391",
    x"3825E2B8",
    x"3825A1F8",
    x"38256151",
    x"382520C4",
    x"3824E050",
    x"38249FF5",
    x"38245FB3",
    x"38241F8A",
    x"3823DF7A",
    x"38239F83",
    x"38235FA6",
    x"38231FE1",
    x"3822E035",
    x"3822A0A2",
    x"38226127",
    x"382221C6",
    x"3821E27D",
    x"3821A34D",
    x"38216435",
    x"38212536",
    x"3820E650",
    x"3820A782",
    x"382068CD",
    x"38202A31",
    x"381FEBAC",
    x"381FAD40",
    x"381F6EED",
    x"381F30B2",
    x"381EF28F",
    x"381EB484",
    x"381E7692",
    x"381E38B8",
    x"381DFAF5",
    x"381DBD4C",
    x"381D7FBA",
    x"381D4240",
    x"381D04DE",
    x"381CC794",
    x"381C8A62",
    x"381C4D48",
    x"381C1045",
    x"381BD35B",
    x"381B9688",
    x"381B59CD",
    x"381B1D2A",
    x"381AE09F",
    x"381AA42B",
    x"381A67CE",
    x"381A2B8A",
    x"3819EF5C",
    x"3819B347",
    x"38197748",
    x"38193B61",
    x"3818FF92",
    x"3818C3DA",
    x"38188839",
    x"38184CAF",
    x"3818113D",
    x"3817D5E2",
    x"38179A9E",
    x"38175F71",
    x"3817245B",
    x"3816E95D",
    x"3816AE75",
    x"381673A4",
    x"381638EB",
    x"3815FE48",
    x"3815C3BC",
    x"38158947",
    x"38154EE9",
    x"381514A1",
    x"3814DA70",
    x"3814A057",
    x"38146653",
    x"38142C67",
    x"3813F291",
    x"3813B8D1",
    x"38137F28",
    x"38134596",
    x"38130C1A",
    x"3812D2B4",
    x"38129965",
    x"3812602C",
    x"3812270A",
    x"3811EDFE",
    x"3811B508",
    x"38117C28",
    x"3811435F",
    x"38110AAC",
    x"3810D20F",
    x"38109988",
    x"38106117",
    x"381028BC",
    x"380FF077",
    x"380FB848",
    x"380F802F",
    x"380F482C",
    x"380F103F",
    x"380ED867",
    x"380EA0A5",
    x"380E68FA",
    x"380E3163",
    x"380DF9E3",
    x"380DC278",
    x"380D8B23",
    x"380D53E3",
    x"380D1CB9",
    x"380CE5A5",
    x"380CAEA6",
    x"380C77BD",
    x"380C40E9",
    x"380C0A2A",
    x"380BD381",
    x"380B9CED",
    x"380B666E",
    x"380B3005",
    x"380AF9B0",
    x"380AC371",
    x"380A8D48",
    x"380A5733",
    x"380A2134",
    x"3809EB49",
    x"3809B574",
    x"38097FB3",
    x"38094A08",
    x"38091472",
    x"3808DEF0",
    x"3808A983",
    x"3808742C",
    x"38083EE9",
    x"380809BA",
    x"3807D4A1",
    x"38079F9C",
    x"38076AAC",
    x"380735D1",
    x"3807010A",
    x"3806CC58",
    x"380697BB",
    x"38066332",
    x"38062EBD",
    x"3805FA5D",
    x"3805C611",
    x"380591DA",
    x"38055DB7",
    x"380529A9",
    x"3804F5AF",
    x"3804C1C9",
    x"38048DF8",
    x"38045A3A",
    x"38042691",
    x"3803F2FC",
    x"3803BF7B",
    x"38038C0E",
    x"380358B6",
    x"38032571",
    x"3802F240",
    x"3802BF24",
    x"38028C1B",
    x"38025926",
    x"38022645",
    x"3801F378",
    x"3801C0BF",
    x"38018E1A",
    x"38015B88",
    x"3801290A",
    x"3800F6A0",
    x"3800C44A",
    x"38009207",
    x"38005FD8",
    x"38002DBC",
    x"37FFF768",
    x"37FF937F",
    x"37FF2FBC",
    x"37FECC21",
    x"37FE68AD",
    x"37FE055F",
    x"37FDA239",
    x"37FD3F39",
    x"37FCDC5F",
    x"37FC79AC",
    x"37FC1720",
    x"37FBB4BA",
    x"37FB527B",
    x"37FAF062",
    x"37FA8E6F",
    x"37FA2CA3",
    x"37F9CAFC",
    x"37F9697C",
    x"37F90822",
    x"37F8A6EE",
    x"37F845DF",
    x"37F7E4F7",
    x"37F78435",
    x"37F72398",
    x"37F6C321",
    x"37F662CF",
    x"37F602A3",
    x"37F5A29D",
    x"37F542BC",
    x"37F4E301",
    x"37F4836B",
    x"37F423FA",
    x"37F3C4AF",
    x"37F36589",
    x"37F30688",
    x"37F2A7AC",
    x"37F248F5",
    x"37F1EA63",
    x"37F18BF5",
    x"37F12DAD",
    x"37F0CF8A",
    x"37F0718B",
    x"37F013B1",
    x"37EFB5FC",
    x"37EF586B",
    x"37EEFAFF",
    x"37EE9DB7",
    x"37EE4093",
    x"37EDE394",
    x"37ED86B9",
    x"37ED2A03",
    x"37ECCD71",
    x"37EC7102",
    x"37EC14B8",
    x"37EBB892",
    x"37EB5C90",
    x"37EB00B2",
    x"37EAA4F8",
    x"37EA4961",
    x"37E9EDEE",
    x"37E9929F",
    x"37E93774",
    x"37E8DC6C",
    x"37E88187",
    x"37E826C7",
    x"37E7CC29",
    x"37E771AF",
    x"37E71758",
    x"37E6BD25",
    x"37E66315",
    x"37E60927",
    x"37E5AF5D",
    x"37E555B6",
    x"37E4FC32",
    x"37E4A2D1",
    x"37E44993",
    x"37E3F078",
    x"37E3977F",
    x"37E33EA9",
    x"37E2E5F6",
    x"37E28D66",
    x"37E234F8",
    x"37E1DCAC",
    x"37E18483",
    x"37E12C7D",
    x"37E0D499",
    x"37E07CD7",
    x"37E02537",
    x"37DFCDBA",
    x"37DF765E",
    x"37DF1F25",
    x"37DEC80E",
    x"37DE7119",
    x"37DE1A46",
    x"37DDC394",
    x"37DD6D05",
    x"37DD1697",
    x"37DCC04B",
    x"37DC6A21",
    x"37DC1418",
    x"37DBBE31",
    x"37DB686C",
    x"37DB12C8",
    x"37DABD45",
    x"37DA67E4",
    x"37DA12A4",
    x"37D9BD85",
    x"37D96888",
    x"37D913AB",
    x"37D8BEF0",
    x"37D86A56",
    x"37D815DD",
    x"37D7C185",
    x"37D76D4E",
    x"37D71938",
    x"37D6C542",
    x"37D6716E",
    x"37D61DBA",
    x"37D5CA26",
    x"37D576B4",
    x"37D52362",
    x"37D4D030",
    x"37D47D1F",
    x"37D42A2E",
    x"37D3D75E",
    x"37D384AE",
    x"37D3321E",
    x"37D2DFAF",
    x"37D28D5F",
    x"37D23B30",
    x"37D1E921",
    x"37D19732",
    x"37D14563",
    x"37D0F3B4",
    x"37D0A225",
    x"37D050B5",
    x"37CFFF66",
    x"37CFAE36",
    x"37CF5D26",
    x"37CF0C35",
    x"37CEBB64",
    x"37CE6AB3",
    x"37CE1A21",
    x"37CDC9AE",
    x"37CD795B",
    x"37CD2927",
    x"37CCD913",
    x"37CC891E",
    x"37CC3948",
    x"37CBE991",
    x"37CB99F9",
    x"37CB4A81",
    x"37CAFB27",
    x"37CAABEC",
    x"37CA5CD1",
    x"37CA0DD4",
    x"37C9BEF6",
    x"37C97037",
    x"37C92196",
    x"37C8D314",
    x"37C884B1",
    x"37C8366D",
    x"37C7E847",
    x"37C79A3F",
    x"37C74C56",
    x"37C6FE8C",
    x"37C6B0DF",
    x"37C66351",
    x"37C615E2",
    x"37C5C890",
    x"37C57B5D",
    x"37C52E48",
    x"37C4E151",
    x"37C49478",
    x"37C447BD",
    x"37C3FB20",
    x"37C3AEA1",
    x"37C3623F",
    x"37C315FC",
    x"37C2C9D6",
    x"37C27DCE",
    x"37C231E4",
    x"37C1E617",
    x"37C19A68",
    x"37C14ED6",
    x"37C10362",
    x"37C0B80C",
    x"37C06CD3",
    x"37C021B7",
    x"37BFD6B8",
    x"37BF8BD7",
    x"37BF4113",
    x"37BEF66C",
    x"37BEABE2",
    x"37BE6176",
    x"37BE1726",
    x"37BDCCF4",
    x"37BD82DE",
    x"37BD38E6",
    x"37BCEF0A",
    x"37BCA54B",
    x"37BC5BA9",
    x"37BC1223",
    x"37BBC8BA",
    x"37BB7F6E",
    x"37BB363F",
    x"37BAED2C",
    x"37BAA436",
    x"37BA5B5C",
    x"37BA129E",
    x"37B9C9FD",
    x"37B98178",
    x"37B93910",
    x"37B8F0C4",
    x"37B8A894",
    x"37B86080",
    x"37B81888",
    x"37B7D0AD",
    x"37B788ED",
    x"37B7414A",
    x"37B6F9C2",
    x"37B6B257",
    x"37B66B07",
    x"37B623D3",
    x"37B5DCBB",
    x"37B595BF",
    x"37B54EDE",
    x"37B50819",
    x"37B4C170",
    x"37B47AE2",
    x"37B43470",
    x"37B3EE19",
    x"37B3A7DE",
    x"37B361BE",
    x"37B31BB9",
    x"37B2D5D0",
    x"37B29002",
    x"37B24A50",
    x"37B204B8",
    x"37B1BF3C",
    x"37B179DB",
    x"37B13495",
    x"37B0EF6A",
    x"37B0AA5A",
    x"37B06564",
    x"37B0208A",
    x"37AFDBCB",
    x"37AF9727",
    x"37AF529D",
    x"37AF0E2E",
    x"37AEC9DA",
    x"37AE85A0",
    x"37AE4181",
    x"37ADFD7D",
    x"37ADB993",
    x"37AD75C4",
    x"37AD320F",
    x"37ACEE75",
    x"37ACAAF5",
    x"37AC678F",
    x"37AC2444",
    x"37ABE113",
    x"37AB9DFC",
    x"37AB5B00",
    x"37AB181D",
    x"37AAD555",
    x"37AA92A7",
    x"37AA5012",
    x"37AA0D98",
    x"37A9CB38",
    x"37A988F1",
    x"37A946C5",
    x"37A904B2",
    x"37A8C2B9",
    x"37A880DA",
    x"37A83F14",
    x"37A7FD68",
    x"37A7BBD6",
    x"37A77A5E",
    x"37A738FF",
    x"37A6F7B9",
    x"37A6B68D",
    x"37A6757A",
    x"37A63481",
    x"37A5F3A1",
    x"37A5B2DB",
    x"37A5722E",
    x"37A5319A",
    x"37A4F11F",
    x"37A4B0BD",
    x"37A47075",
    x"37A43045",
    x"37A3F02F",
    x"37A3B032",
    x"37A3704D",
    x"37A33082",
    x"37A2F0D0",
    x"37A2B136",
    x"37A271B5",
    x"37A2324D",
    x"37A1F2FE",
    x"37A1B3C7",
    x"37A174A9",
    x"37A135A4",
    x"37A0F6B7",
    x"37A0B7E3",
    x"37A07928",
    x"37A03A85",
    x"379FFBFA",
    x"379FBD88",
    x"379F7F2E",
    x"379F40EC",
    x"379F02C3",
    x"379EC4B2",
    x"379E86BA",
    x"379E48D9",
    x"379E0B11",
    x"379DCD60",
    x"379D8FC8",
    x"379D5248",
    x"379D14E0",
    x"379CD790",
    x"379C9A57",
    x"379C5D37",
    x"379C202F",
    x"379BE33E",
    x"379BA665",
    x"379B69A4",
    x"379B2CFA",
    x"379AF069",
    x"379AB3EF",
    x"379A778C",
    x"379A3B41",
    x"3799FF0E",
    x"3799C2F2",
    x"379986EE",
    x"37994B01",
    x"37990F2B",
    x"3798D36D",
    x"379897C6",
    x"37985C36",
    x"379820BE",
    x"3797E55D",
    x"3797AA12",
    x"37976EE0",
    x"379733C4",
    x"3796F8BF",
    x"3796BDD2",
    x"379682FB",
    x"3796483B",
    x"37960D92",
    x"3795D301",
    x"37959886",
    x"37955E21",
    x"379523D4",
    x"3794E99D",
    x"3794AF7D",
    x"37947574",
    x"37943B82",
    x"379401A6",
    x"3793C7E0",
    x"37938E32",
    x"37935499",
    x"37931B18",
    x"3792E1AC",
    x"3792A857",
    x"37926F19",
    x"379235F0",
    x"3791FCDE",
    x"3791C3E3",
    x"37918AFD",
    x"3791522E",
    x"37911975",
    x"3790E0D2",
    x"3790A846",
    x"37906FCF",
    x"3790376E",
    x"378FFF24",
    x"378FC6EF",
    x"378F8ED0",
    x"378F56C7",
    x"378F1ED4",
    x"378EE6F7",
    x"378EAF30",
    x"378E777E",
    x"378E3FE2",
    x"378E085C",
    x"378DD0EC",
    x"378D9991",
    x"378D624C",
    x"378D2B1C",
    x"378CF402",
    x"378CBCFE",
    x"378C860F",
    x"378C4F35",
    x"378C1871",
    x"378BE1C2",
    x"378BAB28",
    x"378B74A4",
    x"378B3E35",
    x"378B07DC",
    x"378AD197",
    x"378A9B68",
    x"378A654E",
    x"378A2F49",
    x"3789F959",
    x"3789C37E",
    x"37898DB8",
    x"37895807",
    x"3789226B",
    x"3788ECE4",
    x"3788B772",
    x"37888215",
    x"37884CCC",
    x"37881799",
    x"3787E27A",
    x"3787AD70",
    x"3787787A",
    x"3787439A",
    x"37870ECE",
    x"3786DA16",
    x"3786A573",
    x"378670E5",
    x"37863C6B",
    x"37860806",
    x"3785D3B5",
    x"37859F78",
    x"37856B50",
    x"3785373C",
    x"3785033D",
    x"3784CF52",
    x"37849B7B",
    x"378467B8",
    x"3784340A",
    x"37840070",
    x"3783CCEA",
    x"37839978",
    x"3783661A",
    x"378332D0",
    x"3782FF9A",
    x"3782CC78",
    x"3782996A",
    x"37826670",
    x"3782338A",
    x"378200B8",
    x"3781CDFA",
    x"37819B4F",
    x"378168B8",
    x"37813635",
    x"378103C6",
    x"3780D16A",
    x"37809F22",
    x"37806CEE",
    x"37803ACD",
    x"378008C0",
    x"377FAD8D",
    x"377F49C0",
    x"377EE61B",
    x"377E829D",
    x"377E1F45",
    x"377DBC14",
    x"377D590A",
    x"377CF627",
    x"377C936A",
    x"377C30D3",
    x"377BCE64",
    x"377B6C1A",
    x"377B09F7",
    x"377AA7FA",
    x"377A4624",
    x"3779E474",
    x"377982E9",
    x"37792185",
    x"3778C047",
    x"37785F2F",
    x"3777FE3D",
    x"37779D70",
    x"37773CCA",
    x"3776DC49",
    x"37767BEE",
    x"37761BB8",
    x"3775BBA8",
    x"37755BBD",
    x"3774FBF8",
    x"37749C59",
    x"37743CDE",
    x"3773DD89",
    x"37737E59",
    x"37731F4E",
    x"3772C069",
    x"377261A8",
    x"3772030C",
    x"3771A496",
    x"37714644",
    x"3770E817",
    x"37708A0E",
    x"37702C2B",
    x"376FCE6C",
    x"376F70D1",
    x"376F135C",
    x"376EB60A",
    x"376E58DD",
    x"376DFBD5",
    x"376D9EF1",
    x"376D4231",
    x"376CE595",
    x"376C891D",
    x"376C2CCA",
    x"376BD09A",
    x"376B748F",
    x"376B18A7",
    x"376ABCE4",
    x"376A6144",
    x"376A05C8",
    x"3769AA6F",
    x"37694F3A",
    x"3768F429",
    x"3768993C",
    x"37683E71",
    x"3767E3CB",
    x"37678947",
    x"37672EE8",
    x"3766D4AB",
    x"37667A91",
    x"3766209B",
    x"3765C6C8",
    x"37656D18",
    x"3765138B",
    x"3764BA20",
    x"376460D9",
    x"376407B5",
    x"3763AEB3",
    x"376355D4",
    x"3762FD18",
    x"3762A47F",
    x"37624C08",
    x"3761F3B3",
    x"37619B81",
    x"37614372",
    x"3760EB84",
    x"376093BA",
    x"37603C11",
    x"375FE48B",
    x"375F8D26",
    x"375F35E4",
    x"375EDEC4",
    x"375E87C6",
    x"375E30EA",
    x"375DDA30",
    x"375D8398",
    x"375D2D21",
    x"375CD6CC",
    x"375C8099",
    x"375C2A88",
    x"375BD498",
    x"375B7ECA",
    x"375B291D",
    x"375AD392",
    x"375A7E28",
    x"375A28DF",
    x"3759D3B8",
    x"37597EB2",
    x"375929CD",
    x"3758D509",
    x"37588066",
    x"37582BE5",
    x"3757D784",
    x"37578344",
    x"37572F26",
    x"3756DB27",
    x"3756874A",
    x"3756338E",
    x"3755DFF2",
    x"37558C77",
    x"3755391C",
    x"3754E5E2",
    x"375492C9",
    x"37543FCF",
    x"3753ECF7",
    x"37539A3E",
    x"375347A6",
    x"3752F52E",
    x"3752A2D7",
    x"3752509F",
    x"3751FE88",
    x"3751AC90",
    x"37515AB9",
    x"37510901",
    x"3750B76A",
    x"375065F2",
    x"3750149A",
    x"374FC362",
    x"374F7249",
    x"374F2151",
    x"374ED077",
    x"374E7FBE",
    x"374E2F24",
    x"374DDEA9",
    x"374D8E4E",
    x"374D3E12",
    x"374CEDF5",
    x"374C9DF8",
    x"374C4E1A",
    x"374BFE5B",
    x"374BAEBB",
    x"374B5F3A",
    x"374B0FD9",
    x"374AC096",
    x"374A7172",
    x"374A226D",
    x"3749D387",
    x"374984C0",
    x"37493617",
    x"3748E78E",
    x"37489923",
    x"37484AD6",
    x"3747FCA8",
    x"3747AE99",
    x"374760A8",
    x"374712D5",
    x"3746C521",
    x"3746778B",
    x"37462A13",
    x"3745DCBA",
    x"37458F7F",
    x"37454262",
    x"3744F563",
    x"3744A882",
    x"37445BBF",
    x"37440F1B",
    x"3743C294",
    x"3743762B",
    x"374329DF",
    x"3742DDB2",
    x"374291A2",
    x"374245B0",
    x"3741F9DC",
    x"3741AE25",
    x"3741628C",
    x"37411710",
    x"3740CBB2",
    x"37408071",
    x"3740354D",
    x"373FEA47",
    x"373F9F5E",
    x"373F5493",
    x"373F09E4",
    x"373EBF53",
    x"373E74DF",
    x"373E2A87",
    x"373DE04D",
    x"373D9630",
    x"373D4C30",
    x"373D024D",
    x"373CB886",
    x"373C6EDD",
    x"373C2550",
    x"373BDBDF",
    x"373B928C",
    x"373B4955",
    x"373B003A",
    x"373AB73D",
    x"373A6E5B",
    x"373A2596",
    x"3739DCEE",
    x"37399462",
    x"37394BF2",
    x"3739039E",
    x"3738BB67",
    x"3738734C",
    x"37382B4D",
    x"3737E36A",
    x"37379BA3",
    x"373753F9",
    x"37370C6A",
    x"3736C4F7",
    x"37367DA0",
    x"37363665",
    x"3735EF45",
    x"3735A842",
    x"3735615A",
    x"37351A8E",
    x"3734D3DD",
    x"37348D48",
    x"373446CF",
    x"37340071",
    x"3733BA2E",
    x"37337407",
    x"37332DFC",
    x"3732E80B",
    x"3732A236",
    x"37325C7D",
    x"373216DE",
    x"3731D15B",
    x"37318BF3",
    x"373146A5",
    x"37310173",
    x"3730BC5C",
    x"37307760",
    x"3730327F",
    x"372FEDB9",
    x"372FA90D",
    x"372F647D",
    x"372F2007",
    x"372EDBAC",
    x"372E976B",
    x"372E5345",
    x"372E0F3A",
    x"372DCB49",
    x"372D8773",
    x"372D43B8",
    x"372D0016",
    x"372CBC8F",
    x"372C7923",
    x"372C35D1",
    x"372BF299",
    x"372BAF7B",
    x"372B6C78",
    x"372B298F",
    x"372AE6BF",
    x"372AA40A",
    x"372A616F",
    x"372A1EEE",
    x"3729DC87",
    x"37299A3A",
    x"37295807",
    x"372915ED",
    x"3728D3ED",
    x"37289207",
    x"3728503B",
    x"37280E89",
    x"3727CCF0",
    x"37278B71",
    x"37274A0B",
    x"372708BF",
    x"3726C78C",
    x"37268673",
    x"37264573",
    x"3726048D",
    x"3725C3BF",
    x"3725830C",
    x"37254271",
    x"372501F0",
    x"3724C188",
    x"37248139",
    x"37244103",
    x"372400E6",
    x"3723C0E2",
    x"372380F7",
    x"37234125",
    x"3723016C",
    x"3722C1CC",
    x"37228245",
    x"372242D6",
    x"37220380",
    x"3721C443",
    x"3721851F",
    x"37214613",
    x"37210720",
    x"3720C846",
    x"37208984",
    x"37204ADA",
    x"37200C49",
    x"371FCDD1",
    x"371F8F71",
    x"371F5129",
    x"371F12F9",
    x"371ED4E2",
    x"371E96E3",
    x"371E58FC",
    x"371E1B2D",
    x"371DDD77",
    x"371D9FD8",
    x"371D6252",
    x"371D24E3",
    x"371CE78D",
    x"371CAA4F",
    x"371C6D28",
    x"371C3019",
    x"371BF322",
    x"371BB643",
    x"371B797C",
    x"371B3CCC",
    x"371B0034",
    x"371AC3B4",
    x"371A874C",
    x"371A4AFB",
    x"371A0EC1",
    x"3719D29F",
    x"37199694",
    x"37195AA1",
    x"37191EC6",
    x"3718E301",
    x"3718A754",
    x"37186BBF",
    x"37183040",
    x"3717F4D9",
    x"3717B989",
    x"37177E50",
    x"3717432E",
    x"37170823",
    x"3716CD30",
    x"37169253",
    x"3716578D",
    x"37161CDF",
    x"3715E247",
    x"3715A7C6",
    x"37156D5C",
    x"37153308",
    x"3714F8CC",
    x"3714BEA6",
    x"37148497",
    x"37144A9E",
    x"371410BD",
    x"3713D6F1",
    x"37139D3D",
    x"3713639E",
    x"37132A17",
    x"3712F0A6",
    x"3712B74B",
    x"37127E06",
    x"371244D8",
    x"37120BC1",
    x"3711D2BF",
    x"371199D4",
    x"371160FF",
    x"37112840",
    x"3710EF97",
    x"3710B705",
    x"37107E88",
    x"37104622",
    x"37100DD2",
    x"370FD597",
    x"370F9D73",
    x"370F6564",
    x"370F2D6C",
    x"370EF589",
    x"370EBDBC",
    x"370E8605",
    x"370E4E63",
    x"370E16D7",
    x"370DDF61",
    x"370DA801",
    x"370D70B6",
    x"370D3981",
    x"370D0261",
    x"370CCB57",
    x"370C9462",
    x"370C5D83",
    x"370C26B9",
    x"370BF005",
    x"370BB966",
    x"370B82DC",
    x"370B4C67",
    x"370B1608",
    x"370ADFBE",
    x"370AA989",
    x"370A736A",
    x"370A3D5F",
    x"370A076A",
    x"3709D189",
    x"37099BBE",
    x"37096608",
    x"37093066",
    x"3708FADA",
    x"3708C562",
    x"37089000",
    x"37085AB2",
    x"37082579",
    x"3707F054",
    x"3707BB45",
    x"3707864A",
    x"37075164",
    x"37071C93",
    x"3706E7D6",
    x"3706B32D",
    x"37067E9A",
    x"37064A1A",
    x"370615B0",
    x"3705E15A",
    x"3705AD18",
    x"370578EA",
    x"370544D1",
    x"370510CC",
    x"3704DCDC",
    x"3704A900",
    x"37047538",
    x"37044184",
    x"37040DE5",
    x"3703DA59",
    x"3703A6E2",
    x"3703737F",
    x"37034030",
    x"37030CF5",
    x"3702D9CE",
    x"3702A6BB",
    x"370273BC",
    x"370240D0",
    x"37020DF9",
    x"3701DB35",
    x"3701A886",
    x"370175EA",
    x"37014362",
    x"370110ED",
    x"3700DE8C",
    x"3700AC3F",
    x"37007A06",
    x"370047E0",
    x"370015CE",
    x"36FFC79E",
    x"36FF63C7",
    x"36FF0018",
    x"36FE9C8F",
    x"36FE392D",
    x"36FDD5F2",
    x"36FD72DE",
    x"36FD0FF1",
    x"36FCAD2A",
    x"36FC4A89",
    x"36FBE80F",
    x"36FB85BC",
    x"36FB238F",
    x"36FAC188",
    x"36FA5FA8",
    x"36F9FDED",
    x"36F99C59",
    x"36F93AEB",
    x"36F8D9A3",
    x"36F87881",
    x"36F81785",
    x"36F7B6AF",
    x"36F755FE",
    x"36F6F574",
    x"36F6950F",
    x"36F634CF",
    x"36F5D4B5",
    x"36F574C1",
    x"36F514F2",
    x"36F4B549",
    x"36F455C4",
    x"36F3F666",
    x"36F3972C",
    x"36F33817",
    x"36F2D928",
    x"36F27A5E",
    x"36F21BB8",
    x"36F1BD38",
    x"36F15EDD",
    x"36F100A6",
    x"36F0A294",
    x"36F044A7",
    x"36EFE6DE",
    x"36EF893B",
    x"36EF2BBB",
    x"36EECE60",
    x"36EE712A",
    x"36EE1418",
    x"36EDB72A",
    x"36ED5A61",
    x"36ECFDBC",
    x"36ECA13B",
    x"36EC44DE",
    x"36EBE8A5",
    x"36EB8C90",
    x"36EB309F",
    x"36EAD4D2",
    x"36EA7929",
    x"36EA1DA3",
    x"36E9C241",
    x"36E96703",
    x"36E90BE9",
    x"36E8B0F2",
    x"36E8561F",
    x"36E7FB6F",
    x"36E7A0E2",
    x"36E74679",
    x"36E6EC33",
    x"36E69211",
    x"36E63811",
    x"36E5DE35",
    x"36E5847B",
    x"36E52AE5",
    x"36E4D172",
    x"36E47822",
    x"36E41EF4",
    x"36E3C5E9",
    x"36E36D01",
    x"36E3143C",
    x"36E2BB9A",
    x"36E2631A",
    x"36E20ABC",
    x"36E1B281",
    x"36E15A69",
    x"36E10273",
    x"36E0AA9F",
    x"36E052ED",
    x"36DFFB5E",
    x"36DFA3F1",
    x"36DF4CA6",
    x"36DEF57D",
    x"36DE9E76",
    x"36DE4791",
    x"36DDF0CE",
    x"36DD9A2D",
    x"36DD43AE",
    x"36DCED50",
    x"36DC9714",
    x"36DC40FA",
    x"36DBEB01",
    x"36DB952A",
    x"36DB3F75",
    x"36DAE9E1",
    x"36DA946E",
    x"36DA3F1D",
    x"36D9E9ED",
    x"36D994DE",
    x"36D93FF1",
    x"36D8EB24",
    x"36D89679",
    x"36D841EF",
    x"36D7ED85",
    x"36D7993D",
    x"36D74516",
    x"36D6F10F",
    x"36D69D29",
    x"36D64964",
    x"36D5F5C0",
    x"36D5A23C",
    x"36D54ED9",
    x"36D4FB97",
    x"36D4A875",
    x"36D45573",
    x"36D40292",
    x"36D3AFD1",
    x"36D35D30",
    x"36D30AB0",
    x"36D2B850",
    x"36D26610",
    x"36D213F0",
    x"36D1C1F0",
    x"36D17011",
    x"36D11E51",
    x"36D0CCB1",
    x"36D07B31",
    x"36D029D1",
    x"36CFD890",
    x"36CF8770",
    x"36CF366E",
    x"36CEE58D",
    x"36CE94CB",
    x"36CE4429",
    x"36CDF3A6",
    x"36CDA342",
    x"36CD52FE",
    x"36CD02DA",
    x"36CCB2D4",
    x"36CC62EE",
    x"36CC1327",
    x"36CBC37F",
    x"36CB73F6",
    x"36CB248C",
    x"36CAD541",
    x"36CA8616",
    x"36CA3709",
    x"36C9E81B",
    x"36C9994B",
    x"36C94A9B",
    x"36C8FC09",
    x"36C8AD96",
    x"36C85F41",
    x"36C8110B",
    x"36C7C2F4",
    x"36C774FB",
    x"36C72721",
    x"36C6D965",
    x"36C68BC7",
    x"36C63E47",
    x"36C5F0E6",
    x"36C5A3A3",
    x"36C5567E",
    x"36C50978",
    x"36C4BC8F",
    x"36C46FC4",
    x"36C42318",
    x"36C3D689",
    x"36C38A18",
    x"36C33DC5",
    x"36C2F190",
    x"36C2A578",
    x"36C2597E",
    x"36C20DA2",
    x"36C1C1E4",
    x"36C17643",
    x"36C12ABF",
    x"36C0DF59",
    x"36C09411",
    x"36C048E6",
    x"36BFFDD8",
    x"36BFB2E7",
    x"36BF6814",
    x"36BF1D5E",
    x"36BED2C5",
    x"36BE8849",
    x"36BE3DEB",
    x"36BDF3A9",
    x"36BDA984",
    x"36BD5F7C",
    x"36BD1592",
    x"36BCCBC4",
    x"36BC8212",
    x"36BC387E",
    x"36BBEF06",
    x"36BBA5AB",
    x"36BB5C6D",
    x"36BB134B",
    x"36BACA46",
    x"36BA815D",
    x"36BA3891",
    x"36B9EFE1",
    x"36B9A74D",
    x"36B95ED6",
    x"36B9167B",
    x"36B8CE3C",
    x"36B8861A",
    x"36B83E14",
    x"36B7F629",
    x"36B7AE5B",
    x"36B766A9",
    x"36B71F13",
    x"36B6D799",
    x"36B6903B",
    x"36B648F8",
    x"36B601D2",
    x"36B5BAC7",
    x"36B573D8",
    x"36B52D04",
    x"36B4E64D",
    x"36B49FB0",
    x"36B45930",
    x"36B412CB",
    x"36B3CC81",
    x"36B38653",
    x"36B34040",
    x"36B2FA49",
    x"36B2B46D",
    x"36B26EAC",
    x"36B22906",
    x"36B1E37C",
    x"36B19E0C",
    x"36B158B8",
    x"36B1137F",
    x"36B0CE61",
    x"36B0895E",
    x"36B04476",
    x"36AFFFA8",
    x"36AFBAF6",
    x"36AF765E",
    x"36AF31E1",
    x"36AEED7F",
    x"36AEA938",
    x"36AE650B",
    x"36AE20F9",
    x"36ADDD01",
    x"36AD9924",
    x"36AD5562",
    x"36AD11B9",
    x"36ACCE2C",
    x"36AC8AB8",
    x"36AC475F",
    x"36AC0421",
    x"36ABC0FC",
    x"36AB7DF2",
    x"36AB3B02",
    x"36AAF82C",
    x"36AAB570",
    x"36AA72CE",
    x"36AA3046",
    x"36A9EDD8",
    x"36A9AB84",
    x"36A9694A",
    x"36A9272A",
    x"36A8E524",
    x"36A8A337",
    x"36A86164",
    x"36A81FAB",
    x"36A7DE0B",
    x"36A79C85",
    x"36A75B19",
    x"36A719C6",
    x"36A6D88D",
    x"36A6976D",
    x"36A65667",
    x"36A61579",
    x"36A5D4A6",
    x"36A593EB",
    x"36A5534A",
    x"36A512C2",
    x"36A4D254",
    x"36A491FE",
    x"36A451C1",
    x"36A4119E",
    x"36A3D194",
    x"36A391A2",
    x"36A351CA",
    x"36A3120A",
    x"36A2D264",
    x"36A292D6",
    x"36A25361",
    x"36A21405",
    x"36A1D4C1",
    x"36A19597",
    x"36A15685",
    x"36A1178B",
    x"36A0D8AA",
    x"36A099E2",
    x"36A05B32",
    x"36A01C9A",
    x"369FDE1C",
    x"369F9FB5",
    x"369F6167",
    x"369F2331",
    x"369EE513",
    x"369EA70E",
    x"369E6921",
    x"369E2B4C",
    x"369DED8F",
    x"369DAFEA",
    x"369D725D",
    x"369D34E9",
    x"369CF78C",
    x"369CBA47",
    x"369C7D1B",
    x"369C4006",
    x"369C0308",
    x"369BC623",
    x"369B8956",
    x"369B4CA0",
    x"369B1002",
    x"369AD37B",
    x"369A970D",
    x"369A5AB5",
    x"369A1E76",
    x"3699E24E",
    x"3699A63D",
    x"36996A44",
    x"36992E62",
    x"3698F297",
    x"3698B6E4",
    x"36987B49",
    x"36983FC4",
    x"36980457",
    x"3697C901",
    x"36978DC2",
    x"3697529A",
    x"36971789",
    x"3696DC8F",
    x"3696A1AD",
    x"369666E1",
    x"36962C2C",
    x"3695F18F",
    x"3695B708",
    x"36957C98",
    x"3695423E",
    x"369507FC",
    x"3694CDD0",
    x"369493BB",
    x"369459BD",
    x"36941FD5",
    x"3693E604",
    x"3693AC49",
    x"369372A5",
    x"36933918",
    x"3692FFA1",
    x"3692C640",
    x"36928CF6",
    x"369253C2",
    x"36921AA4",
    x"3691E19D",
    x"3691A8AC",
    x"36916FD1",
    x"3691370D",
    x"3690FE5E",
    x"3690C5C6",
    x"36908D44",
    x"369054D7",
    x"36901C81",
    x"368FE441",
    x"368FAC17",
    x"368F7403",
    x"368F3C04",
    x"368F041C",
    x"368ECC49",
    x"368E948C",
    x"368E5CE5",
    x"368E2554",
    x"368DEDD8",
    x"368DB672",
    x"368D7F21",
    x"368D47E6",
    x"368D10C1",
    x"368CD9B1",
    x"368CA2B7",
    x"368C6BD2",
    x"368C3503",
    x"368BFE49",
    x"368BC7A4",
    x"368B9115",
    x"368B5A9B",
    x"368B2436",
    x"368AEDE6",
    x"368AB7AC",
    x"368A8187",
    x"368A4B77",
    x"368A157C",
    x"3689DF96",
    x"3689A9C5",
    x"3689740A",
    x"36893E63",
    x"368908D1",
    x"3688D354",
    x"36889DEC",
    x"36886898",
    x"3688335A",
    x"3687FE30",
    x"3687C91B",
    x"3687941B",
    x"36875F30",
    x"36872A59",
    x"3686F597",
    x"3686C0E9",
    x"36868C50",
    x"368657CB",
    x"3686235B",
    x"3685EF00",
    x"3685BAB8",
    x"36858686",
    x"36855267",
    x"36851E5D",
    x"3684EA68",
    x"3684B686",
    x"368482B9",
    x"36844F00",
    x"36841B5B",
    x"3683E7CB",
    x"3683B44E",
    x"368380E6",
    x"36834D91",
    x"36831A51",
    x"3682E725",
    x"3682B40D",
    x"36828108",
    x"36824E18",
    x"36821B3B",
    x"3681E873",
    x"3681B5BE",
    x"3681831D",
    x"3681508F",
    x"36811E16",
    x"3680EBB0",
    x"3680B95D",
    x"3680871F",
    x"368054F4",
    x"368022DC",
    x"367FE1B1",
    x"367F7DD1",
    x"367F1A17",
    x"367EB684",
    x"367E5318",
    x"367DEFD3",
    x"367D8CB5",
    x"367D29BD",
    x"367CC6EC",
    x"367C6442",
    x"367C01BE",
    x"367B9F60",
    x"367B3D29",
    x"367ADB19",
    x"367A792E",
    x"367A176A",
    x"3679B5CC",
    x"36795454",
    x"3678F302",
    x"367891D6",
    x"367830D0",
    x"3677CFF0",
    x"36776F36",
    x"36770EA1",
    x"3676AE32",
    x"36764DE9",
    x"3675EDC5",
    x"36758DC7",
    x"36752DEE",
    x"3674CE3B",
    x"36746EAD",
    x"36740F45",
    x"3673B001",
    x"367350E3",
    x"3672F1EA",
    x"36729316",
    x"36723467",
    x"3671D5DD",
    x"36717778",
    x"36711938",
    x"3670BB1C",
    x"36705D26",
    x"366FFF54",
    x"366FA1A6",
    x"366F441D",
    x"366EE6B9",
    x"366E8979",
    x"366E2C5E",
    x"366DCF66",
    x"366D7293",
    x"366D15E5",
    x"366CB95A",
    x"366C5CF4",
    x"366C00B2",
    x"366BA493",
    x"366B4899",
    x"366AECC3",
    x"366A9110",
    x"366A3581",
    x"3669DA16",
    x"36697ECF",
    x"366923AB",
    x"3668C8AB",
    x"36686DCE",
    x"36681315",
    x"3667B880",
    x"36675E0D",
    x"366703BE",
    x"3666A992",
    x"36664F8A",
    x"3665F5A4",
    x"36659BE2",
    x"36654242",
    x"3664E8C6",
    x"36648F6C",
    x"36643636",
    x"3663DD22",
    x"36638431",
    x"36632B63",
    x"3662D2B7",
    x"36627A2E",
    x"366221C8",
    x"3661C984",
    x"36617162",
    x"36611963",
    x"3660C186",
    x"366069CC",
    x"36601234",
    x"365FBABE",
    x"365F636A",
    x"365F0C38",
    x"365EB528",
    x"365E5E3A",
    x"365E076F",
    x"365DB0C5",
    x"365D5A3C",
    x"365D03D6",
    x"365CAD91",
    x"365C576E",
    x"365C016D",
    x"365BAB8D",
    x"365B55CF",
    x"365B0032",
    x"365AAAB7",
    x"365A555D",
    x"365A0024",
    x"3659AB0D",
    x"36595616",
    x"36590141",
    x"3658AC8E",
    x"365857FB",
    x"36580389",
    x"3657AF38",
    x"36575B08",
    x"365706F9",
    x"3656B30A",
    x"36565F3D",
    x"36560B90",
    x"3655B804",
    x"36556498",
    x"3655114D",
    x"3654BE23",
    x"36546B19",
    x"3654182F",
    x"3653C566",
    x"365372BD",
    x"36532034",
    x"3652CDCC",
    x"36527B83",
    x"3652295B",
    x"3651D753",
    x"3651856B",
    x"365133A3",
    x"3650E1FA",
    x"36509072",
    x"36503F0A",
    x"364FEDC1",
    x"364F9C98",
    x"364F4B8E",
    x"364EFAA5",
    x"364EA9DB",
    x"364E5930",
    x"364E08A5",
    x"364DB839",
    x"364D67ED",
    x"364D17C0",
    x"364CC7B2",
    x"364C77C4",
    x"364C27F5",
    x"364BD845",
    x"364B88B4",
    x"364B3942",
    x"364AE9EF",
    x"364A9ABB",
    x"364A4BA6",
    x"3649FCB0",
    x"3649ADD9",
    x"36495F20",
    x"36491086",
    x"3648C20B",
    x"364873AF",
    x"36482571",
    x"3647D752",
    x"36478951",
    x"36473B6E",
    x"3646EDAA",
    x"3646A005",
    x"3646527D",
    x"36460514",
    x"3645B7C9",
    x"36456A9D",
    x"36451D8E",
    x"3644D09D",
    x"364483CB",
    x"36443716",
    x"3643EA80",
    x"36439E07",
    x"364351AC",
    x"3643056F",
    x"3642B950",
    x"36426D4F",
    x"3642216B",
    x"3641D5A5",
    x"364189FC",
    x"36413E71",
    x"3640F303",
    x"3640A7B3",
    x"36405C80",
    x"3640116B",
    x"363FC672",
    x"363F7B98",
    x"363F30DA",
    x"363EE639",
    x"363E9BB6",
    x"363E5150",
    x"363E0706",
    x"363DBCDA",
    x"363D72CB",
    x"363D28D8",
    x"363CDF03",
    x"363C954A",
    x"363C4BAE",
    x"363C022F",
    x"363BB8CD",
    x"363B6F87",
    x"363B265D",
    x"363ADD51",
    x"363A9461",
    x"363A4B8D",
    x"363A02D5",
    x"3639BA3B",
    x"363971BC",
    x"3639295A",
    x"3638E114",
    x"363898EA",
    x"363850DC",
    x"363808EB",
    x"3637C115",
    x"3637795C",
    x"363731BE",
    x"3636EA3D",
    x"3636A2D7",
    x"36365B8E",
    x"36361460",
    x"3635CD4E",
    x"36358657",
    x"36353F7D",
    x"3634F8BE",
    x"3634B21A",
    x"36346B93",
    x"36342526",
    x"3633DED6",
    x"363398A0",
    x"36335286",
    x"36330C88",
    x"3632C6A5",
    x"363280DD",
    x"36323B30",
    x"3631F59E",
    x"3631B028",
    x"36316ACD",
    x"3631258C",
    x"3630E067",
    x"36309B5D",
    x"3630566E",
    x"3630119A",
    x"362FCCE0",
    x"362F8842",
    x"362F43BE",
    x"362EFF55",
    x"362EBB06",
    x"362E76D2",
    x"362E32B9",
    x"362DEEBB",
    x"362DAAD7",
    x"362D670D",
    x"362D235E",
    x"362CDFCA",
    x"362C9C4F",
    x"362C58F0",
    x"362C15AA",
    x"362BD27F",
    x"362B8F6E",
    x"362B4C77",
    x"362B099A",
    x"362AC6D7",
    x"362A842E",
    x"362A41A0",
    x"3629FF2B",
    x"3629BCD0",
    x"36297A90",
    x"36293869",
    x"3628F65C",
    x"3628B468",
    x"3628728F",
    x"362830CF",
    x"3627EF28",
    x"3627AD9C",
    x"36276C29",
    x"36272ACF",
    x"3626E98F",
    x"3626A869",
    x"3626675C",
    x"36262668",
    x"3625E58E",
    x"3625A4CD",
    x"36256425",
    x"36252396",
    x"3624E321",
    x"3624A2C5",
    x"36246282",
    x"36242258",
    x"3623E247",
    x"3623A24F",
    x"36236270",
    x"362322AA",
    x"3622E2FD",
    x"3622A369",
    x"362263EE",
    x"3622248B",
    x"3621E541",
    x"3621A610",
    x"362166F7",
    x"362127F7",
    x"3620E910",
    x"3620AA41",
    x"36206B8B",
    x"36202CED",
    x"361FEE68",
    x"361FAFFB",
    x"361F71A6",
    x"361F336A",
    x"361EF546",
    x"361EB73A",
    x"361E7947",
    x"361E3B6C",
    x"361DFDA9",
    x"361DBFFE",
    x"361D826B",
    x"361D44F0",
    x"361D078D",
    x"361CCA42",
    x"361C8D0F",
    x"361C4FF4",
    x"361C12F0",
    x"361BD605",
    x"361B9931",
    x"361B5C75",
    x"361B1FD1",
    x"361AE344",
    x"361AA6CF",
    x"361A6A72",
    x"361A2E2C",
    x"3619F1FE",
    x"3619B5E7",
    x"361979E8",
    x"36193E00",
    x"3619022F",
    x"3618C676",
    x"36188AD4",
    x"36184F4A",
    x"361813D6",
    x"3617D87A",
    x"36179D35",
    x"36176207",
    x"361726F0",
    x"3616EBF1",
    x"3616B108",
    x"36167636",
    x"36163B7C",
    x"361600D8",
    x"3615C64B",
    x"36158BD5",
    x"36155176",
    x"3615172D",
    x"3614DCFC",
    x"3614A2E1",
    x"361468DC",
    x"36142EEF",
    x"3613F518",
    x"3613BB57",
    x"361381AD",
    x"3613481A",
    x"36130E9D",
    x"3612D537",
    x"36129BE6",
    x"361262AD",
    x"36122989",
    x"3611F07C",
    x"3611B785",
    x"36117EA5",
    x"361145DB",
    x"36110D26",
    x"3610D488",
    x"36109C00",
    x"3610638E",
    x"36102B32",
    x"360FF2ED",
    x"360FBABD",
    x"360F82A3",
    x"360F4A9F",
    x"360F12B0",
    x"360EDAD8",
    x"360EA315",
    x"360E6B69",
    x"360E33D1",
    x"360DFC50",
    x"360DC4E4",
    x"360D8D8E",
    x"360D564E",
    x"360D1F23",
    x"360CE80D",
    x"360CB10D",
    x"360C7A23",
    x"360C434E",
    x"360C0C8E",
    x"360BD5E4",
    x"360B9F4F",
    x"360B68D0",
    x"360B3265",
    x"360AFC10",
    x"360AC5D1",
    x"360A8FA6",
    x"360A5990",
    x"360A2390",
    x"3609EDA4",
    x"3609B7CE",
    x"3609820D",
    x"36094C61",
    x"360916C9",
    x"3608E147",
    x"3608ABD9",
    x"36087680",
    x"3608413D",
    x"36080C0E",
    x"3607D6F3",
    x"3607A1EE",
    x"36076CFD",
    x"36073820",
    x"36070359",
    x"3606CEA6",
    x"36069A07",
    x"3606657D",
    x"36063108",
    x"3605FCA7",
    x"3605C85B",
    x"36059423",
    x"36055FFF",
    x"36052BF0",
    x"3604F7F5",
    x"3604C40E",
    x"3604903B",
    x"36045C7D",
    x"360428D3",
    x"3603F53D",
    x"3603C1BC",
    x"36038E4E",
    x"36035AF4",
    x"360327AF",
    x"3602F47D",
    x"3602C160",
    x"36028E56",
    x"36025B61",
    x"3602287F",
    x"3601F5B1",
    x"3601C2F7",
    x"36019051",
    x"36015DBE",
    x"36012B3F",
    x"3600F8D4",
    x"3600C67D",
    x"36009439",
    x"36006209",
    x"36002FED",
    x"35FFFBC7",
    x"35FF97DD",
    x"35FF3419",
    x"35FED07C",
    x"35FE6D06",
    x"35FE09B7",
    x"35FDA68E",
    x"35FD438D",
    x"35FCE0B1",
    x"35FC7DFD",
    x"35FC1B6F",
    x"35FBB908",
    x"35FB56C6",
    x"35FAF4AC",
    x"35FA92B7",
    x"35FA30E9",
    x"35F9CF41",
    x"35F96DBF",
    x"35F90C63",
    x"35F8AB2D",
    x"35F84A1E",
    x"35F7E934",
    x"35F7886F",
    x"35F727D1",
    x"35F6C758",
    x"35F66705",
    x"35F606D8",
    x"35F5A6D0",
    x"35F546ED",
    x"35F4E730",
    x"35F48799",
    x"35F42826",
    x"35F3C8D9",
    x"35F369B1",
    x"35F30AAF",
    x"35F2ABD1",
    x"35F24D18",
    x"35F1EE85",
    x"35F19016",
    x"35F131CC",
    x"35F0D3A7",
    x"35F075A7",
    x"35F017CB",
    x"35EFBA14",
    x"35EF5C82",
    x"35EEFF14",
    x"35EEA1CB",
    x"35EE44A6",
    x"35EDE7A5",
    x"35ED8AC9",
    x"35ED2E10",
    x"35ECD17D",
    x"35EC750D",
    x"35EC18C1",
    x"35EBBC99",
    x"35EB6096",
    x"35EB04B6",
    x"35EAA8FA",
    x"35EA4D62",
    x"35E9F1EE",
    x"35E9969D",
    x"35E93B70",
    x"35E8E066",
    x"35E88581",
    x"35E82ABE",
    x"35E7D01F",
    x"35E775A4",
    x"35E71B4B",
    x"35E6C116",
    x"35E66704",
    x"35E60D16",
    x"35E5B34A",
    x"35E559A2",
    x"35E5001C",
    x"35E4A6BA",
    x"35E44D7A",
    x"35E3F45D",
    x"35E39B63",
    x"35E3428C",
    x"35E2E9D7",
    x"35E29145",
    x"35E238D5",
    x"35E1E088",
    x"35E1885E",
    x"35E13056",
    x"35E0D870",
    x"35E080AD",
    x"35E0290C",
    x"35DFD18D",
    x"35DF7A30",
    x"35DF22F5",
    x"35DECBDD",
    x"35DE74E6",
    x"35DE1E11",
    x"35DDC75E",
    x"35DD70CD",
    x"35DD1A5E",
    x"35DCC411",
    x"35DC6DE5",
    x"35DC17DB",
    x"35DBC1F2",
    x"35DB6C2B",
    x"35DB1686",
    x"35DAC102",
    x"35DA6B9F",
    x"35DA165E",
    x"35D9C13E",
    x"35D96C3F",
    x"35D91761",
    x"35D8C2A4",
    x"35D86E09",
    x"35D8198E",
    x"35D7C535",
    x"35D770FC",
    x"35D71CE5",
    x"35D6C8EE",
    x"35D67518",
    x"35D62162",
    x"35D5CDCE",
    x"35D57A59",
    x"35D52706",
    x"35D4D3D3",
    x"35D480C0",
    x"35D42DCE",
    x"35D3DAFD",
    x"35D3884B",
    x"35D335BA",
    x"35D2E349",
    x"35D290F9",
    x"35D23EC8",
    x"35D1ECB8",
    x"35D19AC7",
    x"35D148F7",
    x"35D0F746",
    x"35D0A5B5",
    x"35D05445",
    x"35D002F4",
    x"35CFB1C2",
    x"35CF60B1",
    x"35CF0FBF",
    x"35CEBEEC",
    x"35CE6E3A",
    x"35CE1DA6",
    x"35CDCD32",
    x"35CD7CDE",
    x"35CD2CA9",
    x"35CCDC93",
    x"35CC8C9C",
    x"35CC3CC5",
    x"35CBED0D",
    x"35CB9D74",
    x"35CB4DFA",
    x"35CAFE9F",
    x"35CAAF63",
    x"35CA6046",
    x"35CA1148",
    x"35C9C268",
    x"35C973A8",
    x"35C92506",
    x"35C8D683",
    x"35C8881E",
    x"35C839D9",
    x"35C7EBB1",
    x"35C79DA8",
    x"35C74FBE",
    x"35C701F2",
    x"35C6B444",
    x"35C666B5",
    x"35C61944",
    x"35C5CBF1",
    x"35C57EBD",
    x"35C531A6",
    x"35C4E4AE",
    x"35C497D4",
    x"35C44B17",
    x"35C3FE79",
    x"35C3B1F9",
    x"35C36596",
    x"35C31951",
    x"35C2CD2A",
    x"35C28121",
    x"35C23535",
    x"35C1E967",
    x"35C19DB7",
    x"35C15224",
    x"35C106AF",
    x"35C0BB57",
    x"35C0701C",
    x"35C024FF",
    x"35BFDA00",
    x"35BF8F1D",
    x"35BF4458",
    x"35BEF9B0",
    x"35BEAF25",
    x"35BE64B7",
    x"35BE1A66",
    x"35BDD032",
    x"35BD861B",
    x"35BD3C21",
    x"35BCF244",
    x"35BCA884",
    x"35BC5EE1",
    x"35BC155A",
    x"35BBCBF0",
    x"35BB82A3",
    x"35BB3972",
    x"35BAF05E",
    x"35BAA766",
    x"35BA5E8B",
    x"35BA15CC",
    x"35B9CD2A",
    x"35B984A4",
    x"35B93C3A",
    x"35B8F3ED",
    x"35B8ABBC",
    x"35B863A7",
    x"35B81BAE",
    x"35B7D3D1",
    x"35B78C10",
    x"35B7446C",
    x"35B6FCE3",
    x"35B6B576",
    x"35B66E25",
    x"35B626F0",
    x"35B5DFD7",
    x"35B598D9",
    x"35B551F7",
    x"35B50B31",
    x"35B4C486",
    x"35B47DF7",
    x"35B43784",
    x"35B3F12C",
    x"35B3AAF0",
    x"35B364CE",
    x"35B31EC9",
    x"35B2D8DE",
    x"35B2930F",
    x"35B24D5B",
    x"35B207C3",
    x"35B1C245",
    x"35B17CE3",
    x"35B1379C",
    x"35B0F270",
    x"35B0AD5E",
    x"35B06868",
    x"35B0238D",
    x"35AFDECC",
    x"35AF9A27",
    x"35AF559C",
    x"35AF112C",
    x"35AECCD6",
    x"35AE889C",
    x"35AE447C",
    x"35AE0076",
    x"35ADBC8B",
    x"35AD78BB",
    x"35AD3505",
    x"35ACF16A",
    x"35ACADE8",
    x"35AC6A82",
    x"35AC2735",
    x"35ABE403",
    x"35ABA0EB",
    x"35AB5DED",
    x"35AB1B0A",
    x"35AAD840",
    x"35AA9591",
    x"35AA52FB",
    x"35AA1080",
    x"35A9CE1E",
    x"35A98BD7",
    x"35A949A9",
    x"35A90795",
    x"35A8C59B",
    x"35A883BB",
    x"35A841F4",
    x"35A80047",
    x"35A7BEB4",
    x"35A77D3A",
    x"35A73BDA",
    x"35A6FA94",
    x"35A6B966",
    x"35A67853",
    x"35A63758",
    x"35A5F677",
    x"35A5B5B0",
    x"35A57501",
    x"35A5346C",
    x"35A4F3F1",
    x"35A4B38E",
    x"35A47344",
    x"35A43314",
    x"35A3F2FC",
    x"35A3B2FE",
    x"35A37318",
    x"35A3334C",
    x"35A2F398",
    x"35A2B3FE",
    x"35A2747C",
    x"35A23513",
    x"35A1F5C2",
    x"35A1B68B",
    x"35A1776C",
    x"35A13865",
    x"35A0F978",
    x"35A0BAA2",
    x"35A07BE6",
    x"35A03D42",
    x"359FFEB6",
    x"359FC043",
    x"359F81E8",
    x"359F43A5",
    x"359F057B",
    x"359EC769",
    x"359E896F",
    x"359E4B8D",
    x"359E0DC4",
    x"359DD013",
    x"359D9279",
    x"359D54F8",
    x"359D178F",
    x"359CDA3E",
    x"359C9D04",
    x"359C5FE3",
    x"359C22DA",
    x"359BE5E8",
    x"359BA90E",
    x"359B6C4C",
    x"359B2FA1",
    x"359AF30F",
    x"359AB693",
    x"359A7A30",
    x"359A3DE4",
    x"359A01B0",
    x"3599C593",
    x"3599898D",
    x"35994D9F",
    x"359911C9",
    x"3598D609",
    x"35989A61",
    x"35985ED1",
    x"35982357",
    x"3597E7F5",
    x"3597ACAA",
    x"35977176",
    x"35973659",
    x"3596FB54",
    x"3596C065",
    x"3596858D",
    x"35964ACD",
    x"35961023",
    x"3595D590",
    x"35959B14",
    x"359560AF",
    x"35952660",
    x"3594EC29",
    x"3594B208",
    x"359477FE",
    x"35943E0A",
    x"3594042D",
    x"3593CA67",
    x"359390B7",
    x"3593571E",
    x"35931D9B",
    x"3592E42F",
    x"3592AAD9",
    x"35927199",
    x"35923870",
    x"3591FF5D",
    x"3591C660",
    x"35918D7A",
    x"359154AA",
    x"35911BF0",
    x"3590E34C",
    x"3590AABE",
    x"35907247",
    x"359039E5",
    x"35900199",
    x"358FC964",
    x"358F9144",
    x"358F593A",
    x"358F2146",
    x"358EE968",
    x"358EB1A0",
    x"358E79EE",
    x"358E4251",
    x"358E0ACA",
    x"358DD358",
    x"358D9BFD",
    x"358D64B6",
    x"358D2D86",
    x"358CF66B",
    x"358CBF65",
    x"358C8875",
    x"358C519B",
    x"358C1AD6",
    x"358BE426",
    x"358BAD8B",
    x"358B7706",
    x"358B4096",
    x"358B0A3C",
    x"358AD3F6",
    x"358A9DC6",
    x"358A67AB",
    x"358A31A5",
    x"3589FBB4",
    x"3589C5D8",
    x"35899012",
    x"35895A60",
    x"358924C3",
    x"3588EF3B",
    x"3588B9C8",
    x"3588846A",
    x"35884F21",
    x"358819EC",
    x"3587E4CC",
    x"3587AFC1",
    x"35877ACB",
    x"358745E9",
    x"3587111C",
    x"3586DC64",
    x"3586A7C0",
    x"35867331",
    x"35863EB6",
    x"35860A50",
    x"3585D5FE",
    x"3585A1C1",
    x"35856D98",
    x"35853983",
    x"35850583",
    x"3584D197",
    x"35849DBF",
    x"358469FC",
    x"3584364C",
    x"358402B1",
    x"3583CF2A",
    x"35839BB7",
    x"35836859",
    x"3583350E",
    x"358301D7",
    x"3582CEB4",
    x"35829BA6",
    x"358268AB",
    x"358235C4",
    x"358202F1",
    x"3581D032",
    x"35819D86",
    x"35816AEE",
    x"3581386B",
    x"358105FA",
    x"3580D39E",
    x"3580A155",
    x"35806F20",
    x"35803CFE",
    x"35800AF0",
    x"357FB1EB",
    x"357F4E1D",
    x"357EEA76",
    x"357E86F6",
    x"357E239D",
    x"357DC06A",
    x"357D5D5E",
    x"357CFA79",
    x"357C97BB",
    x"357C3523",
    x"357BD2B1",
    x"357B7066",
    x"357B0E41",
    x"357AAC43",
    x"357A4A6B",
    x"3579E8B9",
    x"3579872D",
    x"357925C7",
    x"3578C487",
    x"3578636E",
    x"3578027A",
    x"3577A1AC",
    x"35774103",
    x"3576E081",
    x"35768024",
    x"35761FED",
    x"3575BFDB",
    x"35755FEF",
    x"35750028",
    x"3574A087",
    x"3574410B",
    x"3573E1B4",
    x"35738282",
    x"35732376",
    x"3572C48F",
    x"357265CC",
    x"3572072F",
    x"3571A8B7",
    x"35714A63",
    x"3570EC35",
    x"35708E2B",
    x"35703045",
    x"356FD285",
    x"356F74E9",
    x"356F1772",
    x"356EBA1F",
    x"356E5CF0",
    x"356DFFE6",
    x"356DA300",
    x"356D463F",
    x"356CE9A1",
    x"356C8D28",
    x"356C30D3",
    x"356BD4A2",
    x"356B7895",
    x"356B1CAC",
    x"356AC0E6",
    x"356A6545",
    x"356A09C7",
    x"3569AE6D",
    x"35695337",
    x"3568F824",
    x"35689D35",
    x"35684269",
    x"3567E7C1",
    x"35678D3C",
    x"356732DB",
    x"3566D89D",
    x"35667E82",
    x"3566248A",
    x"3565CAB5",
    x"35657103",
    x"35651775",
    x"3564BE09",
    x"356464C0",
    x"35640B9A",
    x"3563B297",
    x"356359B7",
    x"356300F9",
    x"3562A85E",
    x"35624FE6",
    x"3561F790",
    x"35619F5C",
    x"3561474B",
    x"3560EF5C",
    x"35609790",
    x"35603FE6",
    x"355FE85E",
    x"355F90F8",
    x"355F39B5",
    x"355EE293",
    x"355E8B94",
    x"355E34B6",
    x"355DDDFB",
    x"355D8761",
    x"355D30E9",
    x"355CDA93",
    x"355C845E",
    x"355C2E4B",
    x"355BD85A",
    x"355B828A",
    x"355B2CDC",
    x"355AD74F",
    x"355A81E4",
    x"355A2C9A",
    x"3559D771",
    x"35598269",
    x"35592D83",
    x"3558D8BE",
    x"35588419",
    x"35582F96",
    x"3557DB34",
    x"355786F3",
    x"355732D3",
    x"3556DED3",
    x"35568AF5",
    x"35563737",
    x"3555E39A",
    x"3555901D",
    x"35553CC1",
    x"3554E986",
    x"3554966B",
    x"35544370",
    x"3553F096",
    x"35539DDC",
    x"35534B42",
    x"3552F8C9",
    x"3552A670",
    x"35525437",
    x"3552021E",
    x"3551B025",
    x"35515E4D",
    x"35510C94",
    x"3550BAFB",
    x"35506982",
    x"35501828",
    x"354FC6EF",
    x"354F75D5",
    x"354F24DB",
    x"354ED400",
    x"354E8345",
    x"354E32AA",
    x"354DE22E",
    x"354D91D1",
    x"354D4194",
    x"354CF176",
    x"354CA177",
    x"354C5197",
    x"354C01D7",
    x"354BB236",
    x"354B62B4",
    x"354B1351",
    x"354AC40D",
    x"354A74E8",
    x"354A25E1",
    x"3549D6FA",
    x"35498832",
    x"35493988",
    x"3548EAFD",
    x"35489C90",
    x"35484E42",
    x"35480013",
    x"3547B202",
    x"35476410",
    x"3547163C",
    x"3546C886",
    x"35467AEF",
    x"35462D76",
    x"3545E01C",
    x"354592DF",
    x"354545C1",
    x"3544F8C1",
    x"3544ABDF",
    x"35445F1A",
    x"35441274",
    x"3543C5EC",
    x"35437982",
    x"35432D35",
    x"3542E106",
    x"354294F5",
    x"35424902",
    x"3541FD2C",
    x"3541B174",
    x"354165DA",
    x"35411A5D",
    x"3540CEFD",
    x"354083BB",
    x"35403896",
    x"353FED8F",
    x"353FA2A4",
    x"353F57D8",
    x"353F0D28",
    x"353EC295",
    x"353E7820",
    x"353E2DC7",
    x"353DE38C",
    x"353D996E",
    x"353D4F6C",
    x"353D0588",
    x"353CBBC0",
    x"353C7215",
    x"353C2887",
    x"353BDF15",
    x"353B95C0",
    x"353B4C88",
    x"353B036D",
    x"353ABA6D",
    x"353A718B",
    x"353A28C5",
    x"3539E01B",
    x"3539978E",
    x"35394F1D",
    x"353906C8",
    x"3538BE8F",
    x"35387673",
    x"35382E73",
    x"3537E68F",
    x"35379EC7",
    x"3537571B",
    x"35370F8B",
    x"3536C816",
    x"353680BE",
    x"35363982",
    x"3535F261",
    x"3535AB5C",
    x"35356473",
    x"35351DA6",
    x"3534D6F4",
    x"3534905E",
    x"353449E3",
    x"35340384",
    x"3533BD41",
    x"35337718",
    x"3533310C",
    x"3532EB1A",
    x"3532A544",
    x"35325F89",
    x"353219E9",
    x"3531D465",
    x"35318EFB",
    x"353149AD",
    x"3531047A",
    x"3530BF61",
    x"35307A64",
    x"35303582",
    x"352FF0BA",
    x"352FAC0E",
    x"352F677C",
    x"352F2305",
    x"352EDEA9",
    x"352E9A67",
    x"352E5640",
    x"352E1234",
    x"352DCE42",
    x"352D8A6A",
    x"352D46AE",
    x"352D030B",
    x"352CBF83",
    x"352C7C16",
    x"352C38C2",
    x"352BF589",
    x"352BB26A",
    x"352B6F66",
    x"352B2C7B",
    x"352AE9AB",
    x"352AA6F5",
    x"352A6459",
    x"352A21D6",
    x"3529DF6E",
    x"35299D20",
    x"35295AEB",
    x"352918D1",
    x"3528D6D0",
    x"352894E9",
    x"3528531C",
    x"35281168",
    x"3527CFCE",
    x"35278E4E",
    x"35274CE7",
    x"35270B99",
    x"3526CA66",
    x"3526894B",
    x"3526484A",
    x"35260763",
    x"3525C695",
    x"352585E0",
    x"35254544",
    x"352504C2",
    x"3524C458",
    x"35248408",
    x"352443D1",
    x"352403B3",
    x"3523C3AE",
    x"352383C2",
    x"352343EF",
    x"35230435",
    x"3522C494",
    x"3522850C",
    x"3522459C",
    x"35220645",
    x"3521C707",
    x"352187E2",
    x"352148D5",
    x"352109E1",
    x"3520CB05",
    x"35208C42",
    x"35204D98",
    x"35200F06",
    x"351FD08C",
    x"351F922B",
    x"351F53E2",
    x"351F15B1",
    x"351ED799",
    x"351E9999",
    x"351E5BB1",
    x"351E1DE1",
    x"351DE029",
    x"351DA28A",
    x"351D6502",
    x"351D2793",
    x"351CEA3B",
    x"351CACFC",
    x"351C6FD4",
    x"351C32C5",
    x"351BF5CD",
    x"351BB8EC",
    x"351B7C24",
    x"351B3F73",
    x"351B02DB",
    x"351AC659",
    x"351A89F0",
    x"351A4D9D",
    x"351A1163",
    x"3519D540",
    x"35199934",
    x"35195D40",
    x"35192163",
    x"3518E59E",
    x"3518A9F0",
    x"35186E59",
    x"351832DA",
    x"3517F772",
    x"3517BC21",
    x"351780E7",
    x"351745C4",
    x"35170AB8",
    x"3516CFC3",
    x"351694E6",
    x"35165A1F",
    x"35161F6F",
    x"3515E4D6",
    x"3515AA55",
    x"35156FE9",
    x"35153595",
    x"3514FB58",
    x"3514C131",
    x"35148721",
    x"35144D27",
    x"35141344",
    x"3513D978",
    x"35139FC2",
    x"35136623",
    x"35132C9B",
    x"3512F328",
    x"3512B9CD",
    x"35128087",
    x"35124758",
    x"35120E3F",
    x"3511D53D",
    x"35119C51",
    x"3511637B",
    x"35112ABB",
    x"3510F212",
    x"3510B97E",
    x"35108101",
    x"35104899",
    x"35101048",
    x"350FD80C",
    x"350F9FE7",
    x"350F67D8",
    x"350F2FDE",
    x"350EF7FA",
    x"350EC02C",
    x"350E8874",
    x"350E50D2",
    x"350E1945",
    x"350DE1CE",
    x"350DAA6C",
    x"350D7321",
    x"350D3BEA",
    x"350D04CA",
    x"350CCDBF",
    x"350C96C9",
    x"350C5FE9",
    x"350C291E",
    x"350BF269",
    x"350BBBC9",
    x"350B853E",
    x"350B4EC9",
    x"350B1868",
    x"350AE21E",
    x"350AABE8",
    x"350A75C7",
    x"350A3FBC",
    x"350A09C5",
    x"3509D3E4",
    x"35099E18",
    x"35096861",
    x"350932BE",
    x"3508FD31",
    x"3508C7B9",
    x"35089255",
    x"35085D06",
    x"350827CC",
    x"3507F2A7",
    x"3507BD97",
    x"3507889B",
    x"350753B4",
    x"35071EE2",
    x"3506EA24",
    x"3506B57B",
    x"350680E6",
    x"35064C66",
    x"350617FA",
    x"3505E3A3",
    x"3505AF60",
    x"35057B32",
    x"35054718",
    x"35051313",
    x"3504DF21",
    x"3504AB44",
    x"3504777B",
    x"350443C7",
    x"35041027",
    x"3503DC9A",
    x"3503A922",
    x"350375BE",
    x"3503426E",
    x"35030F32",
    x"3502DC0A",
    x"3502A8F6",
    x"350275F6",
    x"3502430A",
    x"35021032",
    x"3501DD6D",
    x"3501AABD",
    x"35017820",
    x"35014597",
    x"35011322",
    x"3500E0C0",
    x"3500AE72",
    x"35007C38",
    x"35004A11",
    x"350017FE",
    x"34FFCBFD",
    x"34FF6824",
    x"34FF0473",
    x"34FEA0E9",
    x"34FE3D86",
    x"34FDDA49",
    x"34FD7733",
    x"34FD1444",
    x"34FCB17B",
    x"34FC4ED9",
    x"34FBEC5D",
    x"34FB8A08",
    x"34FB27DA",
    x"34FAC5D1",
    x"34FA63EF",
    x"34FA0233",
    x"34F9A09D",
    x"34F93F2E",
    x"34F8DDE4",
    x"34F87CC0",
    x"34F81BC2",
    x"34F7BAEB",
    x"34F75A38",
    x"34F6F9AC",
    x"34F69945",
    x"34F63904",
    x"34F5D8E9",
    x"34F578F3",
    x"34F51922",
    x"34F4B977",
    x"34F459F1",
    x"34F3FA91",
    x"34F39B56",
    x"34F33C3F",
    x"34F2DD4E",
    x"34F27E83",
    x"34F21FDC",
    x"34F1C15A",
    x"34F162FD",
    x"34F104C4",
    x"34F0A6B1",
    x"34F048C2",
    x"34EFEAF8",
    x"34EF8D52",
    x"34EF2FD2",
    x"34EED275",
    x"34EE753D",
    x"34EE1829",
    x"34EDBB3A",
    x"34ED5E6F",
    x"34ED01C8",
    x"34ECA546",
    x"34EC48E7",
    x"34EBECAD",
    x"34EB9096",
    x"34EB34A4",
    x"34EAD8D5",
    x"34EA7D2A",
    x"34EA21A3",
    x"34E9C640",
    x"34E96B00",
    x"34E90FE4",
    x"34E8B4EC",
    x"34E85A17",
    x"34E7FF66",
    x"34E7A4D8",
    x"34E74A6D",
    x"34E6F025",
    x"34E69601",
    x"34E63C00",
    x"34E5E222",
    x"34E58868",
    x"34E52ED0",
    x"34E4D55B",
    x"34E47C09",
    x"34E422DA",
    x"34E3C9CE",
    x"34E370E4",
    x"34E3181E",
    x"34E2BF79",
    x"34E266F8",
    x"34E20E99",
    x"34E1B65D",
    x"34E15E43",
    x"34E1064B",
    x"34E0AE76",
    x"34E056C3",
    x"34DFFF32",
    x"34DFA7C3",
    x"34DF5077",
    x"34DEF94C",
    x"34DEA244",
    x"34DE4B5E",
    x"34DDF499",
    x"34DD9DF6",
    x"34DD4776",
    x"34DCF117",
    x"34DC9AD9",
    x"34DC44BE",
    x"34DBEEC4",
    x"34DB98EB",
    x"34DB4334",
    x"34DAED9F",
    x"34DA982A",
    x"34DA42D8",
    x"34D9EDA6",
    x"34D99896",
    x"34D943A7",
    x"34D8EED9",
    x"34D89A2C",
    x"34D845A1",
    x"34D7F136",
    x"34D79CEC",
    x"34D748C3",
    x"34D6F4BB",
    x"34D6A0D4",
    x"34D64D0E",
    x"34D5F968",
    x"34D5A5E3",
    x"34D5527E",
    x"34D4FF3A",
    x"34D4AC17",
    x"34D45914",
    x"34D40631",
    x"34D3B36F",
    x"34D360CD",
    x"34D30E4B",
    x"34D2BBEA",
    x"34D269A9",
    x"34D21787",
    x"34D1C586",
    x"34D173A5",
    x"34D121E4",
    x"34D0D042",
    x"34D07EC1",
    x"34D02D5F",
    x"34CFDC1E",
    x"34CF8AFB",
    x"34CF39F9",
    x"34CEE916",
    x"34CE9853",
    x"34CE47AF",
    x"34CDF72B",
    x"34CDA6C6",
    x"34CD5681",
    x"34CD065A",
    x"34CCB654",
    x"34CC666C",
    x"34CC16A4",
    x"34CBC6FA",
    x"34CB7770",
    x"34CB2805",
    x"34CAD8B9",
    x"34CA898C",
    x"34CA3A7D",
    x"34C9EB8E",
    x"34C99CBD",
    x"34C94E0B",
    x"34C8FF78",
    x"34C8B104",
    x"34C862AE",
    x"34C81477",
    x"34C7C65E",
    x"34C77864",
    x"34C72A88",
    x"34C6DCCA",
    x"34C68F2B",
    x"34C641AB",
    x"34C5F448",
    x"34C5A704",
    x"34C559DE",
    x"34C50CD6",
    x"34C4BFEC",
    x"34C47320",
    x"34C42672",
    x"34C3D9E2",
    x"34C38D6F",
    x"34C3411B",
    x"34C2F4E4",
    x"34C2A8CC",
    x"34C25CD1",
    x"34C210F3",
    x"34C1C533",
    x"34C17991",
    x"34C12E0C",
    x"34C0E2A5",
    x"34C0975B",
    x"34C04C2F",
    x"34C00120",
    x"34BFB62E",
    x"34BF6B59",
    x"34BF20A2",
    x"34BED608",
    x"34BE8B8B",
    x"34BE412B",
    x"34BDF6E8",
    x"34BDACC2",
    x"34BD62B9",
    x"34BD18CD",
    x"34BCCEFD",
    x"34BC854B",
    x"34BC3BB5",
    x"34BBF23C",
    x"34BBA8E0",
    x"34BB5FA0",
    x"34BB167D",
    x"34BACD77",
    x"34BA848D",
    x"34BA3BBF",
    x"34B9F30E",
    x"34B9AA79",
    x"34B96201",
    x"34B919A5",
    x"34B8D165",
    x"34B88941",
    x"34B8413A",
    x"34B7F94E",
    x"34B7B17F",
    x"34B769CC",
    x"34B72234",
    x"34B6DAB9",
    x"34B69359",
    x"34B64C16",
    x"34B604EE",
    x"34B5BDE2",
    x"34B576F1",
    x"34B5301D",
    x"34B4E964",
    x"34B4A2C7",
    x"34B45C45",
    x"34B415DE",
    x"34B3CF94",
    x"34B38964",
    x"34B34350",
    x"34B2FD58",
    x"34B2B77A",
    x"34B271B8",
    x"34B22C11",
    x"34B1E686",
    x"34B1A115",
    x"34B15BC0",
    x"34B11686",
    x"34B0D166",
    x"34B08C62",
    x"34B04779",
    x"34B002AA",
    x"34AFBDF7",
    x"34AF795E",
    x"34AF34E0",
    x"34AEF07C",
    x"34AEAC34",
    x"34AE6806",
    x"34AE23F3",
    x"34ADDFFA",
    x"34AD9C1C",
    x"34AD5858",
    x"34AD14AF",
    x"34ACD120",
    x"34AC8DAB",
    x"34AC4A51",
    x"34AC0711",
    x"34ABC3EB",
    x"34AB80E0",
    x"34AB3DEF",
    x"34AAFB18",
    x"34AAB85B",
    x"34AA75B8",
    x"34AA332F",
    x"34A9F0C0",
    x"34A9AE6A",
    x"34A96C2F",
    x"34A92A0E",
    x"34A8E806",
    x"34A8A619",
    x"34A86445",
    x"34A8228A",
    x"34A7E0EA",
    x"34A79F63",
    x"34A75DF5",
    x"34A71CA1",
    x"34A6DB67",
    x"34A69A46",
    x"34A6593E",
    x"34A61850",
    x"34A5D77B",
    x"34A596C0",
    x"34A5561D",
    x"34A51594",
    x"34A4D525",
    x"34A494CE",
    x"34A45490",
    x"34A4146C",
    x"34A3D460",
    x"34A3946E",
    x"34A35494",
    x"34A314D4",
    x"34A2D52C",
    x"34A2959D",
    x"34A25627",
    x"34A216CA",
    x"34A1D785",
    x"34A19859",
    x"34A15946",
    x"34A11A4C",
    x"34A0DB6A",
    x"34A09CA0",
    x"34A05DEF",
    x"34A01F57",
    x"349FE0D7",
    x"349FA26F",
    x"349F6420",
    x"349F25E9",
    x"349EE7CA",
    x"349EA9C4",
    x"349E6BD6",
    x"349E2E00",
    x"349DF042",
    x"349DB29C",
    x"349D750E",
    x"349D3798",
    x"349CFA3B",
    x"349CBCF5",
    x"349C7FC7",
    x"349C42B1",
    x"349C05B3",
    x"349BC8CD",
    x"349B8BFE",
    x"349B4F47",
    x"349B12A8",
    x"349AD621",
    x"349A99B1",
    x"349A5D59",
    x"349A2118",
    x"3499E4EF",
    x"3499A8DD",
    x"34996CE3",
    x"34993100",
    x"3498F535",
    x"3498B980",
    x"34987DE4",
    x"3498425E",
    x"349806F0",
    x"3497CB99",
    x"34979059",
    x"34975530",
    x"34971A1E",
    x"3496DF23",
    x"3496A440",
    x"34966973",
    x"34962EBD",
    x"3495F41F",
    x"3495B997",
    x"34957F26",
    x"349544CB",
    x"34950A88",
    x"3494D05B",
    x"34949645",
    x"34945C46",
    x"3494225D",
    x"3493E88B",
    x"3493AECF",
    x"3493752A",
    x"34933B9C",
    x"34930224",
    x"3492C8C2",
    x"34928F77",
    x"34925642",
    x"34921D23",
    x"3491E41B",
    x"3491AB29",
    x"3491724D",
    x"34913988",
    x"349100D8",
    x"3490C83F",
    x"34908FBC",
    x"3490574F",
    x"34901EF8",
    x"348FE6B7",
    x"348FAE8B",
    x"348F7676",
    x"348F3E77",
    x"348F068D",
    x"348ECEBA",
    x"348E96FC",
    x"348E5F54",
    x"348E27C1",
    x"348DF045",
    x"348DB8DE",
    x"348D818C",
    x"348D4A51",
    x"348D132A",
    x"348CDC1A",
    x"348CA51E",
    x"348C6E39",
    x"348C3768",
    x"348C00AD",
    x"348BCA08",
    x"348B9377",
    x"348B5CFC",
    x"348B2697",
    x"348AF046",
    x"348ABA0B",
    x"348A83E5",
    x"348A4DD4",
    x"348A17D8",
    x"3489E1F1",
    x"3489AC20",
    x"34897663",
    x"348940BB",
    x"34890B28",
    x"3488D5AA",
    x"3488A041",
    x"34886AED",
    x"348835AE",
    x"34880083",
    x"3487CB6D",
    x"3487966C",
    x"34876180",
    x"34872CA8",
    x"3486F7E5",
    x"3486C336",
    x"34868E9C",
    x"34865A17",
    x"348625A6",
    x"3485F14A",
    x"3485BD01",
    x"348588CE",
    x"348554AF",
    x"348520A4",
    x"3484ECAD",
    x"3484B8CB",
    x"348484FD",
    x"34845143",
    x"34841D9D",
    x"3483EA0C",
    x"3483B68E",
    x"34838325",
    x"34834FD0",
    x"34831C8F",
    x"3482E962",
    x"3482B648",
    x"34828343",
    x"34825052",
    x"34821D74",
    x"3481EAAB",
    x"3481B7F5",
    x"34818553",
    x"348152C5",
    x"3481204A",
    x"3480EDE4",
    x"3480BB91",
    x"34808951",
    x"34805725",
    x"3480250D",
    x"347FE611",
    x"347F822E",
    x"347F1E73",
    x"347EBADE",
    x"347E5771",
    x"347DF42A",
    x"347D910A",
    x"347D2E11",
    x"347CCB3E",
    x"347C6892",
    x"347C060C",
    x"347BA3AD",
    x"347B4174",
    x"347ADF62",
    x"347A7D76",
    x"347A1BB0",
    x"3479BA10",
    x"34795897",
    x"3478F743",
    x"34789615",
    x"3478350E",
    x"3477D42C",
    x"34777370",
    x"347712DA",
    x"3476B269",
    x"3476521E",
    x"3475F1F9",
    x"347591F9",
    x"3475321F",
    x"3474D26A",
    x"347472DB",
    x"34741370",
    x"3473B42B",
    x"3473550C",
    x"3472F611",
    x"3472973B",
    x"3472388B",
    x"3471D9FF",
    x"34717B98",
    x"34711D57",
    x"3470BF3A",
    x"34706141",
    x"3470036E",
    x"346FA5BE",
    x"346F4834",
    x"346EEACE",
    x"346E8D8D",
    x"346E306F",
    x"346DD377",
    x"346D76A2",
    x"346D19F2",
    x"346CBD66",
    x"346C60FE",
    x"346C04BA",
    x"346BA89A",
    x"346B4C9E",
    x"346AF0C6",
    x"346A9512",
    x"346A3982",
    x"3469DE15",
    x"346982CC",
    x"346927A7",
    x"3468CCA5",
    x"346871C7",
    x"3468170D",
    x"3467BC75",
    x"34676201",
    x"346707B1",
    x"3466AD83",
    x"34665379",
    x"3465F992",
    x"34659FCE",
    x"3465462D",
    x"3464ECAF",
    x"34649354",
    x"34643A1C",
    x"3463E107",
    x"34638814",
    x"34632F44",
    x"3462D697",
    x"34627E0D",
    x"346225A5",
    x"3461CD5F",
    x"3461753C",
    x"34611D3C",
    x"3460C55E",
    x"34606DA2",
    x"34601608",
    x"345FBE90",
    x"345F673B",
    x"345F1008",
    x"345EB8F6",
    x"345E6207",
    x"345E0B3A",
    x"345DB48E",
    x"345D5E05",
    x"345D079D",
    x"345CB157",
    x"345C5B32",
    x"345C0530",
    x"345BAF4E",
    x"345B598F",
    x"345B03F0",
    x"345AAE73",
    x"345A5918",
    x"345A03DE",
    x"3459AEC5",
    x"345959CD",
    x"345904F7",
    x"3458B041",
    x"34585BAD",
    x"3458073A",
    x"3457B2E7",
    x"34575EB6",
    x"34570AA5",
    x"3456B6B6",
    x"345662E7",
    x"34560F38",
    x"3455BBAB",
    x"3455683E",
    x"345514F1",
    x"3454C1C5",
    x"34546EBA",
    x"34541BCF",
    x"3453C904",
    x"3453765A",
    x"345323D0",
    x"3452D166",
    x"34527F1C",
    x"34522CF2",
    x"3451DAE9",
    x"345188FF",
    x"34513736",
    x"3450E58C",
    x"34509403",
    x"34504299",
    x"344FF14E",
    x"344FA024",
    x"344F4F19",
    x"344EFE2E",
    x"344EAD63",
    x"344E5CB7",
    x"344E0C2A",
    x"344DBBBD",
    x"344D6B70",
    x"344D1B41",
    x"344CCB32",
    x"344C7B43",
    x"344C2B72",
    x"344BDBC1",
    x"344B8C2E",
    x"344B3CBB",
    x"344AED67",
    x"344A9E32",
    x"344A4F1B",
    x"344A0024",
    x"3449B14B",
    x"34496291",
    x"344913F6",
    x"3448C57A",
    x"3448771C",
    x"344828DD",
    x"3447DABC",
    x"34478CBA",
    x"34473ED6",
    x"3446F111",
    x"3446A36A",
    x"344655E1",
    x"34460876",
    x"3445BB2A",
    x"34456DFC",
    x"344520EC",
    x"3444D3FA",
    x"34448727",
    x"34443A71",
    x"3443EDD9",
    x"3443A15F",
    x"34435503",
    x"344308C5",
    x"3442BCA4",
    x"344270A1",
    x"344224BC",
    x"3441D8F4",
    x"34418D4B",
    x"344141BE",
    x"3440F64F",
    x"3440AAFE",
    x"34405FCA",
    x"344014B3",
    x"343FC9B9",
    x"343F7EDD",
    x"343F341E",
    x"343EE97C",
    x"343E9EF8",
    x"343E5490",
    x"343E0A46",
    x"343DC018",
    x"343D7608",
    x"343D2C14",
    x"343CE23D",
    x"343C9883",
    x"343C4EE6",
    x"343C0566",
    x"343BBC02",
    x"343B72BB",
    x"343B2990",
    x"343AE082",
    x"343A9791",
    x"343A4EBC",
    x"343A0603",
    x"3439BD67",
    x"343974E7",
    x"34392C84",
    x"3438E43C",
    x"34389C11",
    x"34385402",
    x"34380C10",
    x"3437C439",
    x"34377C7E",
    x"343734E0",
    x"3436ED5D",
    x"3436A5F6",
    x"34365EAB",
    x"3436177C",
    x"3435D069",
    x"34358972",
    x"34354296",
    x"3434FBD5",
    x"3434B531",
    x"34346EA8",
    x"3434283A",
    x"3433E1E8",
    x"34339BB2",
    x"34335597",
    x"34330F97",
    x"3432C9B3",
    x"343283E9",
    x"34323E3C",
    x"3431F8A9",
    x"3431B331",
    x"34316DD5",
    x"34312893",
    x"3430E36D",
    x"34309E62",
    x"34305971",
    x"3430149C",
    x"342FCFE1",
    x"342F8B41",
    x"342F46BC",
    x"342F0252",
    x"342EBE03",
    x"342E79CE",
    x"342E35B3",
    x"342DF1B4",
    x"342DADCF",
    x"342D6A04",
    x"342D2654",
    x"342CE2BE",
    x"342C9F43",
    x"342C5BE2",
    x"342C189B",
    x"342BD56E",
    x"342B925C",
    x"342B4F64",
    x"342B0C86",
    x"342AC9C2",
    x"342A8718",
    x"342A4489",
    x"342A0213",
    x"3429BFB7",
    x"34297D75",
    x"34293B4D",
    x"3428F93F",
    x"3428B74A",
    x"3428756F",
    x"342833AE",
    x"3427F207",
    x"3427B079",
    x"34276F05",
    x"34272DAB",
    x"3426EC6A",
    x"3426AB42",
    x"34266A34",
    x"3426293F",
    x"3425E863",
    x"3425A7A1",
    x"342566F8",
    x"34252669",
    x"3424E5F2",
    x"3424A595",
    x"34246551",
    x"34242526",
    x"3423E514",
    x"3423A51B",
    x"3423653B",
    x"34232574",
    x"3422E5C6",
    x"3422A630",
    x"342266B4",
    x"34222750",
    x"3421E805",
    x"3421A8D3",
    x"342169B9",
    x"34212AB8",
    x"3420EBD0",
    x"3420AD00",
    x"34206E49",
    x"34202FAA",
    x"341FF124",
    x"341FB2B6",
    x"341F7460",
    x"341F3623",
    x"341EF7FE",
    x"341EB9F1",
    x"341E7BFC",
    x"341E3E20",
    x"341E005C",
    x"341DC2B0",
    x"341D851C",
    x"341D47A0",
    x"341D0A3C",
    x"341CCCF0",
    x"341C8FBC",
    x"341C529F",
    x"341C159B",
    x"341BD8AE",
    x"341B9BDA",
    x"341B5F1D",
    x"341B2277",
    x"341AE5EA",
    x"341AA974",
    x"341A6D15",
    x"341A30CF",
    x"3419F49F",
    x"3419B887",
    x"34197C87",
    x"3419409E",
    x"341904CD",
    x"3418C912",
    x"34188D6F",
    x"341851E4",
    x"3418166F",
    x"3417DB12",
    x"34179FCC",
    x"3417649D",
    x"34172986",
    x"3416EE85",
    x"3416B39B",
    x"341678C9",
    x"34163E0D",
    x"34160368",
    x"3415C8DA",
    x"34158E63",
    x"34155403",
    x"341519BA",
    x"3414DF87",
    x"3414A56B",
    x"34146B66",
    x"34143177",
    x"3413F79F",
    x"3413BDDE",
    x"34138433",
    x"34134A9E",
    x"34131120",
    x"3412D7B9",
    x"34129E68",
    x"3412652D",
    x"34122C09",
    x"3411F2FB",
    x"3411BA03",
    x"34118121",
    x"34114856",
    x"34110FA1",
    x"3410D702",
    x"34109E79",
    x"34106606",
    x"34102DA9",
    x"340FF562",
    x"340FBD31",
    x"340F8516",
    x"340F4D11",
    x"340F1522",
    x"340EDD49",
    x"340EA585",
    x"340E6DD8",
    x"340E3640",
    x"340DFEBD",
    x"340DC751",
    x"340D8FF9",
    x"340D58B8",
    x"340D218C",
    x"340CEA76",
    x"340CB375",
    x"340C7C8A",
    x"340C45B4",
    x"340C0EF3",
    x"340BD848",
    x"340BA1B2",
    x"340B6B32",
    x"340B34C6",
    x"340AFE70",
    x"340AC830",
    x"340A9204",
    x"340A5BEE",
    x"340A25EC",
    x"3409F000",
    x"3409BA29",
    x"34098466",
    x"34094EB9",
    x"34091921",
    x"3408E39E",
    x"3408AE2F",
    x"340878D5",
    x"34084391",
    x"34080E61",
    x"3407D945",
    x"3407A43F",
    x"34076F4D",
    x"34073A70",
    x"340705A7",
    x"3406D0F4",
    x"34069C54",
    x"340667C9",
    x"34063353",
    x"3405FEF1",
    x"3405CAA4",
    x"3405966B",
    x"34056246",
    x"34052E36",
    x"3404FA3A",
    x"3404C653",
    x"3404927F",
    x"34045EC0",
    x"34042B15",
    x"3403F77F",
    x"3403C3FC",
    x"3403908D",
    x"34035D33",
    x"340329ED",
    x"3402F6BA",
    x"3402C39C",
    x"34029091",
    x"34025D9B",
    x"34022AB8",
    x"3401F7E9",
    x"3401C52F",
    x"34019287",
    x"34015FF4",
    x"34012D74",
    x"3400FB09",
    x"3400C8B0",
    x"3400966C",
    x"3400643B",
    x"3400321D",
    x"34000014",
    x"33FF9C3B",
    x"33FF3875",
    x"33FED4D7",
    x"33FE715F",
    x"33FE0E0E",
    x"33FDAAE4",
    x"33FD47E0",
    x"33FCE504",
    x"33FC824E",
    x"33FC1FBE",
    x"33FBBD55",
    x"33FB5B12",
    x"33FAF8F6",
    x"33FA96FF",
    x"33FA3530",
    x"33F9D386",
    x"33F97202",
    x"33F910A5",
    x"33F8AF6D",
    x"33F84E5C",
    x"33F7ED70",
    x"33F78CAA",
    x"33F72C0A",
    x"33F6CB90",
    x"33F66B3B",
    x"33F60B0C",
    x"33F5AB02",
    x"33F54B1E",
    x"33F4EB60",
    x"33F48BC6",
    x"33F42C53",
    x"33F3CD04",
    x"33F36DDA",
    x"33F30ED6",
    x"33F2AFF7",
    x"33F2513C",
    x"33F1F2A7",
    x"33F19437",
    x"33F135EB",
    x"33F0D7C5",
    x"33F079C3",
    x"33F01BE6",
    x"33EFBE2D",
    x"33EF6099",
    x"33EF032A",
    x"33EEA5DF",
    x"33EE48B8",
    x"33EDEBB6",
    x"33ED8ED8",
    x"33ED321E",
    x"33ECD589",
    x"33EC7917",
    x"33EC1CCA",
    x"33EBC0A1",
    x"33EB649B",
    x"33EB08BA",
    x"33EAACFD",
    x"33EA5163",
    x"33E9F5ED",
    x"33E99A9B",
    x"33E93F6C",
    x"33E8E461",
    x"33E8897A",
    x"33E82EB6",
    x"33E7D415",
    x"33E77998",
    x"33E71F3E",
    x"33E6C508",
    x"33E66AF4",
    x"33E61104",
    x"33E5B737",
    x"33E55D8D",
    x"33E50406",
    x"33E4AAA2",
    x"33E45161",
    x"33E3F842",
    x"33E39F47",
    x"33E3466E",
    x"33E2EDB8",
    x"33E29524",
    x"33E23CB3",
    x"33E1E465",
    x"33E18C39",
    x"33E1342F",
    x"33E0DC48",
    x"33E08483",
    x"33E02CE0",
    x"33DFD560",
    x"33DF7E02",
    x"33DF26C5",
    x"33DECFAB",
    x"33DE78B3",
    x"33DE21DD",
    x"33DDCB29",
    x"33DD7496",
    x"33DD1E26",
    x"33DCC7D7",
    x"33DC71A9",
    x"33DC1B9E",
    x"33DBC5B4",
    x"33DB6FEB",
    x"33DB1A44",
    x"33DAC4BF",
    x"33DA6F5B",
    x"33DA1A18",
    x"33D9C4F6",
    x"33D96FF6",
    x"33D91B17",
    x"33D8C659",
    x"33D871BC",
    x"33D81D40",
    x"33D7C8E5",
    x"33D774AB",
    x"33D72092",
    x"33D6CC99",
    x"33D678C2",
    x"33D6250B",
    x"33D5D175",
    x"33D57DFF",
    x"33D52AAA",
    x"33D4D776",
    x"33D48462",
    x"33D4316F",
    x"33D3DE9B",
    x"33D38BE9",
    x"33D33956",
    x"33D2E6E4",
    x"33D29492",
    x"33D24260",
    x"33D1F04E",
    x"33D19E5C",
    x"33D14C8A",
    x"33D0FAD8",
    x"33D0A946",
    x"33D057D4",
    x"33D00682",
    x"33CFB54F",
    x"33CF643C",
    x"33CF1349",
    x"33CEC275",
    x"33CE71C1",
    x"33CE212C",
    x"33CDD0B7",
    x"33CD8061",
    x"33CD302A",
    x"33CCE013",
    x"33CC901B",
    x"33CC4043",
    x"33CBF089",
    x"33CBA0EF",
    x"33CB5173",
    x"33CB0217",
    x"33CAB2DA",
    x"33CA63BB",
    x"33CA14BC",
    x"33C9C5DB",
    x"33C97719",
    x"33C92876",
    x"33C8D9F2",
    x"33C88B8C",
    x"33C83D44",
    x"33C7EF1C",
    x"33C7A112",
    x"33C75326",
    x"33C70559",
    x"33C6B7AA",
    x"33C66A19",
    x"33C61CA7",
    x"33C5CF53",
    x"33C5821D",
    x"33C53505",
    x"33C4E80B",
    x"33C49B30",
    x"33C44E72",
    x"33C401D3",
    x"33C3B551",
    x"33C368ED",
    x"33C31CA7",
    x"33C2D07E",
    x"33C28474",
    x"33C23887",
    x"33C1ECB8",
    x"33C1A106",
    x"33C15572",
    x"33C109FB",
    x"33C0BEA2",
    x"33C07366",
    x"33C02848",
    x"33BFDD47",
    x"33BF9263",
    x"33BF479C",
    x"33BEFCF3",
    x"33BEB267",
    x"33BE67F8",
    x"33BE1DA6",
    x"33BDD370",
    x"33BD8958",
    x"33BD3F5D",
    x"33BCF57F",
    x"33BCABBD",
    x"33BC6219",
    x"33BC1891",
    x"33BBCF25",
    x"33BB85D7",
    x"33BB3CA5",
    x"33BAF38F",
    x"33BAAA97",
    x"33BA61BA",
    x"33BA18FA",
    x"33B9D057",
    x"33B987CF",
    x"33B93F65",
    x"33B8F716",
    x"33B8AEE3",
    x"33B866CD",
    x"33B81ED3",
    x"33B7D6F5",
    x"33B78F33",
    x"33B7478D",
    x"33B70003",
    x"33B6B895",
    x"33B67143",
    x"33B62A0D",
    x"33B5E2F2",
    x"33B59BF3",
    x"33B55510",
    x"33B50E49",
    x"33B4C79D",
    x"33B4810D",
    x"33B43A98",
    x"33B3F43F",
    x"33B3AE01",
    x"33B367DF",
    x"33B321D8",
    x"33B2DBED",
    x"33B2961C",
    x"33B25067",
    x"33B20ACE",
    x"33B1C54F",
    x"33B17FEC",
    x"33B13AA3",
    x"33B0F576",
    x"33B0B063",
    x"33B06B6C",
    x"33B0268F",
    x"33AFE1CE",
    x"33AF9D27",
    x"33AF589B",
    x"33AF142A",
    x"33AECFD3",
    x"33AE8B97",
    x"33AE4776",
    x"33AE036F",
    x"33ADBF83",
    x"33AD7BB2",
    x"33AD37FB",
    x"33ACF45E",
    x"33ACB0DC",
    x"33AC6D74",
    x"33AC2A26",
    x"33ABE6F3",
    x"33ABA3DA",
    x"33AB60DB",
    x"33AB1DF6",
    x"33AADB2C",
    x"33AA987B",
    x"33AA55E4",
    x"33AA1368",
    x"33A9D105",
    x"33A98EBD",
    x"33A94C8E",
    x"33A90A79",
    x"33A8C87D",
    x"33A8869C",
    x"33A844D4",
    x"33A80326",
    x"33A7C192",
    x"33A78017",
    x"33A73EB6",
    x"33A6FD6E",
    x"33A6BC40",
    x"33A67B2B",
    x"33A63A30",
    x"33A5F94D",
    x"33A5B885",
    x"33A577D5",
    x"33A5373F",
    x"33A4F6C2",
    x"33A4B65E",
    x"33A47614",
    x"33A435E2",
    x"33A3F5CA",
    x"33A3B5CA",
    x"33A375E3",
    x"33A33616",
    x"33A2F661",
    x"33A2B6C5",
    x"33A27742",
    x"33A237D8",
    x"33A1F887",
    x"33A1B94E",
    x"33A17A2E",
    x"33A13B27",
    x"33A0FC38",
    x"33A0BD62",
    x"33A07EA4",
    x"33A03FFF",
    x"33A00172",
    x"339FC2FD",
    x"339F84A1",
    x"339F465E",
    x"339F0832",
    x"339ECA1F",
    x"339E8C25",
    x"339E4E42",
    x"339E1077",
    x"339DD2C5",
    x"339D952B",
    x"339D57A8",
    x"339D1A3E",
    x"339CDCEC",
    x"339C9FB2",
    x"339C628F",
    x"339C2585",
    x"339BE892",
    x"339BABB7",
    x"339B6EF4",
    x"339B3248",
    x"339AF5B4",
    x"339AB938",
    x"339A7CD4",
    x"339A4087",
    x"339A0451",
    x"3399C833",
    x"33998C2D",
    x"3399503E",
    x"33991466",
    x"3398D8A6",
    x"33989CFD",
    x"3398616B",
    x"339825F1",
    x"3397EA8E",
    x"3397AF41",
    x"3397740D",
    x"339738EF",
    x"3396FDE8",
    x"3396C2F8",
    x"33968820",
    x"33964D5E",
    x"339612B3",
    x"3395D81F",
    x"33959DA2",
    x"3395633C",
    x"339528ED",
    x"3394EEB4",
    x"3394B492",
    x"33947A87",
    x"33944093",
    x"339406B5",
    x"3393CCED",
    x"3393933D",
    x"339359A2",
    x"3393201F",
    x"3392E6B1",
    x"3392AD5A",
    x"3392741A",
    x"33923AF0",
    x"339201DC",
    x"3391C8DE",
    x"33918FF7",
    x"33915726",
    x"33911E6B",
    x"3390E5C6",
    x"3390AD37",
    x"339074BF",
    x"33903C5C",
    x"3390040F",
    x"338FCBD9",
    x"338F93B8",
    x"338F5BAD",
    x"338F23B9",
    x"338EEBDA",
    x"338EB410",
    x"338E7C5D",
    x"338E44BF",
    x"338E0D37",
    x"338DD5C5",
    x"338D9E68",
    x"338D6721",
    x"338D2FF0",
    x"338CF8D4",
    x"338CC1CD",
    x"338C8ADC",
    x"338C5401",
    x"338C1D3A",
    x"338BE68A",
    x"338BAFEE",
    x"338B7968",
    x"338B42F8",
    x"338B0C9C",
    x"338AD656",
    x"338AA025",
    x"338A6A09",
    x"338A3402",
    x"3389FE10",
    x"3389C833",
    x"3389926B",
    x"33895CB9",
    x"3389271B",
    x"3388F192",
    x"3388BC1E",
    x"338886BF",
    x"33885175",
    x"33881C40",
    x"3387E71F",
    x"3387B213",
    x"33877D1C",
    x"33874839",
    x"3387136B",
    x"3386DEB2",
    x"3386AA0D",
    x"3386757D",
    x"33864102",
    x"33860C9A",
    x"3385D848",
    x"3385A409",
    x"33856FE0",
    x"33853BCA",
    x"338507C9",
    x"3384D3DC",
    x"3384A003",
    x"33846C3F",
    x"3384388F",
    x"338404F3",
    x"3383D16B",
    x"33839DF7",
    x"33836A97",
    x"3383374C",
    x"33830414",
    x"3382D0F1",
    x"33829DE1",
    x"33826AE5",
    x"338237FD",
    x"3382052A",
    x"3381D269",
    x"33819FBD",
    x"33816D25",
    x"33813AA0",
    x"3381082F",
    x"3380D5D1",
    x"3380A388",
    x"33807152",
    x"33803F2F",
    x"33800D20",
    x"337FB64A",
    x"337F527A",
    x"337EEED1",
    x"337E8B50",
    x"337E27F5",
    x"337DC4C0",
    x"337D61B3",
    x"337CFECC",
    x"337C9C0C",
    x"337C3972",
    x"337BD6FF",
    x"337B74B2",
    x"337B128C",
    x"337AB08C",
    x"337A4EB2",
    x"3379ECFE",
    x"33798B71",
    x"33792A09",
    x"3378C8C8",
    x"337867AC",
    x"337806B7",
    x"3377A5E7",
    x"3377453D",
    x"3376E4B9",
    x"3376845A",
    x"33762421",
    x"3375C40E",
    x"33756420",
    x"33750458",
    x"3374A4B5",
    x"33744537",
    x"3373E5DF",
    x"337386AC",
    x"3373279D",
    x"3372C8B5",
    x"337269F1",
    x"33720B52",
    x"3371ACD8",
    x"33714E83",
    x"3370F052",
    x"33709247",
    x"33703460",
    x"336FD69E",
    x"336F7900",
    x"336F1B87",
    x"336EBE33",
    x"336E6103",
    x"336E03F7",
    x"336DA710",
    x"336D4A4D",
    x"336CEDAE",
    x"336C9133",
    x"336C34DC",
    x"336BD8AA",
    x"336B7C9B",
    x"336B20B0",
    x"336AC4E9",
    x"336A6946",
    x"336A0DC7",
    x"3369B26C",
    x"33695734",
    x"3368FC1F",
    x"3368A12F",
    x"33684661",
    x"3367EBB8",
    x"33679131",
    x"336736CE",
    x"3366DC8E",
    x"33668272",
    x"33662879",
    x"3365CEA2",
    x"336574EF",
    x"33651B5F",
    x"3364C1F2",
    x"336468A7",
    x"33640F80",
    x"3363B67B",
    x"33635D99",
    x"336304DA",
    x"3362AC3E",
    x"336253C4",
    x"3361FB6C",
    x"3361A337",
    x"33614B25",
    x"3360F334",
    x"33609B67",
    x"336043BB",
    x"335FEC32",
    x"335F94CA",
    x"335F3D85",
    x"335EE662",
    x"335E8F61",
    x"335E3882",
    x"335DE1C5",
    x"335D8B2A",
    x"335D34B0",
    x"335CDE59",
    x"335C8823",
    x"335C320E",
    x"335BDC1C",
    x"335B864A",
    x"335B309B",
    x"335ADB0C",
    x"335A859F",
    x"335A3054",
    x"3359DB2A",
    x"33598621",
    x"33593139",
    x"3358DC72",
    x"335887CD",
    x"33583348",
    x"3357DEE5",
    x"33578AA2",
    x"33573680",
    x"3356E27F",
    x"33568E9F",
    x"33563AE0",
    x"3355E741",
    x"335593C3",
    x"33554066",
    x"3354ED29",
    x"33549A0D",
    x"33544711",
    x"3353F435",
    x"3353A17A",
    x"33534EDF",
    x"3352FC64",
    x"3352AA0A",
    x"335257CF",
    x"335205B5",
    x"3351B3BB",
    x"335161E1",
    x"33511026",
    x"3350BE8C",
    x"33506D11",
    x"33501BB7",
    x"334FCA7C",
    x"334F7961",
    x"334F2865",
    x"334ED789",
    x"334E86CD",
    x"334E3630",
    x"334DE5B2",
    x"334D9554",
    x"334D4516",
    x"334CF4F6",
    x"334CA4F6",
    x"334C5515",
    x"334C0554",
    x"334BB5B1",
    x"334B662E",
    x"334B16C9",
    x"334AC784",
    x"334A785D",
    x"334A2956",
    x"3349DA6D",
    x"33498BA3",
    x"33493CF8",
    x"3348EE6B",
    x"33489FFE",
    x"334851AE",
    x"3348037E",
    x"3347B56C",
    x"33476778",
    x"334719A3",
    x"3346CBEC",
    x"33467E54",
    x"334630D9",
    x"3345E37D",
    x"33459640",
    x"33454920",
    x"3344FC1E",
    x"3344AF3B",
    x"33446276",
    x"334415CE",
    x"3343C944",
    x"33437CD9",
    x"3343308B",
    x"3342E45B",
    x"33429849",
    x"33424C54",
    x"3342007D",
    x"3341B4C3",
    x"33416928",
    x"33411DA9",
    x"3340D248",
    x"33408705",
    x"33403BDF",
    x"333FF0D6",
    x"333FA5EB",
    x"333F5B1D",
    x"333F106C",
    x"333EC5D8",
    x"333E7B61",
    x"333E3107",
    x"333DE6CB",
    x"333D9CAB",
    x"333D52A8",
    x"333D08C2",
    x"333CBEF9",
    x"333C754D",
    x"333C2BBE",
    x"333BE24B",
    x"333B98F5",
    x"333B4FBC",
    x"333B069F",
    x"333ABD9E",
    x"333A74BA",
    x"333A2BF3",
    x"3339E348",
    x"33399ABA",
    x"33395247",
    x"333909F1",
    x"3338C1B7",
    x"3338799A",
    x"33383198",
    x"3337E9B3",
    x"3337A1EA",
    x"33375A3D",
    x"333712AB",
    x"3336CB36",
    x"333683DD",
    x"33363C9F",
    x"3335F57D",
    x"3335AE77",
    x"3335678D",
    x"333520BE",
    x"3334DA0B",
    x"33349374",
    x"33344CF8",
    x"33340698",
    x"3333C053",
    x"33337A2A",
    x"3333341B",
    x"3332EE29",
    x"3332A851",
    x"33326295",
    x"33321CF4",
    x"3331D76F",
    x"33319204",
    x"33314CB5",
    x"33310780",
    x"3330C267",
    x"33307D68",
    x"33303885",
    x"332FF3BC",
    x"332FAF0E",
    x"332F6A7B",
    x"332F2603",
    x"332EE1A6",
    x"332E9D63",
    x"332E593B",
    x"332E152D",
    x"332DD13A",
    x"332D8D62",
    x"332D49A4",
    x"332D0600",
    x"332CC277",
    x"332C7F08",
    x"332C3BB4",
    x"332BF879",
    x"332BB559",
    x"332B7254",
    x"332B2F68",
    x"332AEC97",
    x"332AA9DF",
    x"332A6742",
    x"332A24BF",
    x"3329E255",
    x"3329A006",
    x"33295DD0",
    x"33291BB4",
    x"3328D9B3",
    x"332897CA",
    x"332855FC",
    x"33281447",
    x"3327D2AC",
    x"3327912B",
    x"33274FC3",
    x"33270E74",
    x"3326CD3F",
    x"33268C24",
    x"33264B22",
    x"33260A39",
    x"3325C96A",
    x"332588B4",
    x"33254817",
    x"33250793",
    x"3324C729",
    x"332486D8",
    x"332446A0",
    x"33240681",
    x"3323C67B",
    x"3323868E",
    x"332346BA",
    x"332306FE",
    x"3322C75C",
    x"332287D3",
    x"33224862",
    x"3322090A",
    x"3321C9CB",
    x"33218AA4",
    x"33214B97",
    x"33210CA1",
    x"3320CDC5",
    x"33208F01",
    x"33205055",
    x"332011C2",
    x"331FD347",
    x"331F94E5",
    x"331F569B",
    x"331F1869",
    x"331EDA50",
    x"331E9C4E",
    x"331E5E65",
    x"331E2095",
    x"331DE2DC",
    x"331DA53B",
    x"331D67B3",
    x"331D2A42",
    x"331CECEA",
    x"331CAFA9",
    x"331C7281",
    x"331C3570",
    x"331BF877",
    x"331BBB96",
    x"331B7ECC",
    x"331B421B",
    x"331B0581",
    x"331AC8FE",
    x"331A8C94",
    x"331A5041",
    x"331A1405",
    x"3319D7E1",
    x"33199BD4",
    x"33195FDF",
    x"33192401",
    x"3318E83B",
    x"3318AC8C",
    x"331870F4",
    x"33183574",
    x"3317FA0A",
    x"3317BEB8",
    x"3317837D",
    x"3317485A",
    x"33170D4D",
    x"3316D257",
    x"33169778",
    x"33165CB1",
    x"33162200",
    x"3315E766",
    x"3315ACE3",
    x"33157277",
    x"33153822",
    x"3314FDE3",
    x"3314C3BB",
    x"331489AA",
    x"33144FB0",
    x"331415CC",
    x"3313DBFF",
    x"3313A248",
    x"331368A8",
    x"33132F1E",
    x"3312F5AB",
    x"3312BC4E",
    x"33128308",
    x"331249D8",
    x"331210BE",
    x"3311D7BB",
    x"33119ECE",
    x"331165F7",
    x"33112D36",
    x"3310F48C",
    x"3310BBF7",
    x"33108379",
    x"33104B10",
    x"331012BE",
    x"330FDA82",
    x"330FA25B",
    x"330F6A4B",
    x"330F3250",
    x"330EFA6C",
    x"330EC29D",
    x"330E8AE4",
    x"330E5340",
    x"330E1BB2",
    x"330DE43A",
    x"330DACD8",
    x"330D758B",
    x"330D3E54",
    x"330D0733",
    x"330CD027",
    x"330C9930",
    x"330C624F",
    x"330C2B83",
    x"330BF4CD",
    x"330BBE2C",
    x"330B87A0",
    x"330B512A",
    x"330B1AC9",
    x"330AE47D",
    x"330AAE46",
    x"330A7825",
    x"330A4219",
    x"330A0C21",
    x"3309D63F",
    x"3309A072",
    x"33096ABA",
    x"33093517",
    x"3308FF88",
    x"3308CA0F",
    x"330894AA",
    x"33085F5B",
    x"33082A20",
    x"3307F4FA",
    x"3307BFE8",
    x"33078AEC",
    x"33075604",
    x"33072131",
    x"3306EC72",
    x"3306B7C8",
    x"33068332",
    x"33064EB1",
    x"33061A45",
    x"3305E5ED",
    x"3305B1A9",
    x"33057D7A",
    x"3305495F",
    x"33051559",
    x"3304E167",
    x"3304AD89",
    x"330479BF",
    x"3304460A",
    x"33041268",
    x"3303DEDB",
    x"3303AB62",
    x"330377FD",
    x"330344AC",
    x"33031170",
    x"3302DE47",
    x"3302AB32",
    x"33027831",
    x"33024544",
    x"3302126B",
    x"3301DFA6",
    x"3301ACF4",
    x"33017A56",
    x"330147CD",
    x"33011556",
    x"3300E2F4",
    x"3300B0A5",
    x"33007E6A",
    x"33004C42",
    x"33001A2E",
    x"32FFD05C",
    x"32FF6C82",
    x"32FF08CF",
    x"32FEA543",
    x"32FE41DE",
    x"32FDDE9F",
    x"32FD7B88",
    x"32FD1897",
    x"32FCB5CD",
    x"32FC5329",
    x"32FBF0AC",
    x"32FB8E55",
    x"32FB2C24",
    x"32FACA1A",
    x"32FA6836",
    x"32FA0679",
    x"32F9A4E1",
    x"32F94370",
    x"32F8E225",
    x"32F880FF",
    x"32F82000",
    x"32F7BF26",
    x"32F75E72",
    x"32F6FDE4",
    x"32F69D7C",
    x"32F63D39",
    x"32F5DD1C",
    x"32F57D25",
    x"32F51D52",
    x"32F4BDA6",
    x"32F45E1E",
    x"32F3FEBC",
    x"32F39F7F",
    x"32F34068",
    x"32F2E175",
    x"32F282A7",
    x"32F223FF",
    x"32F1C57B",
    x"32F1671D",
    x"32F108E3",
    x"32F0AACE",
    x"32F04CDD",
    x"32EFEF12",
    x"32EF916A",
    x"32EF33E8",
    x"32EED68A",
    x"32EE7950",
    x"32EE1C3B",
    x"32EDBF4A",
    x"32ED627E",
    x"32ED05D5",
    x"32ECA951",
    x"32EC4CF1",
    x"32EBF0B5",
    x"32EB949D",
    x"32EB38A9",
    x"32EADCD9",
    x"32EA812C",
    x"32EA25A4",
    x"32E9CA3F",
    x"32E96EFE",
    x"32E913E0",
    x"32E8B8E6",
    x"32E85E10",
    x"32E8035D",
    x"32E7A8CD",
    x"32E74E61",
    x"32E6F418",
    x"32E699F2",
    x"32E63FEF",
    x"32E5E610",
    x"32E58C54",
    x"32E532BA",
    x"32E4D944",
    x"32E47FF1",
    x"32E426C0",
    x"32E3CDB2",
    x"32E374C7",
    x"32E31BFF",
    x"32E2C359",
    x"32E26AD6",
    x"32E21276",
    x"32E1BA38",
    x"32E1621C",
    x"32E10A23",
    x"32E0B24D",
    x"32E05A98",
    x"32E00306",
    x"32DFAB96",
    x"32DF5448",
    x"32DEFD1C",
    x"32DEA612",
    x"32DE4F2A",
    x"32DDF864",
    x"32DDA1C0",
    x"32DD4B3E",
    x"32DCF4DD",
    x"32DC9E9E",
    x"32DC4881",
    x"32DBF286",
    x"32DB9CAC",
    x"32DB46F3",
    x"32DAF15C",
    x"32DA9BE7",
    x"32DA4692",
    x"32D9F160",
    x"32D99C4E",
    x"32D9475D",
    x"32D8F28E",
    x"32D89DE0",
    x"32D84953",
    x"32D7F4E7",
    x"32D7A09B",
    x"32D74C71",
    x"32D6F868",
    x"32D6A47F",
    x"32D650B7",
    x"32D5FD10",
    x"32D5A989",
    x"32D55623",
    x"32D502DE",
    x"32D4AFB9",
    x"32D45CB5",
    x"32D409D1",
    x"32D3B70D",
    x"32D3646A",
    x"32D311E7",
    x"32D2BF84",
    x"32D26D41",
    x"32D21B1E",
    x"32D1C91C",
    x"32D17739",
    x"32D12577",
    x"32D0D3D4",
    x"32D08251",
    x"32D030EE",
    x"32CFDFAB",
    x"32CF8E87",
    x"32CF3D84",
    x"32CEEC9F",
    x"32CE9BDB",
    x"32CE4B36",
    x"32CDFAB0",
    x"32CDAA4A",
    x"32CD5A03",
    x"32CD09DB",
    x"32CCB9D3",
    x"32CC69EA",
    x"32CC1A20",
    x"32CBCA76",
    x"32CB7AEA",
    x"32CB2B7E",
    x"32CADC30",
    x"32CA8D02",
    x"32CA3DF2",
    x"32C9EF01",
    x"32C9A02F",
    x"32C9517C",
    x"32C902E8",
    x"32C8B472",
    x"32C8661B",
    x"32C817E2",
    x"32C7C9C8",
    x"32C77BCC",
    x"32C72DEF",
    x"32C6E030",
    x"32C69290",
    x"32C6450E",
    x"32C5F7AA",
    x"32C5AA64",
    x"32C55D3D",
    x"32C51034",
    x"32C4C348",
    x"32C4767B",
    x"32C429CC",
    x"32C3DD3A",
    x"32C390C7",
    x"32C34471",
    x"32C2F839",
    x"32C2AC1F",
    x"32C26023",
    x"32C21444",
    x"32C1C883",
    x"32C17CDF",
    x"32C13159",
    x"32C0E5F1",
    x"32C09AA6",
    x"32C04F78",
    x"32C00468",
    x"32BFB975",
    x"32BF6E9F",
    x"32BF23E6",
    x"32BED94B",
    x"32BE8ECC",
    x"32BE446B",
    x"32BDFA27",
    x"32BDB000",
    x"32BD65F5",
    x"32BD1C08",
    x"32BCD237",
    x"32BC8884",
    x"32BC3EED",
    x"32BBF573",
    x"32BBAC15",
    x"32BB62D4",
    x"32BB19B0",
    x"32BAD0A8",
    x"32BA87BD",
    x"32BA3EEE",
    x"32B9F63C",
    x"32B9ADA6",
    x"32B9652C",
    x"32B91CCF",
    x"32B8D48D",
    x"32B88C68",
    x"32B84460",
    x"32B7FC73",
    x"32B7B4A2",
    x"32B76CEE",
    x"32B72555",
    x"32B6DDD9",
    x"32B69678",
    x"32B64F33",
    x"32B6080A",
    x"32B5C0FD",
    x"32B57A0B",
    x"32B53336",
    x"32B4EC7B",
    x"32B4A5DD",
    x"32B45F5A",
    x"32B418F2",
    x"32B3D2A6",
    x"32B38C76",
    x"32B34660",
    x"32B30067",
    x"32B2BA88",
    x"32B274C5",
    x"32B22F1D",
    x"32B1E990",
    x"32B1A41E",
    x"32B15EC8",
    x"32B1198C",
    x"32B0D46C",
    x"32B08F66",
    x"32B04A7C",
    x"32B005AC",
    x"32AFC0F7",
    x"32AF7C5D",
    x"32AF37DE",
    x"32AEF37A",
    x"32AEAF30",
    x"32AE6B01",
    x"32AE26EC",
    x"32ADE2F2",
    x"32AD9F13",
    x"32AD5B4E",
    x"32AD17A4",
    x"32ACD414",
    x"32AC909E",
    x"32AC4D43",
    x"32AC0A02",
    x"32ABC6DB",
    x"32AB83CE",
    x"32AB40DC",
    x"32AAFE04",
    x"32AABB45",
    x"32AA78A1",
    x"32AA3617",
    x"32A9F3A7",
    x"32A9B151",
    x"32A96F14",
    x"32A92CF2",
    x"32A8EAE9",
    x"32A8A8FA",
    x"32A86725",
    x"32A8256A",
    x"32A7E3C8",
    x"32A7A240",
    x"32A760D1",
    x"32A71F7C",
    x"32A6DE41",
    x"32A69D1F",
    x"32A65C16",
    x"32A61B27",
    x"32A5DA51",
    x"32A59994",
    x"32A558F1",
    x"32A51867",
    x"32A4D7F6",
    x"32A4979E",
    x"32A4575F",
    x"32A4173A",
    x"32A3D72D",
    x"32A39739",
    x"32A3575F",
    x"32A3179D",
    x"32A2D7F4",
    x"32A29864",
    x"32A258ED",
    x"32A2198F",
    x"32A1DA49",
    x"32A19B1C",
    x"32A15C08",
    x"32A11D0C",
    x"32A0DE29",
    x"32A09F5F",
    x"32A060AD",
    x"32A02213",
    x"329FE392",
    x"329FA52A",
    x"329F66D9",
    x"329F28A1",
    x"329EEA81",
    x"329EAC7A",
    x"329E6E8B",
    x"329E30B4",
    x"329DF2F5",
    x"329DB54E",
    x"329D77BF",
    x"329D3A48",
    x"329CFCE9",
    x"329CBFA3",
    x"329C8274",
    x"329C455D",
    x"329C085E",
    x"329BCB76",
    x"329B8EA7",
    x"329B51EF",
    x"329B154F",
    x"329AD8C6",
    x"329A9C55",
    x"329A5FFC",
    x"329A23BA",
    x"3299E790",
    x"3299AB7D",
    x"32996F82",
    x"3299339E",
    x"3298F7D2",
    x"3298BC1D",
    x"3298807F",
    x"329844F8",
    x"32980989",
    x"3297CE31",
    x"329792F0",
    x"329757C6",
    x"32971CB3",
    x"3296E1B7",
    x"3296A6D3",
    x"32966C05",
    x"3296314E",
    x"3295F6AF",
    x"3295BC26",
    x"329581B4",
    x"32954758",
    x"32950D14",
    x"3294D2E6",
    x"329498CF",
    x"32945ECF",
    x"329424E5",
    x"3293EB12",
    x"3293B155",
    x"329377AF",
    x"32933E20",
    x"329304A7",
    x"3292CB44",
    x"329291F8",
    x"329258C2",
    x"32921FA3",
    x"3291E699",
    x"3291ADA6",
    x"329174CA",
    x"32913C03",
    x"32910353",
    x"3290CAB9",
    x"32909234",
    x"329059C6",
    x"3290216E",
    x"328FE92C",
    x"328FB100",
    x"328F78EA",
    x"328F40EA",
    x"328F08FF",
    x"328ED12B",
    x"328E996C",
    x"328E61C3",
    x"328E2A2F",
    x"328DF2B2",
    x"328DBB4A",
    x"328D83F7",
    x"328D4CBB",
    x"328D1593",
    x"328CDE82",
    x"328CA786",
    x"328C709F",
    x"328C39CE",
    x"328C0312",
    x"328BCC6B",
    x"328B95DA",
    x"328B5F5E",
    x"328B28F7",
    x"328AF2A6",
    x"328ABC6A",
    x"328A8643",
    x"328A5031",
    x"328A1A34",
    x"3289E44C",
    x"3289AE7A",
    x"328978BC",
    x"32894313",
    x"32890D80",
    x"3288D801",
    x"3288A297",
    x"32886D42",
    x"32883802",
    x"328802D6",
    x"3287CDBF",
    x"328798BD",
    x"328763D0",
    x"32872EF7",
    x"3286FA33",
    x"3286C584",
    x"328690E9",
    x"32865C63",
    x"328627F1",
    x"3285F393",
    x"3285BF4B",
    x"32858B16",
    x"328556F6",
    x"328522EA",
    x"3284EEF3",
    x"3284BB0F",
    x"32848740",
    x"32845386",
    x"32841FDF",
    x"3283EC4D",
    x"3283B8CF",
    x"32838564",
    x"3283520E",
    x"32831ECC",
    x"3282EB9E",
    x"3282B884",
    x"3282857E",
    x"3282528C",
    x"32821FAE",
    x"3281ECE3",
    x"3281BA2D",
    x"3281878A",
    x"328154FB",
    x"3281227F",
    x"3280F018",
    x"3280BDC4",
    x"32808B83",
    x"32805957",
    x"3280273E",
    x"327FEA70",
    x"327F868C",
    x"327F22CF",
    x"327EBF39",
    x"327E5BCA",
    x"327DF881",
    x"327D955F",
    x"327D3264",
    x"327CCF90",
    x"327C6CE2",
    x"327C0A5B",
    x"327BA7FA",
    x"327B45C0",
    x"327AE3AC",
    x"327A81BE",
    x"327A1FF6",
    x"3279BE55",
    x"32795CD9",
    x"3278FB84",
    x"32789A55",
    x"3278394C",
    x"3277D868",
    x"327777AB",
    x"32771713",
    x"3276B6A0",
    x"32765654",
    x"3275F62D",
    x"3275962C",
    x"32753650",
    x"3274D699",
    x"32747708",
    x"3274179C",
    x"3273B856",
    x"32735934",
    x"3272FA38",
    x"32729B61",
    x"32723CAE",
    x"3271DE21",
    x"32717FB9",
    x"32712175",
    x"3270C357",
    x"3270655D",
    x"32700788",
    x"326FA9D7",
    x"326F4C4B",
    x"326EEEE3",
    x"326E91A0",
    x"326E3481",
    x"326DD787",
    x"326D7AB1",
    x"326D1DFF",
    x"326CC172",
    x"326C6508",
    x"326C08C3",
    x"326BACA1",
    x"326B50A4",
    x"326AF4CA",
    x"326A9915",
    x"326A3D83",
    x"3269E214",
    x"326986CA",
    x"32692BA3",
    x"3268D0A0",
    x"326875C0",
    x"32681B04",
    x"3267C06B",
    x"326765F5",
    x"32670BA3",
    x"3266B174",
    x"32665769",
    x"3265FD80",
    x"3265A3BB",
    x"32654A18",
    x"3264F099",
    x"3264973C",
    x"32643E03",
    x"3263E4EC",
    x"32638BF8",
    x"32633326",
    x"3262DA78",
    x"326281EC",
    x"32622982",
    x"3261D13B",
    x"32617917",
    x"32612115",
    x"3260C935",
    x"32607177",
    x"326019DC",
    x"325FC263",
    x"325F6B0C",
    x"325F13D7",
    x"325EBCC5",
    x"325E65D4",
    x"325E0F05",
    x"325DB858",
    x"325D61CD",
    x"325D0B64",
    x"325CB51C",
    x"325C5EF6",
    x"325C08F2",
    x"325BB30F",
    x"325B5D4E",
    x"325B07AE",
    x"325AB230",
    x"325A5CD3",
    x"325A0798",
    x"3259B27D",
    x"32595D84",
    x"325908AC",
    x"3258B3F5",
    x"32585F60",
    x"32580AEB",
    x"3257B697",
    x"32576264",
    x"32570E52",
    x"3256BA61",
    x"32566690",
    x"325612E1",
    x"3255BF52",
    x"32556BE3",
    x"32551895",
    x"3254C568",
    x"3254725B",
    x"32541F6F",
    x"3253CCA3",
    x"325379F7",
    x"3253276B",
    x"3252D500",
    x"325282B5",
    x"3252308A",
    x"3251DE7F",
    x"32518C94",
    x"32513AC9",
    x"3250E91E",
    x"32509793",
    x"32504628",
    x"324FF4DC",
    x"324FA3B0",
    x"324F52A4",
    x"324F01B8",
    x"324EB0EB",
    x"324E603E",
    x"324E0FB0",
    x"324DBF41",
    x"324D6EF2",
    x"324D1EC3",
    x"324CCEB2",
    x"324C7EC1",
    x"324C2EEF",
    x"324BDF3C",
    x"324B8FA9",
    x"324B4034",
    x"324AF0DF",
    x"324AA1A8",
    x"324A5290",
    x"324A0397",
    x"3249B4BD",
    x"32496602",
    x"32491766",
    x"3248C8E8",
    x"32487A89",
    x"32482C48",
    x"3247DE26",
    x"32479023",
    x"3247423E",
    x"3246F477",
    x"3246A6CF",
    x"32465944",
    x"32460BD9",
    x"3245BE8B",
    x"3245715C",
    x"3245244B",
    x"3244D758",
    x"32448A82",
    x"32443DCB",
    x"3243F132",
    x"3243A4B7",
    x"32435859",
    x"32430C1A",
    x"3242BFF8",
    x"324273F4",
    x"3242280D",
    x"3241DC44",
    x"32419099",
    x"3241450C",
    x"3240F99B",
    x"3240AE48",
    x"32406313",
    x"324017FB",
    x"323FCD00",
    x"323F8223",
    x"323F3763",
    x"323EECC0",
    x"323EA23A",
    x"323E57D1",
    x"323E0D85",
    x"323DC356",
    x"323D7944",
    x"323D2F50",
    x"323CE577",
    x"323C9BBC",
    x"323C521E",
    x"323C089C",
    x"323BBF37",
    x"323B75EF",
    x"323B2CC3",
    x"323AE3B4",
    x"323A9AC1",
    x"323A51EB",
    x"323A0931",
    x"3239C094",
    x"32397813",
    x"32392FAE",
    x"3238E765",
    x"32389F39",
    x"32385729",
    x"32380F35",
    x"3237C75D",
    x"32377FA1",
    x"32373801",
    x"3236F07D",
    x"3236A915",
    x"323661C9",
    x"32361A99",
    x"3235D384",
    x"32358C8C",
    x"323545AF",
    x"3234FEED",
    x"3234B847",
    x"323471BD",
    x"32342B4F",
    x"3233E4FB",
    x"32339EC4",
    x"323358A7",
    x"323312A6",
    x"3232CCC1",
    x"323286F6",
    x"32324147",
    x"3231FBB3",
    x"3231B63B",
    x"323170DD",
    x"32312B9A",
    x"3230E673",
    x"3230A166",
    x"32305C75",
    x"3230179E",
    x"322FD2E2",
    x"322F8E41",
    x"322F49BB",
    x"322F0550",
    x"322EC0FF",
    x"322E7CC9",
    x"322E38AE",
    x"322DF4AD",
    x"322DB0C6",
    x"322D6CFB",
    x"322D2949",
    x"322CE5B2",
    x"322CA236",
    x"322C5ED4",
    x"322C1B8C",
    x"322BD85E",
    x"322B954B",
    x"322B5251",
    x"322B0F72",
    x"322ACCAD",
    x"322A8A02",
    x"322A4771",
    x"322A04FB",
    x"3229C29E",
    x"3229805A",
    x"32293E31",
    x"3228FC22",
    x"3228BA2C",
    x"32287850",
    x"3228368E",
    x"3227F4E6",
    x"3227B357",
    x"322771E2",
    x"32273086",
    x"3226EF44",
    x"3226AE1B",
    x"32266D0C",
    x"32262C16",
    x"3225EB39",
    x"3225AA76",
    x"322569CC",
    x"3225293B",
    x"3224E8C4",
    x"3224A865",
    x"32246820",
    x"322427F4",
    x"3223E7E1",
    x"3223A7E7",
    x"32236806",
    x"3223283E",
    x"3222E88E",
    x"3222A8F8",
    x"3222697A",
    x"32222A16",
    x"3221EACA",
    x"3221AB96",
    x"32216C7B",
    x"32212D79",
    x"3220EE90",
    x"3220AFBF",
    x"32207107",
    x"32203267",
    x"321FF3DF",
    x"321FB570",
    x"321F7719",
    x"321F38DB",
    x"321EFAB5",
    x"321EBCA7",
    x"321E7EB2",
    x"321E40D4",
    x"321E030F",
    x"321DC562",
    x"321D87CD",
    x"321D4A50",
    x"321D0CEB",
    x"321CCF9E",
    x"321C9268",
    x"321C554B",
    x"321C1846",
    x"321BDB58",
    x"321B9E82",
    x"321B61C4",
    x"321B251E",
    x"321AE88F",
    x"321AAC18",
    x"321A6FB9",
    x"321A3371",
    x"3219F741",
    x"3219BB28",
    x"32197F26",
    x"3219433D",
    x"3219076A",
    x"3218CBAF",
    x"3218900B",
    x"3218547E",
    x"32181909",
    x"3217DDAB",
    x"3217A264",
    x"32176734",
    x"32172C1B",
    x"3216F119",
    x"3216B62F",
    x"32167B5B",
    x"3216409E",
    x"321605F8",
    x"3215CB6A",
    x"321590F1",
    x"32155690",
    x"32151C46",
    x"3214E212",
    x"3214A7F5",
    x"32146DEF",
    x"321433FF",
    x"3213FA26",
    x"3213C064",
    x"321386B8",
    x"32134D23",
    x"321313A4",
    x"3212DA3B",
    x"3212A0E9",
    x"321267AE",
    x"32122E88",
    x"3211F579",
    x"3211BC80",
    x"3211839E",
    x"32114AD2",
    x"3211121B",
    x"3210D97B",
    x"3210A0F2",
    x"3210687E",
    x"32103020",
    x"320FF7D8",
    x"320FBFA6",
    x"320F878A",
    x"320F4F84",
    x"320F1794",
    x"320EDFBA",
    x"320EA7F5",
    x"320E7047",
    x"320E38AE",
    x"320E012A",
    x"320DC9BD",
    x"320D9265",
    x"320D5B22",
    x"320D23F6",
    x"320CECDE",
    x"320CB5DC",
    x"320C7EF0",
    x"320C4819",
    x"320C1158",
    x"320BDAAC",
    x"320BA415",
    x"320B6D94",
    x"320B3727",
    x"320B00D0",
    x"320ACA8F",
    x"320A9462",
    x"320A5E4B",
    x"320A2849",
    x"3209F25B",
    x"3209BC83",
    x"320986C0",
    x"32095112",
    x"32091B79",
    x"3208E5F4",
    x"3208B085",
    x"32087B2A",
    x"320845E5",
    x"320810B4",
    x"3207DB98",
    x"3207A690",
    x"3207719E",
    x"32073CC0",
    x"320707F6",
    x"3206D341",
    x"32069EA1",
    x"32066A15",
    x"3206359E",
    x"3206013B",
    x"3205CCED",
    x"320598B3",
    x"3205648E",
    x"3205307D",
    x"3204FC80",
    x"3204C898",
    x"320494C3",
    x"32046103",
    x"32042D57",
    x"3203F9C0",
    x"3203C63C",
    x"320392CD",
    x"32035F72",
    x"32032C2A",
    x"3202F8F7",
    x"3202C5D8",
    x"320292CD",
    x"32025FD5",
    x"32022CF2",
    x"3201FA22",
    x"3201C766",
    x"320194BE",
    x"3201622A",
    x"32012FAA",
    x"3200FD3D",
    x"3200CAE4",
    x"3200989E",
    x"3200666C",
    x"3200344E",
    x"32000244",
    x"31FFA099",
    x"31FF3CD2",
    x"31FED931",
    x"31FE75B8",
    x"31FE1265",
    x"31FDAF3A",
    x"31FD4C34",
    x"31FCE956",
    x"31FC869E",
    x"31FC240D",
    x"31FBC1A2",
    x"31FB5F5E",
    x"31FAFD3F",
    x"31FA9B48",
    x"31FA3976",
    x"31F9D7CB",
    x"31F97646",
    x"31F914E6",
    x"31F8B3AD",
    x"31F8529A",
    x"31F7F1AD",
    x"31F790E5",
    x"31F73043",
    x"31F6CFC7",
    x"31F66F71",
    x"31F60F40",
    x"31F5AF35",
    x"31F54F4F",
    x"31F4EF8F",
    x"31F48FF4",
    x"31F4307F",
    x"31F3D12E",
    x"31F37203",
    x"31F312FD",
    x"31F2B41C",
    x"31F25561",
    x"31F1F6CA",
    x"31F19858",
    x"31F13A0B",
    x"31F0DBE2",
    x"31F07DDF",
    x"31F02000",
    x"31EFC246",
    x"31EF64B0",
    x"31EF073F",
    x"31EEA9F3",
    x"31EE4CCA",
    x"31EDEFC7",
    x"31ED92E7",
    x"31ED362C",
    x"31ECD995",
    x"31EC7D22",
    x"31EC20D3",
    x"31EBC4A8",
    x"31EB68A1",
    x"31EB0CBE",
    x"31EAB0FF",
    x"31EA5564",
    x"31E9F9ED",
    x"31E99E99",
    x"31E94369",
    x"31E8E85C",
    x"31E88D73",
    x"31E832AE",
    x"31E7D80B",
    x"31E77D8D",
    x"31E72331",
    x"31E6C8F9",
    x"31E66EE4",
    x"31E614F3",
    x"31E5BB24",
    x"31E56178",
    x"31E507F0",
    x"31E4AE8A",
    x"31E45547",
    x"31E3FC27",
    x"31E3A32A",
    x"31E34A50",
    x"31E2F198",
    x"31E29903",
    x"31E24091",
    x"31E1E841",
    x"31E19013",
    x"31E13808",
    x"31E0E01F",
    x"31E08859",
    x"31E030B5",
    x"31DFD933",
    x"31DF81D3",
    x"31DF2A96",
    x"31DED37A",
    x"31DE7C80",
    x"31DE25A9",
    x"31DDCEF3",
    x"31DD785F",
    x"31DD21ED",
    x"31DCCB9C",
    x"31DC756E",
    x"31DC1F61",
    x"31DBC975",
    x"31DB73AB",
    x"31DB1E03",
    x"31DAC87C",
    x"31DA7316",
    x"31DA1DD2",
    x"31D9C8AF",
    x"31D973AD",
    x"31D91ECC",
    x"31D8CA0D",
    x"31D8756F",
    x"31D820F1",
    x"31D7CC95",
    x"31D77859",
    x"31D7243F",
    x"31D6D045",
    x"31D67C6C",
    x"31D628B4",
    x"31D5D51C",
    x"31D581A5",
    x"31D52E4F",
    x"31D4DB19",
    x"31D48804",
    x"31D4350F",
    x"31D3E23A",
    x"31D38F86",
    x"31D33CF2",
    x"31D2EA7E",
    x"31D2982B",
    x"31D245F8",
    x"31D1F3E4",
    x"31D1A1F1",
    x"31D1501E",
    x"31D0FE6A",
    x"31D0ACD7",
    x"31D05B63",
    x"31D00A10",
    x"31CFB8DB",
    x"31CF67C7",
    x"31CF16D2",
    x"31CEC5FD",
    x"31CE7548",
    x"31CE24B2",
    x"31CDD43B",
    x"31CD83E4",
    x"31CD33AC",
    x"31CCE393",
    x"31CC939A",
    x"31CC43C0",
    x"31CBF405",
    x"31CBA469",
    x"31CB54ED",
    x"31CB058F",
    x"31CAB650",
    x"31CA6731",
    x"31CA1830",
    x"31C9C94E",
    x"31C97A8A",
    x"31C92BE6",
    x"31C8DD60",
    x"31C88EF9",
    x"31C840B0",
    x"31C7F286",
    x"31C7A47B",
    x"31C7568E",
    x"31C708BF",
    x"31C6BB0F",
    x"31C66D7D",
    x"31C6200A",
    x"31C5D2B4",
    x"31C5857D",
    x"31C53864",
    x"31C4EB69",
    x"31C49E8C",
    x"31C451CD",
    x"31C4052C",
    x"31C3B8A9",
    x"31C36C44",
    x"31C31FFC",
    x"31C2D3D3",
    x"31C287C7",
    x"31C23BD9",
    x"31C1F008",
    x"31C1A455",
    x"31C158C0",
    x"31C10D48",
    x"31C0C1ED",
    x"31C076B0",
    x"31C02B90",
    x"31BFE08E",
    x"31BF95A9",
    x"31BF4AE1",
    x"31BF0037",
    x"31BEB5A9",
    x"31BE6B39",
    x"31BE20E5",
    x"31BDD6AF",
    x"31BD8C95",
    x"31BD4299",
    x"31BCF8B9",
    x"31BCAEF7",
    x"31BC6551",
    x"31BC1BC8",
    x"31BBD25B",
    x"31BB890B",
    x"31BB3FD8",
    x"31BAF6C1",
    x"31BAADC7",
    x"31BA64EA",
    x"31BA1C28",
    x"31B9D383",
    x"31B98AFB",
    x"31B9428F",
    x"31B8FA3F",
    x"31B8B20B",
    x"31B869F4",
    x"31B821F9",
    x"31B7DA19",
    x"31B79256",
    x"31B74AAF",
    x"31B70324",
    x"31B6BBB5",
    x"31B67461",
    x"31B62D2A",
    x"31B5E60E",
    x"31B59F0E",
    x"31B5582A",
    x"31B51161",
    x"31B4CAB4",
    x"31B48423",
    x"31B43DAD",
    x"31B3F752",
    x"31B3B114",
    x"31B36AF0",
    x"31B324E8",
    x"31B2DEFB",
    x"31B2992A",
    x"31B25374",
    x"31B20DD9",
    x"31B1C859",
    x"31B182F4",
    x"31B13DAA",
    x"31B0F87C",
    x"31B0B368",
    x"31B06E70",
    x"31B02992",
    x"31AFE4CF",
    x"31AFA027",
    x"31AF5B9A",
    x"31AF1728",
    x"31AED2D0",
    x"31AE8E93",
    x"31AE4A71",
    x"31AE0669",
    x"31ADC27B",
    x"31AD7EA9",
    x"31AD3AF1",
    x"31ACF753",
    x"31ACB3CF",
    x"31AC7066",
    x"31AC2D17",
    x"31ABE9E3",
    x"31ABA6C9",
    x"31AB63C9",
    x"31AB20E3",
    x"31AADE17",
    x"31AA9B65",
    x"31AA58CE",
    x"31AA1650",
    x"31A9D3EC",
    x"31A991A2",
    x"31A94F72",
    x"31A90D5C",
    x"31A8CB60",
    x"31A8897D",
    x"31A847B4",
    x"31A80605",
    x"31A7C470",
    x"31A782F4",
    x"31A74191",
    x"31A70049",
    x"31A6BF19",
    x"31A67E03",
    x"31A63D07",
    x"31A5FC24",
    x"31A5BB5A",
    x"31A57AA9",
    x"31A53A12",
    x"31A4F994",
    x"31A4B92F",
    x"31A478E3",
    x"31A438B0",
    x"31A3F897",
    x"31A3B896",
    x"31A378AF",
    x"31A338E0",
    x"31A2F92A",
    x"31A2B98D",
    x"31A27A09",
    x"31A23A9E",
    x"31A1FB4B",
    x"31A1BC12",
    x"31A17CF0",
    x"31A13DE8",
    x"31A0FEF8",
    x"31A0C021",
    x"31A08162",
    x"31A042BC",
    x"31A0042E",
    x"319FC5B8",
    x"319F875B",
    x"319F4917",
    x"319F0AEA",
    x"319ECCD6",
    x"319E8EDA",
    x"319E50F6",
    x"319E132B",
    x"319DD577",
    x"319D97DC",
    x"319D5A59",
    x"319D1CED",
    x"319CDF9A",
    x"319CA25F",
    x"319C653B",
    x"319C2830",
    x"319BEB3C",
    x"319BAE60",
    x"319B719C",
    x"319B34EF",
    x"319AF85A",
    x"319ABBDD",
    x"319A7F78",
    x"319A432A",
    x"319A06F3",
    x"3199CAD4",
    x"31998ECD",
    x"319952DC",
    x"31991704",
    x"3198DB42",
    x"31989F99",
    x"31986406",
    x"3198288A",
    x"3197ED26",
    x"3197B1D9",
    x"319776A3",
    x"31973B84",
    x"3197007D",
    x"3196C58C",
    x"31968AB2",
    x"31964FF0",
    x"31961544",
    x"3195DAAF",
    x"3195A031",
    x"319565CA",
    x"31952B79",
    x"3194F140",
    x"3194B71D",
    x"31947D11",
    x"3194431B",
    x"3194093C",
    x"3193CF74",
    x"319395C2",
    x"31935C27",
    x"319322A2",
    x"3192E934",
    x"3192AFDC",
    x"3192769B",
    x"31923D6F",
    x"3192045B",
    x"3191CB5C",
    x"31919274",
    x"319159A2",
    x"319120E6",
    x"3190E840",
    x"3190AFB0",
    x"31907737",
    x"31903ED3",
    x"31900685",
    x"318FCE4E",
    x"318F962C",
    x"318F5E21",
    x"318F262B",
    x"318EEE4B",
    x"318EB681",
    x"318E7ECC",
    x"318E472D",
    x"318E0FA5",
    x"318DD831",
    x"318DA0D4",
    x"318D698C",
    x"318D3259",
    x"318CFB3C",
    x"318CC435",
    x"318C8D43",
    x"318C5666",
    x"318C1F9F",
    x"318BE8EE",
    x"318BB251",
    x"318B7BCA",
    x"318B4559",
    x"318B0EFC",
    x"318AD8B5",
    x"318AA283",
    x"318A6C66",
    x"318A365E",
    x"318A006C",
    x"3189CA8E",
    x"318994C5",
    x"31895F12",
    x"31892973",
    x"3188F3E9",
    x"3188BE74",
    x"31888914",
    x"318853C9",
    x"31881E93",
    x"3187E971",
    x"3187B465",
    x"31877F6D",
    x"31874A89",
    x"318715BA",
    x"3186E100",
    x"3186AC5A",
    x"318677C9",
    x"3186434D",
    x"31860EE5",
    x"3185DA91",
    x"3185A652",
    x"31857227",
    x"31853E11",
    x"31850A0F",
    x"3184D621",
    x"3184A247",
    x"31846E82",
    x"31843AD1",
    x"31840734",
    x"3183D3AC",
    x"3183A037",
    x"31836CD6",
    x"3183398A",
    x"31830651",
    x"3182D32D",
    x"3182A01C",
    x"31826D20",
    x"31823A37",
    x"31820762",
    x"3181D4A1",
    x"3181A1F4",
    x"31816F5B",
    x"31813CD5",
    x"31810A63",
    x"3180D805",
    x"3180A5BA",
    x"31807384",
    x"31804160",
    x"31800F50",
    x"317FBAA9",
    x"317F56D7",
    x"317EF32D",
    x"317E8FA9",
    x"317E2C4C",
    x"317DC916",
    x"317D6607",
    x"317D031F",
    x"317CA05D",
    x"317C3DC1",
    x"317BDB4D",
    x"317B78FE",
    x"317B16D6",
    x"317AB4D4",
    x"317A52F9",
    x"3179F143",
    x"31798FB4",
    x"31792E4B",
    x"3178CD08",
    x"31786BEB",
    x"31780AF4",
    x"3177AA22",
    x"31774977",
    x"3176E8F1",
    x"31768891",
    x"31762856",
    x"3175C841",
    x"31756852",
    x"31750888",
    x"3174A8E3",
    x"31744964",
    x"3173EA0A",
    x"31738AD5",
    x"31732BC5",
    x"3172CCDB",
    x"31726E15",
    x"31720F75",
    x"3171B0F9",
    x"317152A2",
    x"3170F470",
    x"31709663",
    x"3170387B",
    x"316FDAB7",
    x"316F7D18",
    x"316F1F9D",
    x"316EC247",
    x"316E6516",
    x"316E0808",
    x"316DAB1F",
    x"316D4E5B",
    x"316CF1BA",
    x"316C953E",
    x"316C38E6",
    x"316BDCB1",
    x"316B80A1",
    x"316B24B5",
    x"316AC8EC",
    x"316A6D48",
    x"316A11C7",
    x"3169B66A",
    x"31695B30",
    x"3169001B",
    x"3168A528",
    x"31684A5A",
    x"3167EFAE",
    x"31679526",
    x"31673AC2",
    x"3166E080",
    x"31668662",
    x"31662C67",
    x"3165D290",
    x"316578DB",
    x"31651F49",
    x"3164C5DA",
    x"31646C8F",
    x"31641366",
    x"3163BA5F",
    x"3163617C",
    x"316308BB",
    x"3162B01D",
    x"316257A2",
    x"3161FF49",
    x"3161A712",
    x"31614EFE",
    x"3160F70C",
    x"31609F3D",
    x"31604790",
    x"315FF005",
    x"315F989C",
    x"315F4156",
    x"315EEA31",
    x"315E932F",
    x"315E3C4E",
    x"315DE590",
    x"315D8EF3",
    x"315D3878",
    x"315CE21F",
    x"315C8BE7",
    x"315C35D2",
    x"315BDFDD",
    x"315B8A0B",
    x"315B345A",
    x"315ADECA",
    x"315A895B",
    x"315A340E",
    x"3159DEE3",
    x"315989D8",
    x"315934EF",
    x"3158E027",
    x"31588B80",
    x"315836FA",
    x"3157E295",
    x"31578E51",
    x"31573A2E",
    x"3156E62B",
    x"3156924A",
    x"31563E89",
    x"3155EAE9",
    x"3155976A",
    x"3155440B",
    x"3154F0CC",
    x"31549DAF",
    x"31544AB1",
    x"3153F7D4",
    x"3153A518",
    x"3153527B",
    x"3152FFFF",
    x"3152ADA3",
    x"31525B67",
    x"3152094C",
    x"3151B750",
    x"31516575",
    x"315113B9",
    x"3150C21D",
    x"315070A1",
    x"31501F45",
    x"314FCE09",
    x"314F7CEC",
    x"314F2BEF",
    x"314EDB12",
    x"314E8A54",
    x"314E39B6",
    x"314DE937",
    x"314D98D8",
    x"314D4897",
    x"314CF877",
    x"314CA875",
    x"314C5893",
    x"314C08D0",
    x"314BB92C",
    x"314B69A7",
    x"314B1A42",
    x"314ACAFB",
    x"314A7BD3",
    x"314A2CCA",
    x"3149DDE0",
    x"31498F15",
    x"31494068",
    x"3148F1DA",
    x"3148A36B",
    x"3148551B",
    x"314806E9",
    x"3147B8D5",
    x"31476AE0",
    x"31471D0A",
    x"3146CF52",
    x"314681B8",
    x"3146343C",
    x"3145E6DF",
    x"314599A0",
    x"31454C7F",
    x"3144FF7C",
    x"3144B297",
    x"314465D1",
    x"31441928",
    x"3143CC9D",
    x"31438030",
    x"314333E1",
    x"3142E7AF",
    x"31429B9C",
    x"31424FA6",
    x"314203CE",
    x"3141B813",
    x"31416C76",
    x"314120F6",
    x"3140D594",
    x"31408A4F",
    x"31403F28",
    x"313FF41E",
    x"313FA931",
    x"313F5E62",
    x"313F13AF",
    x"313EC91A",
    x"313E7EA2",
    x"313E3447",
    x"313DEA09",
    x"313D9FE9",
    x"313D55E5",
    x"313D0BFD",
    x"313CC233",
    x"313C7886",
    x"313C2EF5",
    x"313BE581",
    x"313B9C2A",
    x"313B52EF",
    x"313B09D1",
    x"313AC0CF",
    x"313A77EA",
    x"313A2F22",
    x"3139E675",
    x"31399DE5",
    x"31395572",
    x"31390D1B",
    x"3138C4E0",
    x"31387CC1",
    x"313834BE",
    x"3137ECD8",
    x"3137A50D",
    x"31375D5F",
    x"313715CC",
    x"3136CE56",
    x"313686FB",
    x"31363FBC",
    x"3135F899",
    x"3135B192",
    x"31356AA6",
    x"313523D7",
    x"3134DD22",
    x"3134968A",
    x"3134500D",
    x"313409AB",
    x"3133C365",
    x"31337D3B",
    x"3133372B",
    x"3132F138",
    x"3132AB5F",
    x"313265A2",
    x"31322000",
    x"3131DA79",
    x"3131950D",
    x"31314FBC",
    x"31310A87",
    x"3130C56C",
    x"3130806C",
    x"31303B88",
    x"312FF6BE",
    x"312FB20F",
    x"312F6D7B",
    x"312F2901",
    x"312EE4A3",
    x"312EA05F",
    x"312E5C35",
    x"312E1827",
    x"312DD432",
    x"312D9059",
    x"312D4C9A",
    x"312D08F5",
    x"312CC56B",
    x"312C81FB",
    x"312C3EA5",
    x"312BFB6A",
    x"312BB849",
    x"312B7542",
    x"312B3255",
    x"312AEF82",
    x"312AACCA",
    x"312A6A2B",
    x"312A27A7",
    x"3129E53C",
    x"3129A2EC",
    x"312960B5",
    x"31291E98",
    x"3128DC95",
    x"31289AAC",
    x"312858DC",
    x"31281726",
    x"3127D58A",
    x"31279408",
    x"3127529F",
    x"3127114F",
    x"3126D019",
    x"31268EFC",
    x"31264DF9",
    x"31260D10",
    x"3125CC3F",
    x"31258B88",
    x"31254AEA",
    x"31250A65",
    x"3124C9FA",
    x"312489A8",
    x"3124496E",
    x"3124094E",
    x"3123C947",
    x"31238959",
    x"31234984",
    x"312309C8",
    x"3122CA24",
    x"31228A9A",
    x"31224B28",
    x"31220BCF",
    x"3121CC8F",
    x"31218D67",
    x"31214E58",
    x"31210F62",
    x"3120D084",
    x"312091BF",
    x"31205312",
    x"3120147E",
    x"311FD602",
    x"311F979F",
    x"311F5954",
    x"311F1B21",
    x"311EDD07",
    x"311E9F04",
    x"311E611A",
    x"311E2348",
    x"311DE58F",
    x"311DA7ED",
    x"311D6A64",
    x"311D2CF2",
    x"311CEF98",
    x"311CB257",
    x"311C752D",
    x"311C381B",
    x"311BFB21",
    x"311BBE3F",
    x"311B8175",
    x"311B44C2",
    x"311B0827",
    x"311ACBA3",
    x"311A8F38",
    x"311A52E4",
    x"311A16A7",
    x"3119DA82",
    x"31199E74",
    x"3119627E",
    x"3119269F",
    x"3118EAD8",
    x"3118AF28",
    x"3118738F",
    x"3118380E",
    x"3117FCA3",
    x"3117C150",
    x"31178614",
    x"31174AEF",
    x"31170FE2",
    x"3116D4EB",
    x"31169A0B",
    x"31165F43",
    x"31162491",
    x"3115E9F6",
    x"3115AF72",
    x"31157505",
    x"31153AAF",
    x"3115006F",
    x"3114C646",
    x"31148C34",
    x"31145239",
    x"31141854",
    x"3113DE86",
    x"3113A4CE",
    x"31136B2D",
    x"311331A2",
    x"3112F82E",
    x"3112BED0",
    x"31128589",
    x"31124C58",
    x"3112133D",
    x"3111DA39",
    x"3111A14B",
    x"31116873",
    x"31112FB1",
    x"3110F706",
    x"3110BE70",
    x"311085F1",
    x"31104D88",
    x"31101534",
    x"310FDCF7",
    x"310FA4D0",
    x"310F6CBE",
    x"310F34C3",
    x"310EFCDD",
    x"310EC50D",
    x"310E8D53",
    x"310E55AF",
    x"310E1E20",
    x"310DE6A7",
    x"310DAF44",
    x"310D77F6",
    x"310D40BE",
    x"310D099C",
    x"310CD28F",
    x"310C9B97",
    x"310C64B5",
    x"310C2DE8",
    x"310BF731",
    x"310BC08F",
    x"310B8A03",
    x"310B538C",
    x"310B1D2A",
    x"310AE6DD",
    x"310AB0A5",
    x"310A7A83",
    x"310A4475",
    x"310A0E7D",
    x"3109D89A",
    x"3109A2CC",
    x"31096D13",
    x"3109376F",
    x"310901E0",
    x"3108CC65",
    x"31089700",
    x"310861AF",
    x"31082C74",
    x"3107F74D",
    x"3107C23A",
    x"31078D3D",
    x"31075854",
    x"31072380",
    x"3106EEC0",
    x"3106BA15",
    x"3106857F",
    x"310650FD",
    x"31061C90",
    x"3105E837",
    x"3105B3F2",
    x"31057FC2",
    x"31054BA6",
    x"3105179F",
    x"3104E3AC",
    x"3104AFCD",
    x"31047C03",
    x"3104484C",
    x"310414AA",
    x"3103E11C",
    x"3103ADA2",
    x"31037A3C",
    x"310346EB",
    x"310313AD",
    x"3102E083",
    x"3102AD6E",
    x"31027A6C",
    x"3102477E",
    x"310214A4",
    x"3101E1DE",
    x"3101AF2B",
    x"31017C8D",
    x"31014A02",
    x"3101178B",
    x"3100E528",
    x"3100B2D8",
    x"3100809C",
    x"31004E74",
    x"31001C5F",
    x"30FFD4BB",
    x"30FF70DF",
    x"30FF0D2B",
    x"30FEA99D",
    x"30FE4636",
    x"30FDE2F6",
    x"30FD7FDD",
    x"30FD1CEA",
    x"30FCBA1E",
    x"30FC5779",
    x"30FBF4FA",
    x"30FB92A1",
    x"30FB306F",
    x"30FACE63",
    x"30FA6C7E",
    x"30FA0ABF",
    x"30F9A925",
    x"30F947B2",
    x"30F8E665",
    x"30F8853E",
    x"30F8243D",
    x"30F7C362",
    x"30F762AD",
    x"30F7021D",
    x"30F6A1B3",
    x"30F6416F",
    x"30F5E150",
    x"30F58157",
    x"30F52183",
    x"30F4C1D4",
    x"30F4624B",
    x"30F402E8",
    x"30F3A3A9",
    x"30F34490",
    x"30F2E59B",
    x"30F286CC",
    x"30F22822",
    x"30F1C99D",
    x"30F16B3D",
    x"30F10D01",
    x"30F0AEEA",
    x"30F050F8",
    x"30EFF32B",
    x"30EF9582",
    x"30EF37FE",
    x"30EEDA9F",
    x"30EE7D64",
    x"30EE204D",
    x"30EDC35A",
    x"30ED668C",
    x"30ED09E2",
    x"30ECAD5C",
    x"30EC50FB",
    x"30EBF4BD",
    x"30EB98A3",
    x"30EB3CAE",
    x"30EAE0DC",
    x"30EA852E",
    x"30EA29A4",
    x"30E9CE3E",
    x"30E972FB",
    x"30E917DC",
    x"30E8BCE0",
    x"30E86208",
    x"30E80754",
    x"30E7ACC2",
    x"30E75255",
    x"30E6F80A",
    x"30E69DE3",
    x"30E643DF",
    x"30E5E9FE",
    x"30E59040",
    x"30E536A5",
    x"30E4DD2D",
    x"30E483D8",
    x"30E42AA6",
    x"30E3D197",
    x"30E378AA",
    x"30E31FE1",
    x"30E2C739",
    x"30E26EB5",
    x"30E21653",
    x"30E1BE13",
    x"30E165F6",
    x"30E10DFC",
    x"30E0B623",
    x"30E05E6D",
    x"30E006DA",
    x"30DFAF68",
    x"30DF5819",
    x"30DF00EB",
    x"30DEA9E0",
    x"30DE52F7",
    x"30DDFC2F",
    x"30DDA589",
    x"30DD4F06",
    x"30DCF8A4",
    x"30DCA263",
    x"30DC4C45",
    x"30DBF648",
    x"30DBA06C",
    x"30DB4AB3",
    x"30DAF51A",
    x"30DA9FA3",
    x"30DA4A4D",
    x"30D9F519",
    x"30D9A006",
    x"30D94B14",
    x"30D8F643",
    x"30D8A193",
    x"30D84D05",
    x"30D7F897",
    x"30D7A44B",
    x"30D7501F",
    x"30D6FC14",
    x"30D6A82A",
    x"30D65461",
    x"30D600B8",
    x"30D5AD30",
    x"30D559C9",
    x"30D50682",
    x"30D4B35C",
    x"30D46056",
    x"30D40D70",
    x"30D3BAAB",
    x"30D36806",
    x"30D31582",
    x"30D2C31E",
    x"30D270DA",
    x"30D21EB5",
    x"30D1CCB2",
    x"30D17ACE",
    x"30D1290A",
    x"30D0D765",
    x"30D085E1",
    x"30D0347D",
    x"30CFE338",
    x"30CF9213",
    x"30CF410E",
    x"30CEF029",
    x"30CE9F62",
    x"30CE4EBC",
    x"30CDFE35",
    x"30CDADCD",
    x"30CD5D85",
    x"30CD0D5C",
    x"30CCBD53",
    x"30CC6D68",
    x"30CC1D9D",
    x"30CBCDF1",
    x"30CB7E64",
    x"30CB2EF6",
    x"30CADFA8",
    x"30CA9078",
    x"30CA4167",
    x"30C9F275",
    x"30C9A3A1",
    x"30C954ED",
    x"30C90657",
    x"30C8B7E0",
    x"30C86987",
    x"30C81B4D",
    x"30C7CD32",
    x"30C77F35",
    x"30C73157",
    x"30C6E396",
    x"30C695F5",
    x"30C64871",
    x"30C5FB0C",
    x"30C5ADC5",
    x"30C5609C",
    x"30C51392",
    x"30C4C6A5",
    x"30C479D6",
    x"30C42D26",
    x"30C3E093",
    x"30C3941E",
    x"30C347C7",
    x"30C2FB8E",
    x"30C2AF73",
    x"30C26375",
    x"30C21795",
    x"30C1CBD3",
    x"30C1802E",
    x"30C134A7",
    x"30C0E93D",
    x"30C09DF0",
    x"30C052C1",
    x"30C007B0",
    x"30BFBCBB",
    x"30BF71E4",
    x"30BF272A",
    x"30BEDC8E",
    x"30BE920E",
    x"30BE47AB",
    x"30BDFD66",
    x"30BDB33D",
    x"30BD6932",
    x"30BD1F43",
    x"30BCD571",
    x"30BC8BBD",
    x"30BC4224",
    x"30BBF8A9",
    x"30BBAF4A",
    x"30BB6608",
    x"30BB1CE2",
    x"30BAD3D9",
    x"30BA8AED",
    x"30BA421D",
    x"30B9F969",
    x"30B9B0D2",
    x"30B96857",
    x"30B91FF8",
    x"30B8D7B6",
    x"30B88F90",
    x"30B84786",
    x"30B7FF98",
    x"30B7B7C6",
    x"30B77010",
    x"30B72877",
    x"30B6E0F9",
    x"30B69997",
    x"30B65251",
    x"30B60B26",
    x"30B5C418",
    x"30B57D25",
    x"30B5364E",
    x"30B4EF93",
    x"30B4A8F3",
    x"30B4626F",
    x"30B41C06",
    x"30B3D5B9",
    x"30B38F87",
    x"30B34971",
    x"30B30376",
    x"30B2BD96",
    x"30B277D2",
    x"30B23228",
    x"30B1EC9A",
    x"30B1A728",
    x"30B161D0",
    x"30B11C93",
    x"30B0D771",
    x"30B0926B",
    x"30B04D7F",
    x"30B008AE",
    x"30AFC3F8",
    x"30AF7F5D",
    x"30AF3ADD",
    x"30AEF677",
    x"30AEB22C",
    x"30AE6DFC",
    x"30AE29E6",
    x"30ADE5EB",
    x"30ADA20B",
    x"30AD5E45",
    x"30AD1A99",
    x"30ACD708",
    x"30AC9391",
    x"30AC5034",
    x"30AC0CF2",
    x"30ABC9CA",
    x"30AB86BD",
    x"30AB43C9",
    x"30AB00F0",
    x"30AABE30",
    x"30AA7B8B",
    x"30AA3900",
    x"30A9F68E",
    x"30A9B437",
    x"30A971FA",
    x"30A92FD6",
    x"30A8EDCC",
    x"30A8ABDC",
    x"30A86A06",
    x"30A82849",
    x"30A7E6A7",
    x"30A7A51D",
    x"30A763AE",
    x"30A72257",
    x"30A6E11B",
    x"30A69FF7",
    x"30A65EEE",
    x"30A61DFD",
    x"30A5DD26",
    x"30A59C69",
    x"30A55BC4",
    x"30A51B39",
    x"30A4DAC7",
    x"30A49A6E",
    x"30A45A2E",
    x"30A41A07",
    x"30A3D9FA",
    x"30A39A05",
    x"30A35A29",
    x"30A31A67",
    x"30A2DABD",
    x"30A29B2C",
    x"30A25BB4",
    x"30A21C54",
    x"30A1DD0D",
    x"30A19DDF",
    x"30A15ECA",
    x"30A11FCD",
    x"30A0E0E9",
    x"30A0A21E",
    x"30A0636B",
    x"30A024D0",
    x"309FE64E",
    x"309FA7E4",
    x"309F6993",
    x"309F2B59",
    x"309EED39",
    x"309EAF30",
    x"309E7140",
    x"309E3368",
    x"309DF5A8",
    x"309DB800",
    x"309D7A70",
    x"309D3CF8",
    x"309CFF98",
    x"309CC250",
    x"309C8520",
    x"309C4808",
    x"309C0B08",
    x"309BCE20",
    x"309B914F",
    x"309B5496",
    x"309B17F5",
    x"309ADB6B",
    x"309A9EFA",
    x"309A629F",
    x"309A265C",
    x"3099EA31",
    x"3099AE1E",
    x"30997221",
    x"3099363C",
    x"3098FA6F",
    x"3098BEB9",
    x"3098831A",
    x"30984792",
    x"30980C22",
    x"3097D0C9",
    x"30979587",
    x"30975A5C",
    x"30971F48",
    x"3096E44B",
    x"3096A966",
    x"30966E97",
    x"309633DF",
    x"3095F93F",
    x"3095BEB5",
    x"30958442",
    x"309549E5",
    x"30950FA0",
    x"3094D571",
    x"30949B59",
    x"30946158",
    x"3094276D",
    x"3093ED99",
    x"3093B3DB",
    x"30937A34",
    x"309340A4",
    x"3093072A",
    x"3092CDC6",
    x"30929479",
    x"30925B42",
    x"30922222",
    x"3091E918",
    x"3091B024",
    x"30917746",
    x"30913E7E",
    x"309105CD",
    x"3090CD32",
    x"309094AD",
    x"30905C3E",
    x"309023E5",
    x"308FEBA2",
    x"308FB375",
    x"308F7B5E",
    x"308F435C",
    x"308F0B71",
    x"308ED39B",
    x"308E9BDC",
    x"308E6432",
    x"308E2C9D",
    x"308DF51F",
    x"308DBDB6",
    x"308D8662",
    x"308D4F25",
    x"308D17FD",
    x"308CE0EA",
    x"308CA9ED",
    x"308C7305",
    x"308C3C33",
    x"308C0576",
    x"308BCECF",
    x"308B983D",
    x"308B61C0",
    x"308B2B58",
    x"308AF506",
    x"308ABEC9",
    x"308A88A1",
    x"308A528E",
    x"308A1C90",
    x"3089E6A8",
    x"3089B0D4",
    x"30897B16",
    x"3089456C",
    x"30890FD7",
    x"3088DA58",
    x"3088A4ED",
    x"30886F97",
    x"30883A56",
    x"30880529",
    x"3087D011",
    x"30879B0F",
    x"30876620",
    x"30873147",
    x"3086FC82",
    x"3086C7D1",
    x"30869336",
    x"30865EAE",
    x"30862A3C",
    x"3085F5DD",
    x"3085C194",
    x"30858D5E",
    x"3085593D",
    x"30852531",
    x"3084F138",
    x"3084BD54",
    x"30848984",
    x"308455C9",
    x"30842221",
    x"3083EE8E",
    x"3083BB0F",
    x"308387A4",
    x"3083544D",
    x"3083210A",
    x"3082EDDB",
    x"3082BAC0",
    x"308287B9",
    x"308254C6",
    x"308221E7",
    x"3081EF1C",
    x"3081BC64",
    x"308189C0",
    x"30815730",
    x"308124B4",
    x"3080F24C",
    x"3080BFF7",
    x"30808DB6",
    x"30805B88",
    x"3080296E",
    x"307FEED0",
    x"307F8AEA",
    x"307F272B",
    x"307EC393",
    x"307E6022",
    x"307DFCD8",
    x"307D99B5",
    x"307D36B8",
    x"307CD3E2",
    x"307C7132",
    x"307C0EA9",
    x"307BAC47",
    x"307B4A0B",
    x"307AE7F5",
    x"307A8606",
    x"307A243C",
    x"3079C299",
    x"3079611C",
    x"3078FFC5",
    x"30789E94",
    x"30783D8A",
    x"3077DCA4",
    x"30777BE5",
    x"30771B4C",
    x"3076BAD8",
    x"30765A8A",
    x"3075FA61",
    x"30759A5E",
    x"30753A80",
    x"3074DAC8",
    x"30747B35",
    x"30741BC8",
    x"3073BC80",
    x"30735D5D",
    x"3072FE5F",
    x"30729F86",
    x"307240D2",
    x"3071E243",
    x"307183D9",
    x"30712594",
    x"3070C774",
    x"30706978",
    x"30700BA2",
    x"306FADEF",
    x"306F5062",
    x"306EF2F8",
    x"306E95B4",
    x"306E3894",
    x"306DDB98",
    x"306D7EC0",
    x"306D220D",
    x"306CC57D",
    x"306C6912",
    x"306C0CCB",
    x"306BB0A8",
    x"306B54A9",
    x"306AF8CE",
    x"306A9D17",
    x"306A4183",
    x"3069E614",
    x"30698AC8",
    x"30692F9F",
    x"3068D49A",
    x"306879B9",
    x"30681EFB",
    x"3067C461",
    x"306769EA",
    x"30670F96",
    x"3066B566",
    x"30665B58",
    x"3066016E",
    x"3065A7A7",
    x"30654E03",
    x"3064F482",
    x"30649B24",
    x"306441E9",
    x"3063E8D1",
    x"30638FDB",
    x"30633708",
    x"3062DE58",
    x"306285CB",
    x"30622D60",
    x"3061D517",
    x"30617CF1",
    x"306124ED",
    x"3060CD0C",
    x"3060754D",
    x"30601DB1",
    x"305FC636",
    x"305F6EDE",
    x"305F17A7",
    x"305EC093",
    x"305E69A1",
    x"305E12D1",
    x"305DBC22",
    x"305D6596",
    x"305D0F2B",
    x"305CB8E2",
    x"305C62BA",
    x"305C0CB5",
    x"305BB6D0",
    x"305B610E",
    x"305B0B6D",
    x"305AB5ED",
    x"305A608E",
    x"305A0B51",
    x"3059B636",
    x"3059613B",
    x"30590C62",
    x"3058B7A9",
    x"30586312",
    x"30580E9C",
    x"3057BA47",
    x"30576612",
    x"305711FF",
    x"3056BE0C",
    x"30566A3A",
    x"30561689",
    x"3055C2F9",
    x"30556F89",
    x"30551C3A",
    x"3054C90B",
    x"305475FD",
    x"3054230F",
    x"3053D041",
    x"30537D94",
    x"30532B07",
    x"3052D89A",
    x"3052864E",
    x"30523421",
    x"3051E215",
    x"30519029",
    x"30513E5C",
    x"3050ECB0",
    x"30509B23",
    x"305049B7",
    x"304FF86A",
    x"304FA73D",
    x"304F562F",
    x"304F0541",
    x"304EB473",
    x"304E63C4",
    x"304E1335",
    x"304DC2C5",
    x"304D7275",
    x"304D2244",
    x"304CD232",
    x"304C8240",
    x"304C326C",
    x"304BE2B8",
    x"304B9323",
    x"304B43AD",
    x"304AF456",
    x"304AA51E",
    x"304A5605",
    x"304A070B",
    x"3049B830",
    x"30496973",
    x"30491AD5",
    x"3048CC56",
    x"30487DF6",
    x"30482FB4",
    x"3047E190",
    x"3047938C",
    x"304745A5",
    x"3046F7DD",
    x"3046AA34",
    x"30465CA8",
    x"30460F3B",
    x"3045C1EC",
    x"304574BC",
    x"304527A9",
    x"3044DAB5",
    x"30448DDE",
    x"30444126",
    x"3043F48B",
    x"3043A80F",
    x"30435BB0",
    x"30430F6F",
    x"3042C34C",
    x"30427746",
    x"30422B5F",
    x"3041DF95",
    x"304193E8",
    x"30414859",
    x"3040FCE7",
    x"3040B193",
    x"3040665D",
    x"30401B43",
    x"303FD047",
    x"303F8569",
    x"303F3AA7",
    x"303EF003",
    x"303EA57C",
    x"303E5B12",
    x"303E10C4",
    x"303DC694",
    x"303D7C81",
    x"303D328B",
    x"303CE8B2",
    x"303C9EF5",
    x"303C5556",
    x"303C0BD3",
    x"303BC26C",
    x"303B7923",
    x"303B2FF6",
    x"303AE6E5",
    x"303A9DF1",
    x"303A551A",
    x"303A0C5F",
    x"3039C3C0",
    x"30397B3E",
    x"303932D8",
    x"3038EA8E",
    x"3038A261",
    x"30385A4F",
    x"3038125A",
    x"3037CA81",
    x"303782C4",
    x"30373B23",
    x"3036F39E",
    x"3036AC34",
    x"303664E7",
    x"30361DB6",
    x"3035D6A0",
    x"30358FA6",
    x"303548C8",
    x"30350205",
    x"3034BB5E",
    x"303474D3",
    x"30342E63",
    x"3033E80E",
    x"3033A1D5",
    x"30335BB8",
    x"303315B6",
    x"3032CFCF",
    x"30328A03",
    x"30324453",
    x"3031FEBE",
    x"3031B944",
    x"303173E5",
    x"30312EA2",
    x"3030E979",
    x"3030A46B",
    x"30305F78",
    x"30301AA0",
    x"302FD5E4",
    x"302F9141",
    x"302F4CBA",
    x"302F084D",
    x"302EC3FC",
    x"302E7FC4",
    x"302E3BA8",
    x"302DF7A6",
    x"302DB3BE",
    x"302D6FF1",
    x"302D2C3F",
    x"302CE8A7",
    x"302CA529",
    x"302C61C6",
    x"302C1E7D",
    x"302BDB4E",
    x"302B9839",
    x"302B553F",
    x"302B125F",
    x"302ACF98",
    x"302A8CEC",
    x"302A4A5A",
    x"302A07E2",
    x"3029C584",
    x"30298340",
    x"30294116",
    x"3028FF05",
    x"3028BD0E",
    x"30287B31",
    x"3028396E",
    x"3027F7C5",
    x"3027B635",
    x"302774BE",
    x"30273361",
    x"3026F21E",
    x"3026B0F4",
    x"30266FE4",
    x"30262EED",
    x"3025EE0F",
    x"3025AD4B",
    x"30256CA0",
    x"30252C0E",
    x"3024EB95",
    x"3024AB36",
    x"30246AEF",
    x"30242AC2",
    x"3023EAAE",
    x"3023AAB3",
    x"30236AD1",
    x"30232B07",
    x"3022EB57",
    x"3022ABC0",
    x"30226C41",
    x"30222CDB",
    x"3021ED8E",
    x"3021AE59",
    x"30216F3E",
    x"3021303A",
    x"3020F150",
    x"3020B27E",
    x"302073C4",
    x"30203523",
    x"301FF69B",
    x"301FB82B",
    x"301F79D3",
    x"301F3B94",
    x"301EFD6C",
    x"301EBF5E",
    x"301E8167",
    x"301E4389",
    x"301E05C2",
    x"301DC814",
    x"301D8A7E",
    x"301D4D00",
    x"301D0F9A",
    x"301CD24C",
    x"301C9515",
    x"301C57F7",
    x"301C1AF1",
    x"301BDE02",
    x"301BA12B",
    x"301B646C",
    x"301B27C5",
    x"301AEB35",
    x"301AAEBD",
    x"301A725D",
    x"301A3614",
    x"3019F9E2",
    x"3019BDC8",
    x"301981C6",
    x"301945DB",
    x"30190A07",
    x"3018CE4B",
    x"301892A6",
    x"30185719",
    x"30181BA2",
    x"3017E043",
    x"3017A4FB",
    x"301769CA",
    x"30172EB0",
    x"3016F3AE",
    x"3016B8C2",
    x"30167DED",
    x"3016432F",
    x"30160889",
    x"3015CDF9",
    x"30159380",
    x"3015591E",
    x"30151ED2",
    x"3014E49D",
    x"3014AA80",
    x"30147078",
    x"30143688",
    x"3013FCAE",
    x"3013C2EA",
    x"3013893D",
    x"30134FA7",
    x"30131627",
    x"3012DCBE",
    x"3012A36B",
    x"30126A2E",
    x"30123108",
    x"3011F7F8",
    x"3011BEFE",
    x"3011861A",
    x"30114D4D",
    x"30111496",
    x"3010DBF5",
    x"3010A36A",
    x"30106AF5",
    x"30103297",
    x"300FFA4E",
    x"300FC21B",
    x"300F89FE",
    x"300F51F7",
    x"300F1A06",
    x"300EE22B",
    x"300EAA65",
    x"300E72B6",
    x"300E3B1C",
    x"300E0398",
    x"300DCC29",
    x"300D94D0",
    x"300D5D8D",
    x"300D265F",
    x"300CEF47",
    x"300CB844",
    x"300C8157",
    x"300C4A7F",
    x"300C13BD",
    x"300BDD10",
    x"300BA678",
    x"300B6FF5",
    x"300B3988",
    x"300B0331",
    x"300ACCEE",
    x"300A96C0",
    x"300A60A8",
    x"300A2AA5",
    x"3009F4B7",
    x"3009BEDE",
    x"3009891A",
    x"3009536B",
    x"30091DD0",
    x"3008E84B",
    x"3008B2DB",
    x"30087D80",
    x"30084839",
    x"30081307",
    x"3007DDEA",
    x"3007A8E2",
    x"300773EE",
    x"30073F0F",
    x"30070A45",
    x"3006D58F",
    x"3006A0EE",
    x"30066C61",
    x"300637E9",
    x"30060386",
    x"3005CF37",
    x"30059AFC",
    x"300566D5",
    x"300532C3",
    x"3004FEC6",
    x"3004CADC",
    x"30049707",
    x"30046346",
    x"30042F9A",
    x"3003FC01",
    x"3003C87D",
    x"3003950D",
    x"300361B0",
    x"30032E68",
    x"3002FB34",
    x"3002C814",
    x"30029508",
    x"30026210",
    x"30022F2B",
    x"3001FC5B",
    x"3001C99E",
    x"300196F5",
    x"30016460",
    x"300131DF",
    x"3000FF71",
    x"3000CD17",
    x"30009AD1",
    x"3000689E",
    x"3000367F",
    x"30000474",
    x"2FFFA4F7",
    x"2FFF412E",
    x"2FFEDD8C",
    x"2FFE7A11",
    x"2FFE16BD",
    x"2FFDB38F",
    x"2FFD5089",
    x"2FFCEDA8",
    x"2FFC8AEF",
    x"2FFC285C",
    x"2FFBC5EF",
    x"2FFB63A9",
    x"2FFB0189",
    x"2FFA9F90",
    x"2FFA3DBD",
    x"2FF9DC10",
    x"2FF97A89",
    x"2FF91928",
    x"2FF8B7ED",
    x"2FF856D8",
    x"2FF7F5E9",
    x"2FF79520",
    x"2FF7347D",
    x"2FF6D3FF",
    x"2FF673A7",
    x"2FF61375",
    x"2FF5B368",
    x"2FF55381",
    x"2FF4F3BF",
    x"2FF49422",
    x"2FF434AB",
    x"2FF3D559",
    x"2FF3762C",
    x"2FF31725",
    x"2FF2B842",
    x"2FF25985",
    x"2FF1FAEC",
    x"2FF19C79",
    x"2FF13E2A",
    x"2FF0E000",
    x"2FF081FB",
    x"2FF0241A",
    x"2FEFC65F",
    x"2FEF68C7",
    x"2FEF0B55",
    x"2FEEAE07",
    x"2FEE50DD",
    x"2FEDF3D7",
    x"2FED96F6",
    x"2FED3A39",
    x"2FECDDA1",
    x"2FEC812C",
    x"2FEC24DC",
    x"2FEBC8AF",
    x"2FEB6CA7",
    x"2FEB10C3",
    x"2FEAB502",
    x"2FEA5965",
    x"2FE9FDEC",
    x"2FE9A297",
    x"2FE94765",
    x"2FE8EC57",
    x"2FE8916C",
    x"2FE836A5",
    x"2FE7DC02",
    x"2FE78181",
    x"2FE72724",
    x"2FE6CCEB",
    x"2FE672D4",
    x"2FE618E1",
    x"2FE5BF11",
    x"2FE56564",
    x"2FE50BDA",
    x"2FE4B273",
    x"2FE4592E",
    x"2FE4000D",
    x"2FE3A70E",
    x"2FE34E32",
    x"2FE2F579",
    x"2FE29CE3",
    x"2FE2446E",
    x"2FE1EC1D",
    x"2FE193EE",
    x"2FE13BE1",
    x"2FE0E3F7",
    x"2FE08C2F",
    x"2FE0348A",
    x"2FDFDD06",
    x"2FDF85A5",
    x"2FDF2E66",
    x"2FDED749",
    x"2FDE804E",
    x"2FDE2974",
    x"2FDDD2BD",
    x"2FDD7C28",
    x"2FDD25B4",
    x"2FDCCF62",
    x"2FDC7932",
    x"2FDC2324",
    x"2FDBCD37",
    x"2FDB776B",
    x"2FDB21C1",
    x"2FDACC39",
    x"2FDA76D2",
    x"2FDA218C",
    x"2FD9CC68",
    x"2FD97764",
    x"2FD92282",
    x"2FD8CDC1",
    x"2FD87922",
    x"2FD824A3",
    x"2FD7D045",
    x"2FD77C08",
    x"2FD727EC",
    x"2FD6D3F1",
    x"2FD68016",
    x"2FD62C5D",
    x"2FD5D8C4",
    x"2FD5854B",
    x"2FD531F4",
    x"2FD4DEBC",
    x"2FD48BA6",
    x"2FD438AF",
    x"2FD3E5D9",
    x"2FD39324",
    x"2FD3408E",
    x"2FD2EE19",
    x"2FD29BC4",
    x"2FD2498F",
    x"2FD1F77B",
    x"2FD1A586",
    x"2FD153B1",
    x"2FD101FD",
    x"2FD0B068",
    x"2FD05EF3",
    x"2FD00D9E",
    x"2FCFBC68",
    x"2FCF6B52",
    x"2FCF1A5C",
    x"2FCEC986",
    x"2FCE78CF",
    x"2FCE2837",
    x"2FCDD7BF",
    x"2FCD8767",
    x"2FCD372E",
    x"2FCCE714",
    x"2FCC9719",
    x"2FCC473E",
    x"2FCBF781",
    x"2FCBA7E4",
    x"2FCB5866",
    x"2FCB0907",
    x"2FCAB9C7",
    x"2FCA6AA6",
    x"2FCA1BA4",
    x"2FC9CCC0",
    x"2FC97DFC",
    x"2FC92F56",
    x"2FC8E0CF",
    x"2FC89266",
    x"2FC8441C",
    x"2FC7F5F1",
    x"2FC7A7E4",
    x"2FC759F6",
    x"2FC70C26",
    x"2FC6BE74",
    x"2FC670E1",
    x"2FC6236C",
    x"2FC5D616",
    x"2FC588DD",
    x"2FC53BC3",
    x"2FC4EEC6",
    x"2FC4A1E8",
    x"2FC45528",
    x"2FC40885",
    x"2FC3BC01",
    x"2FC36F9B",
    x"2FC32352",
    x"2FC2D727",
    x"2FC28B1A",
    x"2FC23F2A",
    x"2FC1F358",
    x"2FC1A7A4",
    x"2FC15C0D",
    x"2FC11094",
    x"2FC0C538",
    x"2FC079FA",
    x"2FC02ED9",
    x"2FBFE3D6",
    x"2FBF98EF",
    x"2FBF4E26",
    x"2FBF037A",
    x"2FBEB8EB",
    x"2FBE6E7A",
    x"2FBE2425",
    x"2FBDD9ED",
    x"2FBD8FD3",
    x"2FBD45D5",
    x"2FBCFBF4",
    x"2FBCB230",
    x"2FBC6889",
    x"2FBC1EFE",
    x"2FBBD591",
    x"2FBB8C40",
    x"2FBB430B",
    x"2FBAF9F3",
    x"2FBAB0F8",
    x"2FBA6819",
    x"2FBA1F56",
    x"2FB9D6B0",
    x"2FB98E27",
    x"2FB945B9",
    x"2FB8FD68",
    x"2FB8B533",
    x"2FB86D1B",
    x"2FB8251E",
    x"2FB7DD3E",
    x"2FB79579",
    x"2FB74DD1",
    x"2FB70644",
    x"2FB6BED4",
    x"2FB6777F",
    x"2FB63047",
    x"2FB5E92A",
    x"2FB5A228",
    x"2FB55B43",
    x"2FB51479",
    x"2FB4CDCB",
    x"2FB48738",
    x"2FB440C1",
    x"2FB3FA66",
    x"2FB3B426",
    x"2FB36E01",
    x"2FB327F8",
    x"2FB2E20A",
    x"2FB29C37",
    x"2FB25680",
    x"2FB210E3",
    x"2FB1CB62",
    x"2FB185FD",
    x"2FB140B2",
    x"2FB0FB82",
    x"2FB0B66D",
    x"2FB07173",
    x"2FB02C95",
    x"2FAFE7D1",
    x"2FAFA327",
    x"2FAF5E99",
    x"2FAF1A26",
    x"2FAED5CD",
    x"2FAE918F",
    x"2FAE4D6B",
    x"2FAE0962",
    x"2FADC574",
    x"2FAD81A0",
    x"2FAD3DE6",
    x"2FACFA47",
    x"2FACB6C3",
    x"2FAC7359",
    x"2FAC3009",
    x"2FABECD3",
    x"2FABA9B8",
    x"2FAB66B6",
    x"2FAB23CF",
    x"2FAAE102",
    x"2FAA9E50",
    x"2FAA5BB7",
    x"2FAA1938",
    x"2FA9D6D3",
    x"2FA99488",
    x"2FA95257",
    x"2FA91040",
    x"2FA8CE42",
    x"2FA88C5F",
    x"2FA84A95",
    x"2FA808E4",
    x"2FA7C74E",
    x"2FA785D1",
    x"2FA7446D",
    x"2FA70323",
    x"2FA6C1F3",
    x"2FA680DC",
    x"2FA63FDE",
    x"2FA5FEFA",
    x"2FA5BE2F",
    x"2FA57D7D",
    x"2FA53CE5",
    x"2FA4FC65",
    x"2FA4BBFF",
    x"2FA47BB3",
    x"2FA43B7F",
    x"2FA3FB64",
    x"2FA3BB62",
    x"2FA37B7A",
    x"2FA33BAA",
    x"2FA2FBF3",
    x"2FA2BC55",
    x"2FA27CD0",
    x"2FA23D64",
    x"2FA1FE10",
    x"2FA1BED5",
    x"2FA17FB3",
    x"2FA140A9",
    x"2FA101B8",
    x"2FA0C2E0",
    x"2FA08420",
    x"2FA04579",
    x"2FA006EA",
    x"2F9FC873",
    x"2F9F8A15",
    x"2F9F4BCF",
    x"2F9F0DA2",
    x"2F9ECF8D",
    x"2F9E9190",
    x"2F9E53AB",
    x"2F9E15DE",
    x"2F9DD82A",
    x"2F9D9A8E",
    x"2F9D5D09",
    x"2F9D1F9D",
    x"2F9CE248",
    x"2F9CA50C",
    x"2F9C67E7",
    x"2F9C2ADB",
    x"2F9BEDE6",
    x"2F9BB109",
    x"2F9B7444",
    x"2F9B3796",
    x"2F9AFB00",
    x"2F9ABE82",
    x"2F9A821B",
    x"2F9A45CC",
    x"2F9A0995",
    x"2F99CD75",
    x"2F99916C",
    x"2F99557B",
    x"2F9919A2",
    x"2F98DDDF",
    x"2F98A234",
    x"2F9866A0",
    x"2F982B24",
    x"2F97EFBF",
    x"2F97B471",
    x"2F97793A",
    x"2F973E1A",
    x"2F970311",
    x"2F96C820",
    x"2F968D45",
    x"2F965281",
    x"2F9617D4",
    x"2F95DD3F",
    x"2F95A2C0",
    x"2F956857",
    x"2F952E06",
    x"2F94F3CB",
    x"2F94B9A8",
    x"2F947F9A",
    x"2F9445A4",
    x"2F940BC4",
    x"2F93D1FB",
    x"2F939848",
    x"2F935EAC",
    x"2F932526",
    x"2F92EBB7",
    x"2F92B25E",
    x"2F92791B",
    x"2F923FEF",
    x"2F9206D9",
    x"2F91CDDA",
    x"2F9194F0",
    x"2F915C1D",
    x"2F912360",
    x"2F90EABA",
    x"2F90B229",
    x"2F9079AF",
    x"2F90414A",
    x"2F9008FC",
    x"2F8FD0C3",
    x"2F8F98A0",
    x"2F8F6094",
    x"2F8F289D",
    x"2F8EF0BC",
    x"2F8EB8F1",
    x"2F8E813C",
    x"2F8E499C",
    x"2F8E1212",
    x"2F8DDA9E",
    x"2F8DA33F",
    x"2F8D6BF6",
    x"2F8D34C3",
    x"2F8CFDA5",
    x"2F8CC69D",
    x"2F8C8FAA",
    x"2F8C58CC",
    x"2F8C2204",
    x"2F8BEB52",
    x"2F8BB4B5",
    x"2F8B7E2D",
    x"2F8B47BA",
    x"2F8B115D",
    x"2F8ADB14",
    x"2F8AA4E1",
    x"2F8A6EC4",
    x"2F8A38BB",
    x"2F8A02C7",
    x"2F89CCE9",
    x"2F89971F",
    x"2F89616B",
    x"2F892BCB",
    x"2F88F640",
    x"2F88C0CB",
    x"2F888B6A",
    x"2F88561E",
    x"2F8820E6",
    x"2F87EBC4",
    x"2F87B6B6",
    x"2F8781BD",
    x"2F874CD9",
    x"2F871809",
    x"2F86E34E",
    x"2F86AEA8",
    x"2F867A16",
    x"2F864598",
    x"2F86112F",
    x"2F85DCDB",
    x"2F85A89B",
    x"2F85746F",
    x"2F854058",
    x"2F850C55",
    x"2F84D866",
    x"2F84A48C",
    x"2F8470C6",
    x"2F843D14",
    x"2F840976",
    x"2F83D5EC",
    x"2F83A277",
    x"2F836F15",
    x"2F833BC8",
    x"2F83088F",
    x"2F82D569",
    x"2F82A258",
    x"2F826F5A",
    x"2F823C71",
    x"2F82099B",
    x"2F81D6D9",
    x"2F81A42B",
    x"2F817191",
    x"2F813F0B",
    x"2F810C98",
    x"2F80DA39",
    x"2F80A7ED",
    x"2F8075B5",
    x"2F804391",
    x"2F801181",
    x"2F7FBF07",
    x"2F7F5B34",
    x"2F7EF788",
    x"2F7E9403",
    x"2F7E30A4",
    x"2F7DCD6D",
    x"2F7D6A5C",
    x"2F7D0772",
    x"2F7CA4AE",
    x"2F7C4211",
    x"2F7BDF9A",
    x"2F7B7D4A",
    x"2F7B1B20",
    x"2F7AB91D",
    x"2F7A5740",
    x"2F79F589",
    x"2F7993F8",
    x"2F79328D",
    x"2F78D148",
    x"2F78702A",
    x"2F780F31",
    x"2F77AE5E",
    x"2F774DB1",
    x"2F76ED29",
    x"2F768CC7",
    x"2F762C8B",
    x"2F75CC74",
    x"2F756C83",
    x"2F750CB8",
    x"2F74AD11",
    x"2F744D90",
    x"2F73EE35",
    x"2F738EFE",
    x"2F732FED",
    x"2F72D101",
    x"2F72723A",
    x"2F721398",
    x"2F71B51A",
    x"2F7156C2",
    x"2F70F88F",
    x"2F709A80",
    x"2F703C96",
    x"2F6FDED1",
    x"2F6F8130",
    x"2F6F23B4",
    x"2F6EC65C",
    x"2F6E6929",
    x"2F6E0C1A",
    x"2F6DAF2F",
    x"2F6D5269",
    x"2F6CF5C7",
    x"2F6C9949",
    x"2F6C3CEF",
    x"2F6BE0B9",
    x"2F6B84A7",
    x"2F6B28B9",
    x"2F6ACCF0",
    x"2F6A7149",
    x"2F6A15C7",
    x"2F69BA68",
    x"2F695F2D",
    x"2F690416",
    x"2F68A922",
    x"2F684E52",
    x"2F67F3A5",
    x"2F67991B",
    x"2F673EB5",
    x"2F66E472",
    x"2F668A53",
    x"2F663056",
    x"2F65D67D",
    x"2F657CC7",
    x"2F652334",
    x"2F64C9C3",
    x"2F647076",
    x"2F64174B",
    x"2F63BE44",
    x"2F63655F",
    x"2F630C9C",
    x"2F62B3FD",
    x"2F625B80",
    x"2F620325",
    x"2F61AAED",
    x"2F6152D8",
    x"2F60FAE5",
    x"2F60A314",
    x"2F604B65",
    x"2F5FF3D9",
    x"2F5F9C6F",
    x"2F5F4527",
    x"2F5EEE01",
    x"2F5E96FD",
    x"2F5E401B",
    x"2F5DE95B",
    x"2F5D92BC",
    x"2F5D3C40",
    x"2F5CE5E5",
    x"2F5C8FAC",
    x"2F5C3995",
    x"2F5BE39F",
    x"2F5B8DCB",
    x"2F5B3818",
    x"2F5AE287",
    x"2F5A8D17",
    x"2F5A37C9",
    x"2F59E29C",
    x"2F598D90",
    x"2F5938A5",
    x"2F58E3DC",
    x"2F588F33",
    x"2F583AAC",
    x"2F57E645",
    x"2F579200",
    x"2F573DDB",
    x"2F56E9D8",
    x"2F5695F5",
    x"2F564232",
    x"2F55EE91",
    x"2F559B10",
    x"2F5547B0",
    x"2F54F470",
    x"2F54A151",
    x"2F544E52",
    x"2F53FB74",
    x"2F53A8B5",
    x"2F535618",
    x"2F53039A",
    x"2F52B13D",
    x"2F525F00",
    x"2F520CE3",
    x"2F51BAE6",
    x"2F516909",
    x"2F51174C",
    x"2F50C5AE",
    x"2F507431",
    x"2F5022D4",
    x"2F4FD196",
    x"2F4F8078",
    x"2F4F2F79",
    x"2F4EDE9B",
    x"2F4E8DDC",
    x"2F4E3D3C",
    x"2F4DECBC",
    x"2F4D9C5B",
    x"2F4D4C1A",
    x"2F4CFBF7",
    x"2F4CABF5",
    x"2F4C5C11",
    x"2F4C0C4D",
    x"2F4BBCA7",
    x"2F4B6D21",
    x"2F4B1DBA",
    x"2F4ACE72",
    x"2F4A7F49",
    x"2F4A303F",
    x"2F49E153",
    x"2F499287",
    x"2F4943D9",
    x"2F48F54A",
    x"2F48A6D9",
    x"2F485887",
    x"2F480A54",
    x"2F47BC3F",
    x"2F476E49",
    x"2F472071",
    x"2F46D2B7",
    x"2F46851C",
    x"2F46379F",
    x"2F45EA41",
    x"2F459D00",
    x"2F454FDE",
    x"2F4502DA",
    x"2F44B5F4",
    x"2F44692C",
    x"2F441C82",
    x"2F43CFF6",
    x"2F438387",
    x"2F433737",
    x"2F42EB04",
    x"2F429EEF",
    x"2F4252F8",
    x"2F42071E",
    x"2F41BB62",
    x"2F416FC4",
    x"2F412443",
    x"2F40D8E0",
    x"2F408D9A",
    x"2F404271",
    x"2F3FF766",
    x"2F3FAC78",
    x"2F3F61A7",
    x"2F3F16F3",
    x"2F3ECC5D",
    x"2F3E81E4",
    x"2F3E3787",
    x"2F3DED48",
    x"2F3DA326",
    x"2F3D5921",
    x"2F3D0F38",
    x"2F3CC56D",
    x"2F3C7BBE",
    x"2F3C322C",
    x"2F3BE8B7",
    x"2F3B9F5E",
    x"2F3B5622",
    x"2F3B0D03",
    x"2F3AC400",
    x"2F3A7B1A",
    x"2F3A3250",
    x"2F39E9A3",
    x"2F39A112",
    x"2F39589D",
    x"2F391044",
    x"2F38C808",
    x"2F387FE8",
    x"2F3837E4",
    x"2F37EFFC",
    x"2F37A831",
    x"2F376081",
    x"2F3718ED",
    x"2F36D175",
    x"2F368A1A",
    x"2F3642D9",
    x"2F35FBB5",
    x"2F35B4AD",
    x"2F356DC0",
    x"2F3526EF",
    x"2F34E03A",
    x"2F3499A0",
    x"2F345322",
    x"2F340CBF",
    x"2F33C678",
    x"2F33804C",
    x"2F333A3B",
    x"2F32F446",
    x"2F32AE6D",
    x"2F3268AE",
    x"2F32230B",
    x"2F31DD83",
    x"2F319816",
    x"2F3152C4",
    x"2F310D8D",
    x"2F30C871",
    x"2F308370",
    x"2F303E8B",
    x"2F2FF9C0",
    x"2F2FB50F",
    x"2F2F707A",
    x"2F2F2C00",
    x"2F2EE7A0",
    x"2F2EA35B",
    x"2F2E5F30",
    x"2F2E1B20",
    x"2F2DD72B",
    x"2F2D9350",
    x"2F2D4F90",
    x"2F2D0BEA",
    x"2F2CC85E",
    x"2F2C84ED",
    x"2F2C4197",
    x"2F2BFE5A",
    x"2F2BBB38",
    x"2F2B7830",
    x"2F2B3542",
    x"2F2AF26E",
    x"2F2AAFB5",
    x"2F2A6D15",
    x"2F2A2A8F",
    x"2F29E824",
    x"2F29A5D2",
    x"2F29639A",
    x"2F29217C",
    x"2F28DF78",
    x"2F289D8D",
    x"2F285BBD",
    x"2F281A06",
    x"2F27D868",
    x"2F2796E5",
    x"2F27557B",
    x"2F27142A",
    x"2F26D2F3",
    x"2F2691D5",
    x"2F2650D1",
    x"2F260FE6",
    x"2F25CF14",
    x"2F258E5C",
    x"2F254DBD",
    x"2F250D37",
    x"2F24CCCB",
    x"2F248C77",
    x"2F244C3D",
    x"2F240C1C",
    x"2F23CC14",
    x"2F238C24",
    x"2F234C4E",
    x"2F230C91",
    x"2F22CCEC",
    x"2F228D61",
    x"2F224DEE",
    x"2F220E94",
    x"2F21CF52",
    x"2F21902A",
    x"2F21511A",
    x"2F211222",
    x"2F20D344",
    x"2F20947D",
    x"2F2055D0",
    x"2F20173A",
    x"2F1FD8BD",
    x"2F1F9A59",
    x"2F1F5C0D",
    x"2F1F1DD9",
    x"2F1EDFBE",
    x"2F1EA1BA",
    x"2F1E63CF",
    x"2F1E25FC",
    x"2F1DE841",
    x"2F1DAA9F",
    x"2F1D6D14",
    x"2F1D2FA2",
    x"2F1CF247",
    x"2F1CB504",
    x"2F1C77D9",
    x"2F1C3AC7",
    x"2F1BFDCC",
    x"2F1BC0E8",
    x"2F1B841D",
    x"2F1B4769",
    x"2F1B0ACD",
    x"2F1ACE49",
    x"2F1A91DC",
    x"2F1A5587",
    x"2F1A1949",
    x"2F19DD23",
    x"2F19A114",
    x"2F19651D",
    x"2F19293D",
    x"2F18ED75",
    x"2F18B1C4",
    x"2F18762A",
    x"2F183AA7",
    x"2F17FF3C",
    x"2F17C3E8",
    x"2F1788AB",
    x"2F174D85",
    x"2F171276",
    x"2F16D77F",
    x"2F169C9E",
    x"2F1661D4",
    x"2F162722",
    x"2F15EC86",
    x"2F15B201",
    x"2F157793",
    x"2F153D3B",
    x"2F1502FB",
    x"2F14C8D1",
    x"2F148EBE",
    x"2F1454C2",
    x"2F141ADC",
    x"2F13E10D",
    x"2F13A754",
    x"2F136DB2",
    x"2F133426",
    x"2F12FAB1",
    x"2F12C152",
    x"2F12880A",
    x"2F124ED8",
    x"2F1215BC",
    x"2F11DCB7",
    x"2F11A3C8",
    x"2F116AEF",
    x"2F11322C",
    x"2F10F980",
    x"2F10C0E9",
    x"2F108869",
    x"2F104FFF",
    x"2F1017AB",
    x"2F0FDF6C",
    x"2F0FA744",
    x"2F0F6F32",
    x"2F0F3735",
    x"2F0EFF4F",
    x"2F0EC77E",
    x"2F0E8FC3",
    x"2F0E581D",
    x"2F0E208E",
    x"2F0DE914",
    x"2F0DB1B0",
    x"2F0D7A61",
    x"2F0D4328",
    x"2F0D0C05",
    x"2F0CD4F7",
    x"2F0C9DFE",
    x"2F0C671B",
    x"2F0C304E",
    x"2F0BF996",
    x"2F0BC2F3",
    x"2F0B8C65",
    x"2F0B55ED",
    x"2F0B1F8A",
    x"2F0AE93C",
    x"2F0AB304",
    x"2F0A7CE1",
    x"2F0A46D2",
    x"2F0A10D9",
    x"2F09DAF5",
    x"2F09A526",
    x"2F096F6C",
    x"2F0939C7",
    x"2F090437",
    x"2F08CEBC",
    x"2F089955",
    x"2F086404",
    x"2F082EC7",
    x"2F07F99F",
    x"2F07C48C",
    x"2F078F8E",
    x"2F075AA4",
    x"2F0725CF",
    x"2F06F10F",
    x"2F06BC63",
    x"2F0687CB",
    x"2F065349",
    x"2F061EDA",
    x"2F05EA80",
    x"2F05B63B",
    x"2F05820A",
    x"2F054DED",
    x"2F0519E5",
    x"2F04E5F1",
    x"2F04B212",
    x"2F047E46",
    x"2F044A8F",
    x"2F0416EC",
    x"2F03E35D",
    x"2F03AFE2",
    x"2F037C7C",
    x"2F034929",
    x"2F0315EA",
    x"2F02E2C0",
    x"2F02AFA9",
    x"2F027CA7",
    x"2F0249B8",
    x"2F0216DD",
    x"2F01E416",
    x"2F01B163",
    x"2F017EC3",
    x"2F014C38",
    x"2F0119C0",
    x"2F00E75C",
    x"2F00B50B",
    x"2F0082CE",
    x"2F0050A5",
    x"2F001E8F",
    x"2EFFD91A",
    x"2EFF753D",
    x"2EFF1186",
    x"2EFEADF7",
    x"2EFE4A8E",
    x"2EFDE74D",
    x"2EFD8432",
    x"2EFD213D",
    x"2EFCBE70",
    x"2EFC5BC9",
    x"2EFBF948",
    x"2EFB96EE",
    x"2EFB34BA",
    x"2EFAD2AD",
    x"2EFA70C5",
    x"2EFA0F04",
    x"2EF9AD6A",
    x"2EF94BF5",
    x"2EF8EAA6",
    x"2EF8897E",
    x"2EF8287B",
    x"2EF7C79E",
    x"2EF766E7",
    x"2EF70656",
    x"2EF6A5EA",
    x"2EF645A4",
    x"2EF5E583",
    x"2EF58589",
    x"2EF525B3",
    x"2EF4C603",
    x"2EF46678",
    x"2EF40713",
    x"2EF3A7D3",
    x"2EF348B8",
    x"2EF2E9C2",
    x"2EF28AF1",
    x"2EF22C45",
    x"2EF1CDBF",
    x"2EF16F5D",
    x"2EF11120",
    x"2EF0B307",
    x"2EF05514",
    x"2EEFF745",
    x"2EEF999B",
    x"2EEF3C15",
    x"2EEEDEB4",
    x"2EEE8177",
    x"2EEE245E",
    x"2EEDC76A",
    x"2EED6A9B",
    x"2EED0DEF",
    x"2EECB168",
    x"2EEC5504",
    x"2EEBF8C5",
    x"2EEB9CAA",
    x"2EEB40B3",
    x"2EEAE4E0",
    x"2EEA8930",
    x"2EEA2DA4",
    x"2EE9D23C",
    x"2EE976F8",
    x"2EE91BD7",
    x"2EE8C0DA",
    x"2EE86601",
    x"2EE80B4B",
    x"2EE7B0B8",
    x"2EE75649",
    x"2EE6FBFC",
    x"2EE6A1D4",
    x"2EE647CE",
    x"2EE5EDEC",
    x"2EE5942C",
    x"2EE53A90",
    x"2EE4E116",
    x"2EE487C0",
    x"2EE42E8C",
    x"2EE3D57B",
    x"2EE37C8D",
    x"2EE323C2",
    x"2EE2CB1A",
    x"2EE27293",
    x"2EE21A30",
    x"2EE1C1EF",
    x"2EE169D0",
    x"2EE111D4",
    x"2EE0B9FB",
    x"2EE06243",
    x"2EE00AAE",
    x"2EDFB33B",
    x"2EDF5BEA",
    x"2EDF04BB",
    x"2EDEADAE",
    x"2EDE56C3",
    x"2EDDFFFA",
    x"2EDDA953",
    x"2EDD52CE",
    x"2EDCFC6A",
    x"2EDCA629",
    x"2EDC5009",
    x"2EDBFA0A",
    x"2EDBA42D",
    x"2EDB4E72",
    x"2EDAF8D8",
    x"2EDAA35F",
    x"2EDA4E08",
    x"2ED9F8D2",
    x"2ED9A3BE",
    x"2ED94ECA",
    x"2ED8F9F8",
    x"2ED8A547",
    x"2ED850B7",
    x"2ED7FC48",
    x"2ED7A7FA",
    x"2ED753CD",
    x"2ED6FFC1",
    x"2ED6ABD5",
    x"2ED6580A",
    x"2ED60460",
    x"2ED5B0D7",
    x"2ED55D6E",
    x"2ED50A26",
    x"2ED4B6FE",
    x"2ED463F7",
    x"2ED41110",
    x"2ED3BE4A",
    x"2ED36BA3",
    x"2ED3191D",
    x"2ED2C6B8",
    x"2ED27472",
    x"2ED2224D",
    x"2ED1D047",
    x"2ED17E62",
    x"2ED12C9D",
    x"2ED0DAF7",
    x"2ED08971",
    x"2ED0380C",
    x"2ECFE6C6",
    x"2ECF959F",
    x"2ECF4499",
    x"2ECEF3B2",
    x"2ECEA2EA",
    x"2ECE5242",
    x"2ECE01BA",
    x"2ECDB151",
    x"2ECD6108",
    x"2ECD10DD",
    x"2ECCC0D2",
    x"2ECC70E7",
    x"2ECC211A",
    x"2ECBD16D",
    x"2ECB81DF",
    x"2ECB326F",
    x"2ECAE31F",
    x"2ECA93EE",
    x"2ECA44DC",
    x"2EC9F5E8",
    x"2EC9A713",
    x"2EC9585D",
    x"2EC909C6",
    x"2EC8BB4E",
    x"2EC86CF4",
    x"2EC81EB9",
    x"2EC7D09C",
    x"2EC7829E",
    x"2EC734BE",
    x"2EC6E6FC",
    x"2EC69959",
    x"2EC64BD5",
    x"2EC5FE6E",
    x"2EC5B126",
    x"2EC563FC",
    x"2EC516F0",
    x"2EC4CA02",
    x"2EC47D32",
    x"2EC43080",
    x"2EC3E3EC",
    x"2EC39776",
    x"2EC34B1E",
    x"2EC2FEE3",
    x"2EC2B2C7",
    x"2EC266C8",
    x"2EC21AE6",
    x"2EC1CF23",
    x"2EC1837C",
    x"2EC137F4",
    x"2EC0EC89",
    x"2EC0A13B",
    x"2EC0560B",
    x"2EC00AF8",
    x"2EBFC002",
    x"2EBF752A",
    x"2EBF2A6F",
    x"2EBEDFD1",
    x"2EBE9550",
    x"2EBE4AEC",
    x"2EBE00A5",
    x"2EBDB67B",
    x"2EBD6C6F",
    x"2EBD227F",
    x"2EBCD8AC",
    x"2EBC8EF5",
    x"2EBC455C",
    x"2EBBFBDF",
    x"2EBBB27F",
    x"2EBB693C",
    x"2EBB2015",
    x"2EBAD70B",
    x"2EBA8E1D",
    x"2EBA454C",
    x"2EB9FC97",
    x"2EB9B3FE",
    x"2EB96B82",
    x"2EB92322",
    x"2EB8DADF",
    x"2EB892B7",
    x"2EB84AAC",
    x"2EB802BD",
    x"2EB7BAEA",
    x"2EB77333",
    x"2EB72B98",
    x"2EB6E419",
    x"2EB69CB6",
    x"2EB6556E",
    x"2EB60E43",
    x"2EB5C733",
    x"2EB5803F",
    x"2EB53967",
    x"2EB4F2AA",
    x"2EB4AC09",
    x"2EB46584",
    x"2EB41F1A",
    x"2EB3D8CC",
    x"2EB39299",
    x"2EB34C81",
    x"2EB30685",
    x"2EB2C0A4",
    x"2EB27ADE",
    x"2EB23534",
    x"2EB1EFA5",
    x"2EB1AA31",
    x"2EB164D8",
    x"2EB11F9A",
    x"2EB0DA77",
    x"2EB0956F",
    x"2EB05082",
    x"2EB00BB0",
    x"2EAFC6F9",
    x"2EAF825D",
    x"2EAF3DDB",
    x"2EAEF975",
    x"2EAEB528",
    x"2EAE70F7",
    x"2EAE2CE0",
    x"2EADE8E4",
    x"2EADA502",
    x"2EAD613B",
    x"2EAD1D8E",
    x"2EACD9FC",
    x"2EAC9684",
    x"2EAC5326",
    x"2EAC0FE3",
    x"2EABCCBA",
    x"2EAB89AB",
    x"2EAB46B6",
    x"2EAB03DC",
    x"2EAAC11B",
    x"2EAA7E75",
    x"2EAA3BE8",
    x"2EA9F976",
    x"2EA9B71E",
    x"2EA974DF",
    x"2EA932BA",
    x"2EA8F0AF",
    x"2EA8AEBE",
    x"2EA86CE7",
    x"2EA82B29",
    x"2EA7E985",
    x"2EA7A7FB",
    x"2EA7668A",
    x"2EA72532",
    x"2EA6E3F5",
    x"2EA6A2D0",
    x"2EA661C6",
    x"2EA620D4",
    x"2EA5DFFC",
    x"2EA59F3D",
    x"2EA55E97",
    x"2EA51E0B",
    x"2EA4DD98",
    x"2EA49D3E",
    x"2EA45CFD",
    x"2EA41CD5",
    x"2EA3DCC7",
    x"2EA39CD1",
    x"2EA35CF4",
    x"2EA31D30",
    x"2EA2DD85",
    x"2EA29DF3",
    x"2EA25E7A",
    x"2EA21F19",
    x"2EA1DFD1",
    x"2EA1A0A2",
    x"2EA1618C",
    x"2EA1228E",
    x"2EA0E3A9",
    x"2EA0A4DC",
    x"2EA06628",
    x"2EA0278C",
    x"2E9FE909",
    x"2E9FAA9E",
    x"2E9F6C4C",
    x"2E9F2E12",
    x"2E9EEFF0",
    x"2E9EB1E6",
    x"2E9E73F5",
    x"2E9E361C",
    x"2E9DF85B",
    x"2E9DBAB2",
    x"2E9D7D21",
    x"2E9D3FA8",
    x"2E9D0247",
    x"2E9CC4FE",
    x"2E9C87CD",
    x"2E9C4AB4",
    x"2E9C0DB3",
    x"2E9BD0C9",
    x"2E9B93F8",
    x"2E9B573E",
    x"2E9B1A9B",
    x"2E9ADE11",
    x"2E9AA19E",
    x"2E9A6543",
    x"2E9A28FF",
    x"2E99ECD3",
    x"2E99B0BE",
    x"2E9974C0",
    x"2E9938DB",
    x"2E98FD0C",
    x"2E98C155",
    x"2E9885B5",
    x"2E984A2C",
    x"2E980EBB",
    x"2E97D361",
    x"2E97981E",
    x"2E975CF2",
    x"2E9721DD",
    x"2E96E6E0",
    x"2E96ABF9",
    x"2E967129",
    x"2E963670",
    x"2E95FBCF",
    x"2E95C144",
    x"2E9586D0",
    x"2E954C72",
    x"2E95122C",
    x"2E94D7FC",
    x"2E949DE3",
    x"2E9463E1",
    x"2E9429F5",
    x"2E93F020",
    x"2E93B662",
    x"2E937CBA",
    x"2E934328",
    x"2E9309AD",
    x"2E92D048",
    x"2E9296FA",
    x"2E925DC3",
    x"2E9224A1",
    x"2E91EB96",
    x"2E91B2A1",
    x"2E9179C2",
    x"2E9140FA",
    x"2E910848",
    x"2E90CFAB",
    x"2E909725",
    x"2E905EB5",
    x"2E90265B",
    x"2E8FEE17",
    x"2E8FB5E9",
    x"2E8F7DD1",
    x"2E8F45CF",
    x"2E8F0DE3",
    x"2E8ED60C",
    x"2E8E9E4B",
    x"2E8E66A0",
    x"2E8E2F0B",
    x"2E8DF78C",
    x"2E8DC022",
    x"2E8D88CE",
    x"2E8D518F",
    x"2E8D1A66",
    x"2E8CE352",
    x"2E8CAC54",
    x"2E8C756C",
    x"2E8C3E98",
    x"2E8C07DB",
    x"2E8BD132",
    x"2E8B9A9F",
    x"2E8B6422",
    x"2E8B2DB9",
    x"2E8AF766",
    x"2E8AC128",
    x"2E8A8AFF",
    x"2E8A54EB",
    x"2E8A1EED",
    x"2E89E903",
    x"2E89B32E",
    x"2E897D6F",
    x"2E8947C4",
    x"2E89122F",
    x"2E88DCAE",
    x"2E88A742",
    x"2E8871EC",
    x"2E883CA9",
    x"2E88077C",
    x"2E87D264",
    x"2E879D60",
    x"2E876871",
    x"2E873396",
    x"2E86FED0",
    x"2E86CA1F",
    x"2E869582",
    x"2E8660FA",
    x"2E862C87",
    x"2E85F828",
    x"2E85C3DD",
    x"2E858FA6",
    x"2E855B85",
    x"2E852777",
    x"2E84F37E",
    x"2E84BF99",
    x"2E848BC8",
    x"2E84580C",
    x"2E842463",
    x"2E83F0CF",
    x"2E83BD4F",
    x"2E8389E3",
    x"2E83568B",
    x"2E832348",
    x"2E82F018",
    x"2E82BCFC",
    x"2E8289F4",
    x"2E825700",
    x"2E822420",
    x"2E81F154",
    x"2E81BE9C",
    x"2E818BF7",
    x"2E815966",
    x"2E8126E9",
    x"2E80F480",
    x"2E80C22A",
    x"2E808FE8",
    x"2E805DBA",
    x"2E802B9F",
    x"2E7FF32F",
    x"2E7F8F48",
    x"2E7F2B87",
    x"2E7EC7EE",
    x"2E7E647B",
    x"2E7E012F",
    x"2E7D9E0A",
    x"2E7D3B0C",
    x"2E7CD834",
    x"2E7C7583",
    x"2E7C12F8",
    x"2E7BB094",
    x"2E7B4E56",
    x"2E7AEC3F",
    x"2E7A8A4E",
    x"2E7A2883",
    x"2E79C6DE",
    x"2E79655F",
    x"2E790407",
    x"2E78A2D4",
    x"2E7841C7",
    x"2E77E0E1",
    x"2E778020",
    x"2E771F85",
    x"2E76BF0F",
    x"2E765EBF",
    x"2E75FE95",
    x"2E759E90",
    x"2E753EB1",
    x"2E74DEF7",
    x"2E747F63",
    x"2E741FF4",
    x"2E73C0AA",
    x"2E736185",
    x"2E730286",
    x"2E72A3AB",
    x"2E7244F6",
    x"2E71E665",
    x"2E7187FA",
    x"2E7129B3",
    x"2E70CB91",
    x"2E706D94",
    x"2E700FBC",
    x"2E6FB208",
    x"2E6F5479",
    x"2E6EF70E",
    x"2E6E99C8",
    x"2E6E3CA6",
    x"2E6DDFA8",
    x"2E6D82CF",
    x"2E6D261A",
    x"2E6CC989",
    x"2E6C6D1C",
    x"2E6C10D4",
    x"2E6BB4AF",
    x"2E6B58AF",
    x"2E6AFCD2",
    x"2E6AA119",
    x"2E6A4584",
    x"2E69EA13",
    x"2E698EC5",
    x"2E69339B",
    x"2E68D895",
    x"2E687DB2",
    x"2E6822F3",
    x"2E67C857",
    x"2E676DDE",
    x"2E671389",
    x"2E66B957",
    x"2E665F48",
    x"2E66055C",
    x"2E65AB94",
    x"2E6551EE",
    x"2E64F86C",
    x"2E649F0C",
    x"2E6445D0",
    x"2E63ECB6",
    x"2E6393BF",
    x"2E633AEA",
    x"2E62E239",
    x"2E6289A9",
    x"2E62313D",
    x"2E61D8F3",
    x"2E6180CB",
    x"2E6128C6",
    x"2E60D0E4",
    x"2E607923",
    x"2E602185",
    x"2E5FCA09",
    x"2E5F72AF",
    x"2E5F1B77",
    x"2E5EC462",
    x"2E5E6D6E",
    x"2E5E169C",
    x"2E5DBFEC",
    x"2E5D695E",
    x"2E5D12F2",
    x"2E5CBCA7",
    x"2E5C667E",
    x"2E5C1077",
    x"2E5BBA92",
    x"2E5B64CD",
    x"2E5B0F2B",
    x"2E5AB9AA",
    x"2E5A644A",
    x"2E5A0F0B",
    x"2E59B9EE",
    x"2E5964F2",
    x"2E591017",
    x"2E58BB5D",
    x"2E5866C5",
    x"2E58124D",
    x"2E57BDF6",
    x"2E5769C1",
    x"2E5715AC",
    x"2E56C1B8",
    x"2E566DE4",
    x"2E561A32",
    x"2E55C6A0",
    x"2E55732F",
    x"2E551FDE",
    x"2E54CCAE",
    x"2E54799E",
    x"2E5426AF",
    x"2E53D3E0",
    x"2E538131",
    x"2E532EA3",
    x"2E52DC35",
    x"2E5289E7",
    x"2E5237B9",
    x"2E51E5AB",
    x"2E5193BD",
    x"2E5141F0",
    x"2E50F042",
    x"2E509EB4",
    x"2E504D46",
    x"2E4FFBF8",
    x"2E4FAAC9",
    x"2E4F59BA",
    x"2E4F08CB",
    x"2E4EB7FB",
    x"2E4E674B",
    x"2E4E16BB",
    x"2E4DC649",
    x"2E4D75F8",
    x"2E4D25C5",
    x"2E4CD5B2",
    x"2E4C85BE",
    x"2E4C35EA",
    x"2E4BE634",
    x"2E4B969E",
    x"2E4B4726",
    x"2E4AF7CE",
    x"2E4AA895",
    x"2E4A597A",
    x"2E4A0A7F",
    x"2E49BBA2",
    x"2E496CE4",
    x"2E491E45",
    x"2E48CFC5",
    x"2E488163",
    x"2E483320",
    x"2E47E4FB",
    x"2E4796F5",
    x"2E47490D",
    x"2E46FB44",
    x"2E46AD99",
    x"2E46600C",
    x"2E46129E",
    x"2E45C54D",
    x"2E45781B",
    x"2E452B08",
    x"2E44DE12",
    x"2E44913A",
    x"2E444480",
    x"2E43F7E5",
    x"2E43AB67",
    x"2E435F07",
    x"2E4312C4",
    x"2E42C6A0",
    x"2E427A99",
    x"2E422EB0",
    x"2E41E2E5",
    x"2E419737",
    x"2E414BA7",
    x"2E410034",
    x"2E40B4DE",
    x"2E4069A6",
    x"2E401E8C",
    x"2E3FD38F",
    x"2E3F88AF",
    x"2E3F3DEC",
    x"2E3EF346",
    x"2E3EA8BE",
    x"2E3E5E52",
    x"2E3E1404",
    x"2E3DC9D3",
    x"2E3D7FBE",
    x"2E3D35C7",
    x"2E3CEBEC",
    x"2E3CA22E",
    x"2E3C588E",
    x"2E3C0F09",
    x"2E3BC5A2",
    x"2E3B7C57",
    x"2E3B3329",
    x"2E3AEA17",
    x"2E3AA122",
    x"2E3A5849",
    x"2E3A0F8D",
    x"2E39C6ED",
    x"2E397E69",
    x"2E393602",
    x"2E38EDB7",
    x"2E38A588",
    x"2E385D76",
    x"2E38157F",
    x"2E37CDA5",
    x"2E3785E7",
    x"2E373E44",
    x"2E36F6BE",
    x"2E36AF54",
    x"2E366805",
    x"2E3620D2",
    x"2E35D9BB",
    x"2E3592C0",
    x"2E354BE1",
    x"2E35051D",
    x"2E34BE75",
    x"2E3477E8",
    x"2E343177",
    x"2E33EB21",
    x"2E33A4E7",
    x"2E335EC9",
    x"2E3318C5",
    x"2E32D2DD",
    x"2E328D10",
    x"2E32475F",
    x"2E3201C9",
    x"2E31BC4E",
    x"2E3176EE",
    x"2E3131A9",
    x"2E30EC7F",
    x"2E30A770",
    x"2E30627C",
    x"2E301DA3",
    x"2E2FD8E5",
    x"2E2F9441",
    x"2E2F4FB9",
    x"2E2F0B4B",
    x"2E2EC6F8",
    x"2E2E82C0",
    x"2E2E3EA2",
    x"2E2DFA9F",
    x"2E2DB6B6",
    x"2E2D72E8",
    x"2E2D2F34",
    x"2E2CEB9B",
    x"2E2CA81C",
    x"2E2C64B8",
    x"2E2C216E",
    x"2E2BDE3E",
    x"2E2B9B28",
    x"2E2B582C",
    x"2E2B154B",
    x"2E2AD284",
    x"2E2A8FD7",
    x"2E2A4D43",
    x"2E2A0ACA",
    x"2E29C86B",
    x"2E298626",
    x"2E2943FA",
    x"2E2901E8",
    x"2E28BFF1",
    x"2E287E12",
    x"2E283C4E",
    x"2E27FAA3",
    x"2E27B912",
    x"2E27779B",
    x"2E27363D",
    x"2E26F4F8",
    x"2E26B3CD",
    x"2E2672BC",
    x"2E2631C4",
    x"2E25F0E5",
    x"2E25B020",
    x"2E256F73",
    x"2E252EE0",
    x"2E24EE67",
    x"2E24AE06",
    x"2E246DBF",
    x"2E242D90",
    x"2E23ED7B",
    x"2E23AD7F",
    x"2E236D9C",
    x"2E232DD1",
    x"2E22EE20",
    x"2E22AE87",
    x"2E226F07",
    x"2E222FA0",
    x"2E21F052",
    x"2E21B11D",
    x"2E217200",
    x"2E2132FC",
    x"2E20F410",
    x"2E20B53D",
    x"2E207682",
    x"2E2037E0",
    x"2E1FF957",
    x"2E1FBAE6",
    x"2E1F7C8D",
    x"2E1F3E4C",
    x"2E1F0024",
    x"2E1EC214",
    x"2E1E841C",
    x"2E1E463D",
    x"2E1E0875",
    x"2E1DCAC6",
    x"2E1D8D2F",
    x"2E1D4FB0",
    x"2E1D1249",
    x"2E1CD4FA",
    x"2E1C97C2",
    x"2E1C5AA3",
    x"2E1C1D9C",
    x"2E1BE0AC",
    x"2E1BA3D4",
    x"2E1B6714",
    x"2E1B2A6B",
    x"2E1AEDDB",
    x"2E1AB162",
    x"2E1A7500",
    x"2E1A38B6",
    x"2E19FC84",
    x"2E19C069",
    x"2E198466",
    x"2E194879",
    x"2E190CA5",
    x"2E18D0E8",
    x"2E189542",
    x"2E1859B3",
    x"2E181E3C",
    x"2E17E2DB",
    x"2E17A792",
    x"2E176C60",
    x"2E173146",
    x"2E16F642",
    x"2E16BB55",
    x"2E168080",
    x"2E1645C1",
    x"2E160B19",
    x"2E15D088",
    x"2E15960E",
    x"2E155BAB",
    x"2E15215E",
    x"2E14E729",
    x"2E14AD0A",
    x"2E147302",
    x"2E143910",
    x"2E13FF35",
    x"2E13C571",
    x"2E138BC3",
    x"2E13522B",
    x"2E1318AB",
    x"2E12DF40",
    x"2E12A5EC",
    x"2E126CAF",
    x"2E123387",
    x"2E11FA76",
    x"2E11C17C",
    x"2E118897",
    x"2E114FC9",
    x"2E111711",
    x"2E10DE6F",
    x"2E10A5E3",
    x"2E106D6D",
    x"2E10350D",
    x"2E0FFCC4",
    x"2E0FC490",
    x"2E0F8C72",
    x"2E0F546A",
    x"2E0F1C78",
    x"2E0EE49C",
    x"2E0EACD6",
    x"2E0E7525",
    x"2E0E3D8A",
    x"2E0E0605",
    x"2E0DCE95",
    x"2E0D973B",
    x"2E0D5FF7",
    x"2E0D28C8",
    x"2E0CF1AF",
    x"2E0CBAAC",
    x"2E0C83BD",
    x"2E0C4CE5",
    x"2E0C1621",
    x"2E0BDF73",
    x"2E0BA8DB",
    x"2E0B7257",
    x"2E0B3BE9",
    x"2E0B0591",
    x"2E0ACF4D",
    x"2E0A991F",
    x"2E0A6305",
    x"2E0A2D01",
    x"2E09F712",
    x"2E09C138",
    x"2E098B73",
    x"2E0955C3",
    x"2E092028",
    x"2E08EAA2",
    x"2E08B531",
    x"2E087FD5",
    x"2E084A8D",
    x"2E08155A",
    x"2E07E03C",
    x"2E07AB33",
    x"2E07763F",
    x"2E07415F",
    x"2E070C94",
    x"2E06D7DD",
    x"2E06A33B",
    x"2E066EAD",
    x"2E063A34",
    x"2E0605D0",
    x"2E05D180",
    x"2E059D44",
    x"2E05691D",
    x"2E05350A",
    x"2E05010C",
    x"2E04CD21",
    x"2E04994B",
    x"2E04658A",
    x"2E0431DC",
    x"2E03FE43",
    x"2E03CABD",
    x"2E03974C",
    x"2E0363EF",
    x"2E0330A6",
    x"2E02FD71",
    x"2E02CA50",
    x"2E029743",
    x"2E02644A",
    x"2E023165",
    x"2E01FE93",
    x"2E01CBD6",
    x"2E01992C",
    x"2E016696",
    x"2E013414",
    x"2E0101A5",
    x"2E00CF4B",
    x"2E009D03",
    x"2E006AD0",
    x"2E0038B0",
    x"2E0006A4",
    x"2DFFA956",
    x"2DFF458B",
    x"2DFEE1E7",
    x"2DFE7E6A",
    x"2DFE1B14",
    x"2DFDB7E5",
    x"2DFD54DD",
    x"2DFCF1FB",
    x"2DFC8F40",
    x"2DFC2CAB",
    x"2DFBCA3D",
    x"2DFB67F5",
    x"2DFB05D4",
    x"2DFAA3D8",
    x"2DFA4204",
    x"2DF9E055",
    x"2DF97ECC",
    x"2DF91D6A",
    x"2DF8BC2D",
    x"2DF85B17",
    x"2DF7FA26",
    x"2DF7995B",
    x"2DF738B6",
    x"2DF6D837",
    x"2DF677DD",
    x"2DF617A9",
    x"2DF5B79B",
    x"2DF557B2",
    x"2DF4F7EE",
    x"2DF49850",
    x"2DF438D7",
    x"2DF3D984",
    x"2DF37A55",
    x"2DF31B4C",
    x"2DF2BC68",
    x"2DF25DA9",
    x"2DF1FF0F",
    x"2DF1A09A",
    x"2DF14249",
    x"2DF0E41E",
    x"2DF08617",
    x"2DF02835",
    x"2DEFCA78",
    x"2DEF6CDF",
    x"2DEF0F6B",
    x"2DEEB21B",
    x"2DEE54EF",
    x"2DEDF7E8",
    x"2DED9B06",
    x"2DED3E47",
    x"2DECE1AD",
    x"2DEC8537",
    x"2DEC28E5",
    x"2DEBCCB7",
    x"2DEB70AD",
    x"2DEB14C7",
    x"2DEAB905",
    x"2DEA5D66",
    x"2DEA01EC",
    x"2DE9A695",
    x"2DE94B62",
    x"2DE8F052",
    x"2DE89566",
    x"2DE83A9D",
    x"2DE7DFF8",
    x"2DE78576",
    x"2DE72B18",
    x"2DE6D0DC",
    x"2DE676C4",
    x"2DE61CD0",
    x"2DE5C2FE",
    x"2DE5694F",
    x"2DE50FC4",
    x"2DE4B65B",
    x"2DE45D15",
    x"2DE403F2",
    x"2DE3AAF2",
    x"2DE35215",
    x"2DE2F95A",
    x"2DE2A0C2",
    x"2DE2484C",
    x"2DE1EFF9",
    x"2DE197C9",
    x"2DE13FBB",
    x"2DE0E7CF",
    x"2DE09006",
    x"2DE0385E",
    x"2DDFE0DA",
    x"2DDF8977",
    x"2DDF3236",
    x"2DDEDB18",
    x"2DDE841B",
    x"2DDE2D40",
    x"2DDDD688",
    x"2DDD7FF1",
    x"2DDD297C",
    x"2DDCD328",
    x"2DDC7CF7",
    x"2DDC26E7",
    x"2DDBD0F8",
    x"2DDB7B2B",
    x"2DDB2580",
    x"2DDACFF6",
    x"2DDA7A8E",
    x"2DDA2546",
    x"2DD9D020",
    x"2DD97B1C",
    x"2DD92638",
    x"2DD8D176",
    x"2DD87CD5",
    x"2DD82854",
    x"2DD7D3F5",
    x"2DD77FB7",
    x"2DD72B99",
    x"2DD6D79D",
    x"2DD683C1",
    x"2DD63006",
    x"2DD5DC6B",
    x"2DD588F1",
    x"2DD53598",
    x"2DD4E260",
    x"2DD48F47",
    x"2DD43C50",
    x"2DD3E978",
    x"2DD396C1",
    x"2DD3442A",
    x"2DD2F1B4",
    x"2DD29F5E",
    x"2DD24D27",
    x"2DD1FB11",
    x"2DD1A91B",
    x"2DD15745",
    x"2DD1058F",
    x"2DD0B3F9",
    x"2DD06282",
    x"2DD0112C",
    x"2DCFBFF5",
    x"2DCF6EDE",
    x"2DCF1DE6",
    x"2DCECD0E",
    x"2DCE7C56",
    x"2DCE2BBD",
    x"2DCDDB44",
    x"2DCD8AEA",
    x"2DCD3AAF",
    x"2DCCEA94",
    x"2DCC9A98",
    x"2DCC4ABB",
    x"2DCBFAFE",
    x"2DCBAB5F",
    x"2DCB5BE0",
    x"2DCB0C7F",
    x"2DCABD3E",
    x"2DCA6E1C",
    x"2DCA1F18",
    x"2DC9D033",
    x"2DC9816D",
    x"2DC932C6",
    x"2DC8E43E",
    x"2DC895D4",
    x"2DC84789",
    x"2DC7F95C",
    x"2DC7AB4E",
    x"2DC75D5E",
    x"2DC70F8D",
    x"2DC6C1DA",
    x"2DC67445",
    x"2DC626CF",
    x"2DC5D977",
    x"2DC58C3D",
    x"2DC53F21",
    x"2DC4F224",
    x"2DC4A544",
    x"2DC45883",
    x"2DC40BDF",
    x"2DC3BF59",
    x"2DC372F2",
    x"2DC326A8",
    x"2DC2DA7B",
    x"2DC28E6D",
    x"2DC2427C",
    x"2DC1F6A9",
    x"2DC1AAF3",
    x"2DC15F5B",
    x"2DC113E1",
    x"2DC0C884",
    x"2DC07D44",
    x"2DC03222",
    x"2DBFE71D",
    x"2DBF9C35",
    x"2DBF516B",
    x"2DBF06BE",
    x"2DBEBC2E",
    x"2DBE71BB",
    x"2DBE2765",
    x"2DBDDD2C",
    x"2DBD9310",
    x"2DBD4911",
    x"2DBCFF2F",
    x"2DBCB56A",
    x"2DBC6BC1",
    x"2DBC2235",
    x"2DBBD8C6",
    x"2DBB8F74",
    x"2DBB463E",
    x"2DBAFD25",
    x"2DBAB429",
    x"2DBA6B48",
    x"2DBA2285",
    x"2DB9D9DD",
    x"2DB99152",
    x"2DB948E4",
    x"2DB90092",
    x"2DB8B85B",
    x"2DB87041",
    x"2DB82844",
    x"2DB7E062",
    x"2DB7989C",
    x"2DB750F3",
    x"2DB70965",
    x"2DB6C1F3",
    x"2DB67A9E",
    x"2DB63364",
    x"2DB5EC45",
    x"2DB5A543",
    x"2DB55E5C",
    x"2DB51791",
    x"2DB4D0E2",
    x"2DB48A4E",
    x"2DB443D6",
    x"2DB3FD79",
    x"2DB3B738",
    x"2DB37112",
    x"2DB32B07",
    x"2DB2E518",
    x"2DB29F44",
    x"2DB2598C",
    x"2DB213EE",
    x"2DB1CE6C",
    x"2DB18905",
    x"2DB143B9",
    x"2DB0FE88",
    x"2DB0B972",
    x"2DB07477",
    x"2DB02F97",
    x"2DAFEAD2",
    x"2DAFA628",
    x"2DAF6198",
    x"2DAF1D24",
    x"2DAED8CA",
    x"2DAE948A",
    x"2DAE5065",
    x"2DAE0C5B",
    x"2DADC86C",
    x"2DAD8497",
    x"2DAD40DC",
    x"2DACFD3C",
    x"2DACB9B6",
    x"2DAC764B",
    x"2DAC32FA",
    x"2DABEFC3",
    x"2DABACA7",
    x"2DAB69A4",
    x"2DAB26BC",
    x"2DAAE3EE",
    x"2DAAA13A",
    x"2DAA5EA0",
    x"2DAA1C20",
    x"2DA9D9BA",
    x"2DA9976E",
    x"2DA9553C",
    x"2DA91323",
    x"2DA8D125",
    x"2DA88F40",
    x"2DA84D75",
    x"2DA80BC3",
    x"2DA7CA2C",
    x"2DA788AD",
    x"2DA74749",
    x"2DA705FE",
    x"2DA6C4CC",
    x"2DA683B4",
    x"2DA642B5",
    x"2DA601D0",
    x"2DA5C104",
    x"2DA58051",
    x"2DA53FB8",
    x"2DA4FF37",
    x"2DA4BED0",
    x"2DA47E82",
    x"2DA43E4D",
    x"2DA3FE31",
    x"2DA3BE2F",
    x"2DA37E45",
    x"2DA33E74",
    x"2DA2FEBC",
    x"2DA2BF1D",
    x"2DA27F97",
    x"2DA24029",
    x"2DA200D5",
    x"2DA1C199",
    x"2DA18275",
    x"2DA1436B",
    x"2DA10479",
    x"2DA0C59F",
    x"2DA086DE",
    x"2DA04836",
    x"2DA009A6",
    x"2D9FCB2E",
    x"2D9F8CCF",
    x"2D9F4E88",
    x"2D9F105A",
    x"2D9ED243",
    x"2D9E9445",
    x"2D9E5660",
    x"2D9E1892",
    x"2D9DDADC",
    x"2D9D9D3F",
    x"2D9D5FBA",
    x"2D9D224C",
    x"2D9CE4F7",
    x"2D9CA7B9",
    x"2D9C6A94",
    x"2D9C2D86",
    x"2D9BF090",
    x"2D9BB3B2",
    x"2D9B76EC",
    x"2D9B3A3D",
    x"2D9AFDA6",
    x"2D9AC127",
    x"2D9A84BF",
    x"2D9A486F",
    x"2D9A0C37",
    x"2D99D016",
    x"2D99940C",
    x"2D99581A",
    x"2D991C3F",
    x"2D98E07C",
    x"2D98A4D0",
    x"2D98693B",
    x"2D982DBE",
    x"2D97F257",
    x"2D97B708",
    x"2D977BD0",
    x"2D9740B0",
    x"2D9705A6",
    x"2D96CAB3",
    x"2D968FD7",
    x"2D965513",
    x"2D961A65",
    x"2D95DFCE",
    x"2D95A54E",
    x"2D956AE5",
    x"2D953093",
    x"2D94F657",
    x"2D94BC32",
    x"2D948224",
    x"2D94482C",
    x"2D940E4C",
    x"2D93D481",
    x"2D939ACE",
    x"2D936130",
    x"2D9327AA",
    x"2D92EE39",
    x"2D92B4DF",
    x"2D927B9C",
    x"2D92426F",
    x"2D920958",
    x"2D91D058",
    x"2D91976D",
    x"2D915E99",
    x"2D9125DB",
    x"2D90ED34",
    x"2D90B4A2",
    x"2D907C27",
    x"2D9043C1",
    x"2D900B72",
    x"2D8FD338",
    x"2D8F9B15",
    x"2D8F6307",
    x"2D8F2B0F",
    x"2D8EF32D",
    x"2D8EBB61",
    x"2D8E83AB",
    x"2D8E4C0A",
    x"2D8E1480",
    x"2D8DDD0A",
    x"2D8DA5AB",
    x"2D8D6E61",
    x"2D8D372D",
    x"2D8D000E",
    x"2D8CC905",
    x"2D8C9211",
    x"2D8C5B32",
    x"2D8C2469",
    x"2D8BEDB6",
    x"2D8BB718",
    x"2D8B808F",
    x"2D8B4A1B",
    x"2D8B13BD",
    x"2D8ADD74",
    x"2D8AA740",
    x"2D8A7121",
    x"2D8A3B18",
    x"2D8A0523",
    x"2D89CF44",
    x"2D899979",
    x"2D8963C4",
    x"2D892E23",
    x"2D88F898",
    x"2D88C321",
    x"2D888DBF",
    x"2D885872",
    x"2D88233A",
    x"2D87EE17",
    x"2D87B908",
    x"2D87840E",
    x"2D874F29",
    x"2D871A58",
    x"2D86E59C",
    x"2D86B0F5",
    x"2D867C62",
    x"2D8647E4",
    x"2D86137A",
    x"2D85DF24",
    x"2D85AAE3",
    x"2D8576B7",
    x"2D85429F",
    x"2D850E9B",
    x"2D84DAAB",
    x"2D84A6D0",
    x"2D847309",
    x"2D843F56",
    x"2D840BB7",
    x"2D83D82D",
    x"2D83A4B7",
    x"2D837154",
    x"2D833E06",
    x"2D830ACC",
    x"2D82D7A6",
    x"2D82A493",
    x"2D827195",
    x"2D823EAB",
    x"2D820BD4",
    x"2D81D911",
    x"2D81A662",
    x"2D8173C7",
    x"2D814140",
    x"2D810ECC",
    x"2D80DC6C",
    x"2D80AA20",
    x"2D8077E7",
    x"2D8045C2",
    x"2D8013B1",
    x"2D7FC366",
    x"2D7F5F91",
    x"2D7EFBE3",
    x"2D7E985C",
    x"2D7E34FC",
    x"2D7DD1C3",
    x"2D7D6EB0",
    x"2D7D0BC4",
    x"2D7CA8FF",
    x"2D7C4660",
    x"2D7BE3E8",
    x"2D7B8196",
    x"2D7B1F6B",
    x"2D7ABD66",
    x"2D7A5B87",
    x"2D79F9CE",
    x"2D79983C",
    x"2D7936CF",
    x"2D78D589",
    x"2D787468",
    x"2D78136E",
    x"2D77B299",
    x"2D7751EA",
    x"2D76F161",
    x"2D7690FE",
    x"2D7630C0",
    x"2D75D0A8",
    x"2D7570B5",
    x"2D7510E8",
    x"2D74B140",
    x"2D7451BD",
    x"2D73F260",
    x"2D739328",
    x"2D733415",
    x"2D72D527",
    x"2D72765E",
    x"2D7217BB",
    x"2D71B93C",
    x"2D715AE2",
    x"2D70FCAD",
    x"2D709E9C",
    x"2D7040B1",
    x"2D6FE2EA",
    x"2D6F8548",
    x"2D6F27CA",
    x"2D6ECA70",
    x"2D6E6D3C",
    x"2D6E102B",
    x"2D6DB33F",
    x"2D6D5677",
    x"2D6CF9D3",
    x"2D6C9D54",
    x"2D6C40F8",
    x"2D6BE4C1",
    x"2D6B88AE",
    x"2D6B2CBE",
    x"2D6AD0F3",
    x"2D6A754B",
    x"2D6A19C7",
    x"2D69BE67",
    x"2D69632A",
    x"2D690811",
    x"2D68AD1C",
    x"2D68524A",
    x"2D67F79C",
    x"2D679D11",
    x"2D6742A9",
    x"2D66E864",
    x"2D668E43",
    x"2D663445",
    x"2D65DA6A",
    x"2D6580B3",
    x"2D65271E",
    x"2D64CDAC",
    x"2D64745D",
    x"2D641B31",
    x"2D63C228",
    x"2D636941",
    x"2D63107E",
    x"2D62B7DD",
    x"2D625F5E",
    x"2D620702",
    x"2D61AEC9",
    x"2D6156B1",
    x"2D60FEBD",
    x"2D60A6EA",
    x"2D604F3A",
    x"2D5FF7AD",
    x"2D5FA041",
    x"2D5F48F7",
    x"2D5EF1D0",
    x"2D5E9ACA",
    x"2D5E43E7",
    x"2D5DED25",
    x"2D5D9686",
    x"2D5D4008",
    x"2D5CE9AC",
    x"2D5C9371",
    x"2D5C3D58",
    x"2D5BE761",
    x"2D5B918C",
    x"2D5B3BD7",
    x"2D5AE645",
    x"2D5A90D4",
    x"2D5A3B84",
    x"2D59E655",
    x"2D599148",
    x"2D593C5C",
    x"2D58E791",
    x"2D5892E7",
    x"2D583E5E",
    x"2D57E9F6",
    x"2D5795AF",
    x"2D574189",
    x"2D56ED84",
    x"2D56999F",
    x"2D5645DC",
    x"2D55F239",
    x"2D559EB6",
    x"2D554B55",
    x"2D54F814",
    x"2D54A4F3",
    x"2D5451F3",
    x"2D53FF13",
    x"2D53AC53",
    x"2D5359B4",
    x"2D530735",
    x"2D52B4D7",
    x"2D526298",
    x"2D52107A",
    x"2D51BE7B",
    x"2D516C9D",
    x"2D511ADE",
    x"2D50C940",
    x"2D5077C1",
    x"2D502662",
    x"2D4FD523",
    x"2D4F8404",
    x"2D4F3304",
    x"2D4EE224",
    x"2D4E9163",
    x"2D4E40C2",
    x"2D4DF041",
    x"2D4D9FDE",
    x"2D4D4F9C",
    x"2D4CFF78",
    x"2D4CAF74",
    x"2D4C5F8F",
    x"2D4C0FC9",
    x"2D4BC023",
    x"2D4B709B",
    x"2D4B2133",
    x"2D4AD1E9",
    x"2D4A82BF",
    x"2D4A33B3",
    x"2D49E4C6",
    x"2D4995F8",
    x"2D494749",
    x"2D48F8B9",
    x"2D48AA47",
    x"2D485BF4",
    x"2D480DBF",
    x"2D47BFA9",
    x"2D4771B1",
    x"2D4723D8",
    x"2D46D61D",
    x"2D468881",
    x"2D463B03",
    x"2D45EDA3",
    x"2D45A061",
    x"2D45533D",
    x"2D450638",
    x"2D44B950",
    x"2D446C87",
    x"2D441FDC",
    x"2D43D34E",
    x"2D4386DF",
    x"2D433A8D",
    x"2D42EE59",
    x"2D42A243",
    x"2D42564A",
    x"2D420A6F",
    x"2D41BEB2",
    x"2D417312",
    x"2D412790",
    x"2D40DC2B",
    x"2D4090E4",
    x"2D4045BA",
    x"2D3FFAAD",
    x"2D3FAFBE",
    x"2D3F64EC",
    x"2D3F1A37",
    x"2D3ECFA0",
    x"2D3E8525",
    x"2D3E3AC8",
    x"2D3DF087",
    x"2D3DA664",
    x"2D3D5C5D",
    x"2D3D1273",
    x"2D3CC8A7",
    x"2D3C7EF7",
    x"2D3C3563",
    x"2D3BEBED",
    x"2D3BA293",
    x"2D3B5956",
    x"2D3B1035",
    x"2D3AC731",
    x"2D3A7E4A",
    x"2D3A357F",
    x"2D39ECD0",
    x"2D39A43E",
    x"2D395BC8",
    x"2D39136E",
    x"2D38CB30",
    x"2D38830F",
    x"2D383B0A",
    x"2D37F321",
    x"2D37AB54",
    x"2D3763A3",
    x"2D371C0E",
    x"2D36D495",
    x"2D368D38",
    x"2D3645F7",
    x"2D35FED1",
    x"2D35B7C8",
    x"2D3570DA",
    x"2D352A08",
    x"2D34E351",
    x"2D349CB6",
    x"2D345636",
    x"2D340FD3",
    x"2D33C98A",
    x"2D33835D",
    x"2D333D4B",
    x"2D32F755",
    x"2D32B17A",
    x"2D326BBB",
    x"2D322616",
    x"2D31E08D",
    x"2D319B1F",
    x"2D3155CC",
    x"2D311094",
    x"2D30CB77",
    x"2D308675",
    x"2D30418E",
    x"2D2FFCC1",
    x"2D2FB810",
    x"2D2F737A",
    x"2D2F2EFE",
    x"2D2EEA9D",
    x"2D2EA657",
    x"2D2E622B",
    x"2D2E1E1A",
    x"2D2DDA23",
    x"2D2D9647",
    x"2D2D5286",
    x"2D2D0EDF",
    x"2D2CCB52",
    x"2D2C87E0",
    x"2D2C4488",
    x"2D2C014A",
    x"2D2BBE27",
    x"2D2B7B1E",
    x"2D2B382F",
    x"2D2AF55A",
    x"2D2AB29F",
    x"2D2A6FFE",
    x"2D2A2D78",
    x"2D29EB0B",
    x"2D29A8B8",
    x"2D29667F",
    x"2D292460",
    x"2D28E25B",
    x"2D28A06F",
    x"2D285E9D",
    x"2D281CE5",
    x"2D27DB47",
    x"2D2799C2",
    x"2D275857",
    x"2D271705",
    x"2D26D5CD",
    x"2D2694AE",
    x"2D2653A8",
    x"2D2612BC",
    x"2D25D1EA",
    x"2D259130",
    x"2D255090",
    x"2D251009",
    x"2D24CF9C",
    x"2D248F47",
    x"2D244F0C",
    x"2D240EE9",
    x"2D23CEE0",
    x"2D238EF0",
    x"2D234F19",
    x"2D230F5A",
    x"2D22CFB4",
    x"2D229028",
    x"2D2250B4",
    x"2D221159",
    x"2D21D216",
    x"2D2192ED",
    x"2D2153DB",
    x"2D2114E3",
    x"2D20D603",
    x"2D20973C",
    x"2D20588D",
    x"2D2019F7",
    x"2D1FDB79",
    x"2D1F9D13",
    x"2D1F5EC6",
    x"2D1F2091",
    x"2D1EE275",
    x"2D1EA470",
    x"2D1E6684",
    x"2D1E28B0",
    x"2D1DEAF4",
    x"2D1DAD51",
    x"2D1D6FC5",
    x"2D1D3251",
    x"2D1CF4F6",
    x"2D1CB7B2",
    x"2D1C7A86",
    x"2D1C3D72",
    x"2D1C0076",
    x"2D1BC392",
    x"2D1B86C5",
    x"2D1B4A10",
    x"2D1B0D73",
    x"2D1AD0EE",
    x"2D1A9480",
    x"2D1A582A",
    x"2D1A1BEB",
    x"2D19DFC4",
    x"2D19A3B4",
    x"2D1967BC",
    x"2D192BDB",
    x"2D18F012",
    x"2D18B460",
    x"2D1878C5",
    x"2D183D41",
    x"2D1801D5",
    x"2D17C680",
    x"2D178B42",
    x"2D17501B",
    x"2D17150B",
    x"2D16DA13",
    x"2D169F31",
    x"2D166466",
    x"2D1629B3",
    x"2D15EF16",
    x"2D15B490",
    x"2D157A21",
    x"2D153FC8",
    x"2D150587",
    x"2D14CB5C",
    x"2D149148",
    x"2D14574A",
    x"2D141D64",
    x"2D13E393",
    x"2D13A9DA",
    x"2D137037",
    x"2D1336AA",
    x"2D12FD34",
    x"2D12C3D4",
    x"2D128A8B",
    x"2D125158",
    x"2D12183B",
    x"2D11DF35",
    x"2D11A645",
    x"2D116D6B",
    x"2D1134A8",
    x"2D10FBFA",
    x"2D10C363",
    x"2D108AE1",
    x"2D105276",
    x"2D101A21",
    x"2D0FE1E2",
    x"2D0FA9B9",
    x"2D0F71A5",
    x"2D0F39A8",
    x"2D0F01C0",
    x"2D0EC9EE",
    x"2D0E9232",
    x"2D0E5A8C",
    x"2D0E22FC",
    x"2D0DEB81",
    x"2D0DB41C",
    x"2D0D7CCC",
    x"2D0D4592",
    x"2D0D0E6E",
    x"2D0CD75F",
    x"2D0CA065",
    x"2D0C6982",
    x"2D0C32B3",
    x"2D0BFBFA",
    x"2D0BC556",
    x"2D0B8EC8",
    x"2D0B584F",
    x"2D0B21EB",
    x"2D0AEB9C",
    x"2D0AB563",
    x"2D0A7F3E",
    x"2D0A492F",
    x"2D0A1335",
    x"2D09DD50",
    x"2D09A780",
    x"2D0971C5",
    x"2D093C1F",
    x"2D09068E",
    x"2D08D112",
    x"2D089BAB",
    x"2D086659",
    x"2D08311B",
    x"2D07FBF2",
    x"2D07C6DE",
    x"2D0791DF",
    x"2D075CF4",
    x"2D07281E",
    x"2D06F35D",
    x"2D06BEB0",
    x"2D068A18",
    x"2D065594",
    x"2D062125",
    x"2D05ECCA",
    x"2D05B884",
    x"2D058452",
    x"2D055035",
    x"2D051C2B",
    x"2D04E837",
    x"2D04B456",
    x"2D04808A",
    x"2D044CD2",
    x"2D04192E",
    x"2D03E59E",
    x"2D03B222",
    x"2D037EBB",
    x"2D034B67",
    x"2D031828",
    x"2D02E4FC",
    x"2D02B1E5",
    x"2D027EE1",
    x"2D024BF2",
    x"2D021916",
    x"2D01E64E",
    x"2D01B39A",
    x"2D0180FA",
    x"2D014E6D",
    x"2D011BF5",
    x"2D00E98F",
    x"2D00B73E",
    x"2D008500",
    x"2D0052D6",
    x"2D0020C0",
    x"2CFFDD79",
    x"2CFF799A",
    x"2CFF15E2",
    x"2CFEB251",
    x"2CFE4EE7",
    x"2CFDEBA3",
    x"2CFD8887",
    x"2CFD2591",
    x"2CFCC2C1",
    x"2CFC6019",
    x"2CFBFD96",
    x"2CFB9B3A",
    x"2CFB3905",
    x"2CFAD6F6",
    x"2CFA750D",
    x"2CFA134A",
    x"2CF9B1AE",
    x"2CF95038",
    x"2CF8EEE7",
    x"2CF88DBD",
    x"2CF82CB8",
    x"2CF7CBDA",
    x"2CF76B21",
    x"2CF70A8E",
    x"2CF6AA21",
    x"2CF649D9",
    x"2CF5E9B7",
    x"2CF589BB",
    x"2CF529E4",
    x"2CF4CA32",
    x"2CF46AA6",
    x"2CF40B3F",
    x"2CF3ABFD",
    x"2CF34CE0",
    x"2CF2EDE9",
    x"2CF28F16",
    x"2CF23069",
    x"2CF1D1E0",
    x"2CF1737D",
    x"2CF1153E",
    x"2CF0B724",
    x"2CF0592F",
    x"2CEFFB5F",
    x"2CEF9DB3",
    x"2CEF402B",
    x"2CEEE2C9",
    x"2CEE858A",
    x"2CEE2870",
    x"2CEDCB7B",
    x"2CED6EA9",
    x"2CED11FC",
    x"2CECB573",
    x"2CEC590E",
    x"2CEBFCCE",
    x"2CEBA0B1",
    x"2CEB44B8",
    x"2CEAE8E3",
    x"2CEA8D32",
    x"2CEA31A5",
    x"2CE9D63B",
    x"2CE97AF5",
    x"2CE91FD3",
    x"2CE8C4D5",
    x"2CE869F9",
    x"2CE80F42",
    x"2CE7B4AD",
    x"2CE75A3D",
    x"2CE6FFEF",
    x"2CE6A5C5",
    x"2CE64BBD",
    x"2CE5F1D9",
    x"2CE59818",
    x"2CE53E7B",
    x"2CE4E500",
    x"2CE48BA8",
    x"2CE43272",
    x"2CE3D960",
    x"2CE38071",
    x"2CE327A4",
    x"2CE2CEFA",
    x"2CE27672",
    x"2CE21E0D",
    x"2CE1C5CB",
    x"2CE16DAB",
    x"2CE115AD",
    x"2CE0BDD2",
    x"2CE06619",
    x"2CE00E82",
    x"2CDFB70D",
    x"2CDF5FBB",
    x"2CDF088A",
    x"2CDEB17C",
    x"2CDE5A90",
    x"2CDE03C5",
    x"2CDDAD1D",
    x"2CDD5696",
    x"2CDD0031",
    x"2CDCA9EE",
    x"2CDC53CC",
    x"2CDBFDCC",
    x"2CDBA7EE",
    x"2CDB5231",
    x"2CDAFC96",
    x"2CDAA71C",
    x"2CDA51C3",
    x"2CD9FC8C",
    x"2CD9A776",
    x"2CD95281",
    x"2CD8FDAD",
    x"2CD8A8FB",
    x"2CD85469",
    x"2CD7FFF9",
    x"2CD7ABA9",
    x"2CD7577B",
    x"2CD7036D",
    x"2CD6AF80",
    x"2CD65BB4",
    x"2CD60808",
    x"2CD5B47E",
    x"2CD56113",
    x"2CD50DCA",
    x"2CD4BAA1",
    x"2CD46798",
    x"2CD414B0",
    x"2CD3C1E8",
    x"2CD36F40",
    x"2CD31CB9",
    x"2CD2CA52",
    x"2CD2780B",
    x"2CD225E4",
    x"2CD1D3DD",
    x"2CD181F6",
    x"2CD13030",
    x"2CD0DE89",
    x"2CD08D02",
    x"2CD03B9B",
    x"2CCFEA53",
    x"2CCF992B",
    x"2CCF4823",
    x"2CCEF73B",
    x"2CCEA672",
    x"2CCE55C9",
    x"2CCE053F",
    x"2CCDB4D5",
    x"2CCD648A",
    x"2CCD145E",
    x"2CCCC452",
    x"2CCC7465",
    x"2CCC2497",
    x"2CCBD4E8",
    x"2CCB8559",
    x"2CCB35E8",
    x"2CCAE697",
    x"2CCA9764",
    x"2CCA4850",
    x"2CC9F95C",
    x"2CC9AA86",
    x"2CC95BCE",
    x"2CC90D36",
    x"2CC8BEBC",
    x"2CC87061",
    x"2CC82224",
    x"2CC7D406",
    x"2CC78606",
    x"2CC73825",
    x"2CC6EA63",
    x"2CC69CBE",
    x"2CC64F38",
    x"2CC601D0",
    x"2CC5B487",
    x"2CC5675B",
    x"2CC51A4E",
    x"2CC4CD5F",
    x"2CC4808D",
    x"2CC433DA",
    x"2CC3E745",
    x"2CC39ACE",
    x"2CC34E74",
    x"2CC30238",
    x"2CC2B61A",
    x"2CC26A1A",
    x"2CC21E37",
    x"2CC1D272",
    x"2CC186CB",
    x"2CC13B41",
    x"2CC0EFD5",
    x"2CC0A486",
    x"2CC05954",
    x"2CC00E40",
    x"2CBFC349",
    x"2CBF786F",
    x"2CBF2DB3",
    x"2CBEE314",
    x"2CBE9891",
    x"2CBE4E2C",
    x"2CBE03E4",
    x"2CBDB9B9",
    x"2CBD6FAB",
    x"2CBD25BA",
    x"2CBCDBE6",
    x"2CBC922E",
    x"2CBC4893",
    x"2CBBFF16",
    x"2CBBB5B4",
    x"2CBB6C70",
    x"2CBB2347",
    x"2CBADA3C",
    x"2CBA914D",
    x"2CBA487A",
    x"2CB9FFC4",
    x"2CB9B72B",
    x"2CB96EAD",
    x"2CB9264C",
    x"2CB8DE07",
    x"2CB895DF",
    x"2CB84DD2",
    x"2CB805E2",
    x"2CB7BE0E",
    x"2CB77655",
    x"2CB72EB9",
    x"2CB6E739",
    x"2CB69FD4",
    x"2CB6588C",
    x"2CB6115F",
    x"2CB5CA4E",
    x"2CB58359",
    x"2CB53C80",
    x"2CB4F5C2",
    x"2CB4AF20",
    x"2CB46899",
    x"2CB4222E",
    x"2CB3DBDE",
    x"2CB395AA",
    x"2CB34F91",
    x"2CB30994",
    x"2CB2C3B2",
    x"2CB27DEB",
    x"2CB23840",
    x"2CB1F2AF",
    x"2CB1AD3A",
    x"2CB167E0",
    x"2CB122A1",
    x"2CB0DD7D",
    x"2CB09874",
    x"2CB05386",
    x"2CB00EB2",
    x"2CAFC9FA",
    x"2CAF855D",
    x"2CAF40DA",
    x"2CAEFC72",
    x"2CAEB825",
    x"2CAE73F2",
    x"2CAE2FDA",
    x"2CADEBDD",
    x"2CADA7FA",
    x"2CAD6431",
    x"2CAD2084",
    x"2CACDCF0",
    x"2CAC9977",
    x"2CAC5618",
    x"2CAC12D4",
    x"2CABCFA9",
    x"2CAB8C99",
    x"2CAB49A4",
    x"2CAB06C8",
    x"2CAAC406",
    x"2CAA815F",
    x"2CAA3ED1",
    x"2CA9FC5E",
    x"2CA9BA04",
    x"2CA977C4",
    x"2CA9359E",
    x"2CA8F392",
    x"2CA8B1A0",
    x"2CA86FC8",
    x"2CA82E09",
    x"2CA7EC64",
    x"2CA7AAD8",
    x"2CA76966",
    x"2CA7280E",
    x"2CA6E6CF",
    x"2CA6A5A9",
    x"2CA6649D",
    x"2CA623AB",
    x"2CA5E2D1",
    x"2CA5A212",
    x"2CA5616B",
    x"2CA520DD",
    x"2CA4E069",
    x"2CA4A00E",
    x"2CA45FCC",
    x"2CA41FA3",
    x"2CA3DF93",
    x"2CA39F9D",
    x"2CA35FBF",
    x"2CA31FFA",
    x"2CA2E04E",
    x"2CA2A0BA",
    x"2CA26140",
    x"2CA221DE",
    x"2CA1E296",
    x"2CA1A365",
    x"2CA1644E",
    x"2CA1254F",
    x"2CA0E669",
    x"2CA0A79B",
    x"2CA068E6",
    x"2CA02A49",
    x"2C9FEBC5",
    x"2C9FAD59",
    x"2C9F6F05",
    x"2C9F30CA",
    x"2C9EF2A7",
    x"2C9EB49D",
    x"2C9E76AA",
    x"2C9E38D0",
    x"2C9DFB0E",
    x"2C9DBD64",
    x"2C9D7FD2",
    x"2C9D4258",
    x"2C9D04F6",
    x"2C9CC7AC",
    x"2C9C8A7A",
    x"2C9C4D60",
    x"2C9C105D",
    x"2C9BD373",
    x"2C9B96A0",
    x"2C9B59E5",
    x"2C9B1D42",
    x"2C9AE0B6",
    x"2C9AA442",
    x"2C9A67E6",
    x"2C9A2BA1",
    x"2C99EF74",
    x"2C99B35E",
    x"2C997760",
    x"2C993B79",
    x"2C98FFA9",
    x"2C98C3F1",
    x"2C988850",
    x"2C984CC7",
    x"2C981154",
    x"2C97D5F9",
    x"2C979AB5",
    x"2C975F88",
    x"2C972472",
    x"2C96E974",
    x"2C96AE8C",
    x"2C9673BB",
    x"2C963902",
    x"2C95FE5F",
    x"2C95C3D3",
    x"2C95895E",
    x"2C954F00",
    x"2C9514B8",
    x"2C94DA87",
    x"2C94A06D",
    x"2C94666A",
    x"2C942C7D",
    x"2C93F2A7",
    x"2C93B8E8",
    x"2C937F3F",
    x"2C9345AC",
    x"2C930C30",
    x"2C92D2CB",
    x"2C92997C",
    x"2C926043",
    x"2C922720",
    x"2C91EE14",
    x"2C91B51E",
    x"2C917C3F",
    x"2C914375",
    x"2C910AC2",
    x"2C90D225",
    x"2C90999E",
    x"2C90612D",
    x"2C9028D2",
    x"2C8FF08D",
    x"2C8FB85E",
    x"2C8F8045",
    x"2C8F4842",
    x"2C8F1054",
    x"2C8ED87D",
    x"2C8EA0BB",
    x"2C8E690F",
    x"2C8E3179",
    x"2C8DF9F9",
    x"2C8DC28E",
    x"2C8D8B39",
    x"2C8D53F9",
    x"2C8D1CCF",
    x"2C8CE5BB",
    x"2C8CAEBC",
    x"2C8C77D2",
    x"2C8C40FE",
    x"2C8C0A3F",
    x"2C8BD396",
    x"2C8B9D02",
    x"2C8B6683",
    x"2C8B301A",
    x"2C8AF9C6",
    x"2C8AC387",
    x"2C8A8D5D",
    x"2C8A5748",
    x"2C8A2149",
    x"2C89EB5E",
    x"2C89B589",
    x"2C897FC8",
    x"2C894A1D",
    x"2C891487",
    x"2C88DF05",
    x"2C88A998",
    x"2C887440",
    x"2C883EFD",
    x"2C8809CF",
    x"2C87D4B6",
    x"2C879FB1",
    x"2C876AC1",
    x"2C8735E6",
    x"2C87011F",
    x"2C86CC6D",
    x"2C8697CF",
    x"2C866346",
    x"2C862ED2",
    x"2C85FA72",
    x"2C85C626",
    x"2C8591EF",
    x"2C855DCC",
    x"2C8529BD",
    x"2C84F5C3",
    x"2C84C1DD",
    x"2C848E0C",
    x"2C845A4E",
    x"2C8426A5",
    x"2C83F310",
    x"2C83BF8F",
    x"2C838C23",
    x"2C8358CA",
    x"2C832585",
    x"2C82F255",
    x"2C82BF38",
    x"2C828C2F",
    x"2C82593A",
    x"2C822659",
    x"2C81F38C",
    x"2C81C0D3",
    x"2C818E2E",
    x"2C815B9C",
    x"2C81291E",
    x"2C80F6B4",
    x"2C80C45D",
    x"2C80921B",
    x"2C805FEB",
    x"2C802DD0",
    x"2C7FF78F",
    x"2C7F93A6",
    x"2C7F2FE4",
    x"2C7ECC48",
    x"2C7E68D4",
    x"2C7E0586",
    x"2C7DA260",
    x"2C7D3F60",
    x"2C7CDC86",
    x"2C7C79D3",
    x"2C7C1747",
    x"2C7BB4E1",
    x"2C7B52A2",
    x"2C7AF088",
    x"2C7A8E96",
    x"2C7A2CC9",
    x"2C79CB23",
    x"2C7969A2",
    x"2C790848",
    x"2C78A714",
    x"2C784606",
    x"2C77E51D",
    x"2C77845A",
    x"2C7723BE",
    x"2C76C347",
    x"2C7662F5",
    x"2C7602C9",
    x"2C75A2C3",
    x"2C7542E2",
    x"2C74E327",
    x"2C748391",
    x"2C742420",
    x"2C73C4D4",
    x"2C7365AE",
    x"2C7306AD",
    x"2C72A7D1",
    x"2C72491A",
    x"2C71EA88",
    x"2C718C1A",
    x"2C712DD2",
    x"2C70CFAF",
    x"2C7071B0",
    x"2C7013D6",
    x"2C6FB620",
    x"2C6F5890",
    x"2C6EFB23",
    x"2C6E9DDB",
    x"2C6E40B8",
    x"2C6DE3B9",
    x"2C6D86DE",
    x"2C6D2A27",
    x"2C6CCD95",
    x"2C6C7127",
    x"2C6C14DD",
    x"2C6BB8B6",
    x"2C6B5CB4",
    x"2C6B00D6",
    x"2C6AA51C",
    x"2C6A4985",
    x"2C69EE12",
    x"2C6992C3",
    x"2C693797",
    x"2C68DC90",
    x"2C6881AB",
    x"2C6826EA",
    x"2C67CC4D",
    x"2C6771D3",
    x"2C67177C",
    x"2C66BD48",
    x"2C666338",
    x"2C66094B",
    x"2C65AF81",
    x"2C6555DA",
    x"2C64FC55",
    x"2C64A2F4",
    x"2C6449B6",
    x"2C63F09B",
    x"2C6397A2",
    x"2C633ECC",
    x"2C62E619",
    x"2C628D89",
    x"2C62351A",
    x"2C61DCCF",
    x"2C6184A6",
    x"2C612C9F",
    x"2C60D4BB",
    x"2C607CF9",
    x"2C602559",
    x"2C5FCDDC",
    x"2C5F7681",
    x"2C5F1F47",
    x"2C5EC830",
    x"2C5E713B",
    x"2C5E1A68",
    x"2C5DC3B6",
    x"2C5D6D27",
    x"2C5D16B9",
    x"2C5CC06D",
    x"2C5C6A43",
    x"2C5C143A",
    x"2C5BBE53",
    x"2C5B688D",
    x"2C5B12E9",
    x"2C5ABD66",
    x"2C5A6805",
    x"2C5A12C5",
    x"2C59BDA6",
    x"2C5968A9",
    x"2C5913CD",
    x"2C58BF11",
    x"2C586A77",
    x"2C5815FE",
    x"2C57C1A6",
    x"2C576D6F",
    x"2C571959",
    x"2C56C563",
    x"2C56718E",
    x"2C561DDA",
    x"2C55CA47",
    x"2C5576D4",
    x"2C552382",
    x"2C54D051",
    x"2C547D3F",
    x"2C542A4F",
    x"2C53D77E",
    x"2C5384CE",
    x"2C53323F",
    x"2C52DFCF",
    x"2C528D80",
    x"2C523B51",
    x"2C51E941",
    x"2C519752",
    x"2C514583",
    x"2C50F3D4",
    x"2C50A245",
    x"2C5050D5",
    x"2C4FFF86",
    x"2C4FAE56",
    x"2C4F5D45",
    x"2C4F0C55",
    x"2C4EBB84",
    x"2C4E6AD2",
    x"2C4E1A40",
    x"2C4DC9CE",
    x"2C4D797B",
    x"2C4D2947",
    x"2C4CD932",
    x"2C4C893D",
    x"2C4C3967",
    x"2C4BE9B0",
    x"2C4B9A18",
    x"2C4B4AA0",
    x"2C4AFB46",
    x"2C4AAC0B",
    x"2C4A5CF0",
    x"2C4A0DF3",
    x"2C49BF15",
    x"2C497056",
    x"2C4921B5",
    x"2C48D333",
    x"2C4884D0",
    x"2C48368B",
    x"2C47E865",
    x"2C479A5E",
    x"2C474C75",
    x"2C46FEAA",
    x"2C46B0FE",
    x"2C466370",
    x"2C461600",
    x"2C45C8AF",
    x"2C457B7B",
    x"2C452E66",
    x"2C44E16F",
    x"2C449496",
    x"2C4447DB",
    x"2C43FB3E",
    x"2C43AEBF",
    x"2C43625D",
    x"2C43161A",
    x"2C42C9F4",
    x"2C427DEC",
    x"2C423202",
    x"2C41E635",
    x"2C419A86",
    x"2C414EF4",
    x"2C410380",
    x"2C40B829",
    x"2C406CF0",
    x"2C4021D4",
    x"2C3FD6D6",
    x"2C3F8BF4",
    x"2C3F4130",
    x"2C3EF689",
    x"2C3EAC00",
    x"2C3E6193",
    x"2C3E1743",
    x"2C3DCD11",
    x"2C3D82FB",
    x"2C3D3903",
    x"2C3CEF27",
    x"2C3CA568",
    x"2C3C5BC5",
    x"2C3C1240",
    x"2C3BC8D7",
    x"2C3B7F8B",
    x"2C3B365C",
    x"2C3AED49",
    x"2C3AA452",
    x"2C3A5B78",
    x"2C3A12BB",
    x"2C39CA1A",
    x"2C398195",
    x"2C39392C",
    x"2C38F0E0",
    x"2C38A8B0",
    x"2C38609C",
    x"2C3818A5",
    x"2C37D0C9",
    x"2C378909",
    x"2C374166",
    x"2C36F9DE",
    x"2C36B273",
    x"2C366B23",
    x"2C3623EF",
    x"2C35DCD7",
    x"2C3595DA",
    x"2C354EFA",
    x"2C350835",
    x"2C34C18B",
    x"2C347AFE",
    x"2C34348B",
    x"2C33EE34",
    x"2C33A7F9",
    x"2C3361D9",
    x"2C331BD5",
    x"2C32D5EB",
    x"2C32901E",
    x"2C324A6B",
    x"2C3204D3",
    x"2C31BF57",
    x"2C3179F6",
    x"2C3134B0",
    x"2C30EF85",
    x"2C30AA75",
    x"2C306580",
    x"2C3020A5",
    x"2C2FDBE6",
    x"2C2F9742",
    x"2C2F52B8",
    x"2C2F0E49",
    x"2C2EC9F5",
    x"2C2E85BB",
    x"2C2E419C",
    x"2C2DFD98",
    x"2C2DB9AE",
    x"2C2D75DF",
    x"2C2D322A",
    x"2C2CEE90",
    x"2C2CAB10",
    x"2C2C67AA",
    x"2C2C245F",
    x"2C2BE12D",
    x"2C2B9E17",
    x"2C2B5B1A",
    x"2C2B1837",
    x"2C2AD56F",
    x"2C2A92C1",
    x"2C2A502C",
    x"2C2A0DB2",
    x"2C29CB52",
    x"2C29890B",
    x"2C2946DF",
    x"2C2904CC",
    x"2C28C2D3",
    x"2C2880F4",
    x"2C283F2E",
    x"2C27FD82",
    x"2C27BBF0",
    x"2C277A77",
    x"2C273918",
    x"2C26F7D3",
    x"2C26B6A7",
    x"2C267594",
    x"2C26349B",
    x"2C25F3BB",
    x"2C25B2F4",
    x"2C257247",
    x"2C2531B3",
    x"2C24F138",
    x"2C24B0D7",
    x"2C24708E",
    x"2C24305F",
    x"2C23F048",
    x"2C23B04B",
    x"2C237067",
    x"2C23309B",
    x"2C22F0E9",
    x"2C22B14F",
    x"2C2271CE",
    x"2C223266",
    x"2C21F317",
    x"2C21B3E0",
    x"2C2174C2",
    x"2C2135BD",
    x"2C20F6D0",
    x"2C20B7FC",
    x"2C207940",
    x"2C203A9D",
    x"2C1FFC13",
    x"2C1FBDA0",
    x"2C1F7F46",
    x"2C1F4105",
    x"2C1F02DC",
    x"2C1EC4CB",
    x"2C1E86D2",
    x"2C1E48F1",
    x"2C1E0B29",
    x"2C1DCD79",
    x"2C1D8FE0",
    x"2C1D5260",
    x"2C1D14F8",
    x"2C1CD7A8",
    x"2C1C9A6F",
    x"2C1C5D4F",
    x"2C1C2047",
    x"2C1BE356",
    x"2C1BA67D",
    x"2C1B69BC",
    x"2C1B2D12",
    x"2C1AF081",
    x"2C1AB406",
    x"2C1A77A4",
    x"2C1A3B59",
    x"2C19FF25",
    x"2C19C30A",
    x"2C198705",
    x"2C194B18",
    x"2C190F42",
    x"2C18D384",
    x"2C1897DD",
    x"2C185C4D",
    x"2C1820D5",
    x"2C17E574",
    x"2C17AA2A",
    x"2C176EF7",
    x"2C1733DB",
    x"2C16F8D6",
    x"2C16BDE9",
    x"2C168312",
    x"2C164852",
    x"2C160DA9",
    x"2C15D318",
    x"2C15989D",
    x"2C155E38",
    x"2C1523EB",
    x"2C14E9B4",
    x"2C14AF94",
    x"2C14758B",
    x"2C143B98",
    x"2C1401BC",
    x"2C13C7F7",
    x"2C138E48",
    x"2C1354B0",
    x"2C131B2E",
    x"2C12E1C3",
    x"2C12A86E",
    x"2C126F2F",
    x"2C123607",
    x"2C11FCF5",
    x"2C11C3F9",
    x"2C118B14",
    x"2C115245",
    x"2C11198B",
    x"2C10E0E9",
    x"2C10A85C",
    x"2C106FE5",
    x"2C103784",
    x"2C0FFF3A",
    x"2C0FC705",
    x"2C0F8EE6",
    x"2C0F56DD",
    x"2C0F1EEA",
    x"2C0EE70D",
    x"2C0EAF46",
    x"2C0E7794",
    x"2C0E3FF8",
    x"2C0E0872",
    x"2C0DD102",
    x"2C0D99A7",
    x"2C0D6262",
    x"2C0D2B32",
    x"2C0CF418",
    x"2C0CBD13",
    x"2C0C8624",
    x"2C0C4F4A",
    x"2C0C1886",
    x"2C0BE1D7",
    x"2C0BAB3E",
    x"2C0B74BA",
    x"2C0B3E4B",
    x"2C0B07F1",
    x"2C0AD1AC",
    x"2C0A9B7D",
    x"2C0A6563",
    x"2C0A2F5E",
    x"2C09F96E",
    x"2C09C393",
    x"2C098DCD",
    x"2C09581C",
    x"2C092280",
    x"2C08ECF9",
    x"2C08B787",
    x"2C08822A",
    x"2C084CE1",
    x"2C0817AE",
    x"2C07E28F",
    x"2C07AD85",
    x"2C07788F",
    x"2C0743AE",
    x"2C070EE2",
    x"2C06DA2B",
    x"2C06A588",
    x"2C0670FA",
    x"2C063C80",
    x"2C06081A",
    x"2C05D3C9",
    x"2C059F8D",
    x"2C056B65",
    x"2C053751",
    x"2C050351",
    x"2C04CF66",
    x"2C049B8F",
    x"2C0467CD",
    x"2C04341E",
    x"2C040084",
    x"2C03CCFE",
    x"2C03998C",
    x"2C03662E",
    x"2C0332E4",
    x"2C02FFAE",
    x"2C02CC8C",
    x"2C02997E",
    x"2C026684",
    x"2C02339E",
    x"2C0200CC",
    x"2C01CE0E",
    x"2C019B63",
    x"2C0168CC",
    x"2C013649",
    x"2C0103DA",
    x"2C00D17E",
    x"2C009F36",
    x"2C006D02",
    x"2C003AE1",
    x"2C0008D4",
    x"2BFFADB4",
    x"2BFF49E8",
    x"2BFEE642",
    x"2BFE82C4",
    x"2BFE1F6C",
    x"2BFDBC3B",
    x"2BFD5931",
    x"2BFCF64D",
    x"2BFC9391",
    x"2BFC30FA",
    x"2BFBCE8A",
    x"2BFB6C41",
    x"2BFB0A1E",
    x"2BFAA821",
    x"2BFA464A",
    x"2BF9E49A",
    x"2BF98310",
    x"2BF921AC",
    x"2BF8C06D",
    x"2BF85F55",
    x"2BF7FE63",
    x"2BF79D96",
    x"2BF73CF0",
    x"2BF6DC6F",
    x"2BF67C13",
    x"2BF61BDE",
    x"2BF5BBCE",
    x"2BF55BE3",
    x"2BF4FC1E",
    x"2BF49C7E",
    x"2BF43D04",
    x"2BF3DDAE",
    x"2BF37E7E",
    x"2BF31F74",
    x"2BF2C08E",
    x"2BF261CD",
    x"2BF20331",
    x"2BF1A4BB",
    x"2BF14669",
    x"2BF0E83C",
    x"2BF08A33",
    x"2BF02C50",
    x"2BEFCE91",
    x"2BEF70F6",
    x"2BEF1380",
    x"2BEEB62F",
    x"2BEE5902",
    x"2BEDFBF9",
    x"2BED9F15",
    x"2BED4255",
    x"2BECE5B9",
    x"2BEC8942",
    x"2BEC2CEE",
    x"2BEBD0BE",
    x"2BEB74B3",
    x"2BEB18CB",
    x"2BEABD08",
    x"2BEA6168",
    x"2BEA05EB",
    x"2BE9AA93",
    x"2BE94F5E",
    x"2BE8F44D",
    x"2BE8995F",
    x"2BE83E95",
    x"2BE7E3EE",
    x"2BE7896B",
    x"2BE72F0B",
    x"2BE6D4CE",
    x"2BE67AB5",
    x"2BE620BE",
    x"2BE5C6EB",
    x"2BE56D3B",
    x"2BE513AE",
    x"2BE4BA44",
    x"2BE460FC",
    x"2BE407D8",
    x"2BE3AED6",
    x"2BE355F7",
    x"2BE2FD3B",
    x"2BE2A4A1",
    x"2BE24C2A",
    x"2BE1F3D6",
    x"2BE19BA4",
    x"2BE14394",
    x"2BE0EBA7",
    x"2BE093DC",
    x"2BE03C33",
    x"2BDFE4AD",
    x"2BDF8D49",
    x"2BDF3607",
    x"2BDEDEE6",
    x"2BDE87E8",
    x"2BDE310C",
    x"2BDDDA52",
    x"2BDD83BA",
    x"2BDD2D43",
    x"2BDCD6EE",
    x"2BDC80BB",
    x"2BDC2AAA",
    x"2BDBD4BA",
    x"2BDB7EEC",
    x"2BDB293F",
    x"2BDAD3B3",
    x"2BDA7E49",
    x"2BDA2901",
    x"2BD9D3D9",
    x"2BD97ED3",
    x"2BD929EE",
    x"2BD8D52A",
    x"2BD88088",
    x"2BD82C06",
    x"2BD7D7A5",
    x"2BD78365",
    x"2BD72F47",
    x"2BD6DB48",
    x"2BD6876B",
    x"2BD633AF",
    x"2BD5E013",
    x"2BD58C98",
    x"2BD5393D",
    x"2BD4E603",
    x"2BD492E9",
    x"2BD43FF0",
    x"2BD3ED17",
    x"2BD39A5F",
    x"2BD347C7",
    x"2BD2F54F",
    x"2BD2A2F7",
    x"2BD250BF",
    x"2BD1FEA8",
    x"2BD1ACB0",
    x"2BD15AD9",
    x"2BD10921",
    x"2BD0B78A",
    x"2BD06612",
    x"2BD014BA",
    x"2BCFC382",
    x"2BCF7269",
    x"2BCF2170",
    x"2BCED097",
    x"2BCE7FDD",
    x"2BCE2F43",
    x"2BCDDEC8",
    x"2BCD8E6D",
    x"2BCD3E31",
    x"2BCCEE15",
    x"2BCC9E17",
    x"2BCC4E39",
    x"2BCBFE7A",
    x"2BCBAEDA",
    x"2BCB5F59",
    x"2BCB0FF8",
    x"2BCAC0B5",
    x"2BCA7191",
    x"2BCA228C",
    x"2BC9D3A6",
    x"2BC984DF",
    x"2BC93636",
    x"2BC8E7AC",
    x"2BC89941",
    x"2BC84AF5",
    x"2BC7FCC7",
    x"2BC7AEB7",
    x"2BC760C6",
    x"2BC712F4",
    x"2BC6C53F",
    x"2BC677A9",
    x"2BC62A32",
    x"2BC5DCD9",
    x"2BC58F9D",
    x"2BC54280",
    x"2BC4F581",
    x"2BC4A8A0",
    x"2BC45BDE",
    x"2BC40F39",
    x"2BC3C2B2",
    x"2BC37649",
    x"2BC329FD",
    x"2BC2DDD0",
    x"2BC291C0",
    x"2BC245CE",
    x"2BC1F9F9",
    x"2BC1AE43",
    x"2BC162A9",
    x"2BC1172D",
    x"2BC0CBCF",
    x"2BC0808E",
    x"2BC0356B",
    x"2BBFEA64",
    x"2BBF9F7C",
    x"2BBF54B0",
    x"2BBF0A01",
    x"2BBEBF70",
    x"2BBE74FC",
    x"2BBE2AA5",
    x"2BBDE06A",
    x"2BBD964D",
    x"2BBD4C4D",
    x"2BBD026A",
    x"2BBCB8A3",
    x"2BBC6EF9",
    x"2BBC256C",
    x"2BBBDBFC",
    x"2BBB92A9",
    x"2BBB4972",
    x"2BBB0057",
    x"2BBAB759",
    x"2BBA6E78",
    x"2BBA25B3",
    x"2BB9DD0A",
    x"2BB9947E",
    x"2BB94C0E",
    x"2BB903BB",
    x"2BB8BB83",
    x"2BB87368",
    x"2BB82B69",
    x"2BB7E386",
    x"2BB79BC0",
    x"2BB75415",
    x"2BB70C86",
    x"2BB6C513",
    x"2BB67DBC",
    x"2BB63681",
    x"2BB5EF61",
    x"2BB5A85E",
    x"2BB56176",
    x"2BB51AA9",
    x"2BB4D3F9",
    x"2BB48D64",
    x"2BB446EA",
    x"2BB4008C",
    x"2BB3BA4A",
    x"2BB37423",
    x"2BB32E17",
    x"2BB2E827",
    x"2BB2A252",
    x"2BB25C98",
    x"2BB216F9",
    x"2BB1D176",
    x"2BB18C0E",
    x"2BB146C1",
    x"2BB1018F",
    x"2BB0BC77",
    x"2BB0777B",
    x"2BB0329A",
    x"2BAFEDD4",
    x"2BAFA928",
    x"2BAF6498",
    x"2BAF2022",
    x"2BAEDBC6",
    x"2BAE9786",
    x"2BAE5360",
    x"2BAE0F55",
    x"2BADCB64",
    x"2BAD878E",
    x"2BAD43D2",
    x"2BAD0031",
    x"2BACBCAA",
    x"2BAC793D",
    x"2BAC35EB",
    x"2BABF2B3",
    x"2BABAF96",
    x"2BAB6C92",
    x"2BAB29A9",
    x"2BAAE6DA",
    x"2BAAA424",
    x"2BAA6189",
    x"2BAA1F08",
    x"2BA9DCA1",
    x"2BA99A54",
    x"2BA95820",
    x"2BA91607",
    x"2BA8D407",
    x"2BA89221",
    x"2BA85055",
    x"2BA80EA3",
    x"2BA7CD0A",
    x"2BA78B8A",
    x"2BA74A25",
    x"2BA708D8",
    x"2BA6C7A6",
    x"2BA6868C",
    x"2BA6458D",
    x"2BA604A6",
    x"2BA5C3D9",
    x"2BA58325",
    x"2BA5428A",
    x"2BA50209",
    x"2BA4C1A1",
    x"2BA48152",
    x"2BA4411C",
    x"2BA400FF",
    x"2BA3C0FB",
    x"2BA38110",
    x"2BA3413E",
    x"2BA30185",
    x"2BA2C1E5",
    x"2BA2825E",
    x"2BA242EF",
    x"2BA20399",
    x"2BA1C45C",
    x"2BA18538",
    x"2BA1462C",
    x"2BA10739",
    x"2BA0C85F",
    x"2BA0899D",
    x"2BA04AF3",
    x"2BA00C62",
    x"2B9FCDE9",
    x"2B9F8F89",
    x"2B9F5141",
    x"2B9F1312",
    x"2B9ED4FA",
    x"2B9E96FB",
    x"2B9E5914",
    x"2B9E1B46",
    x"2B9DDD8F",
    x"2B9D9FF0",
    x"2B9D626A",
    x"2B9D24FC",
    x"2B9CE7A5",
    x"2B9CAA67",
    x"2B9C6D40",
    x"2B9C3031",
    x"2B9BF33A",
    x"2B9BB65B",
    x"2B9B7994",
    x"2B9B3CE4",
    x"2B9B004C",
    x"2B9AC3CC",
    x"2B9A8763",
    x"2B9A4B12",
    x"2B9A0ED9",
    x"2B99D2B7",
    x"2B9996AC",
    x"2B995AB9",
    x"2B991EDD",
    x"2B98E319",
    x"2B98A76C",
    x"2B986BD6",
    x"2B983057",
    x"2B97F4F0",
    x"2B97B9A0",
    x"2B977E67",
    x"2B974345",
    x"2B97083B",
    x"2B96CD47",
    x"2B96926A",
    x"2B9657A4",
    x"2B961CF6",
    x"2B95E25E",
    x"2B95A7DD",
    x"2B956D73",
    x"2B95331F",
    x"2B94F8E3",
    x"2B94BEBD",
    x"2B9484AE",
    x"2B944AB5",
    x"2B9410D3",
    x"2B93D708",
    x"2B939D53",
    x"2B9363B5",
    x"2B932A2D",
    x"2B92F0BC",
    x"2B92B761",
    x"2B927E1D",
    x"2B9244EF",
    x"2B920BD7",
    x"2B91D2D5",
    x"2B9199EA",
    x"2B916115",
    x"2B912856",
    x"2B90EFAE",
    x"2B90B71B",
    x"2B907E9F",
    x"2B904638",
    x"2B900DE8",
    x"2B8FD5AD",
    x"2B8F9D89",
    x"2B8F657A",
    x"2B8F2D82",
    x"2B8EF59F",
    x"2B8EBDD2",
    x"2B8E861A",
    x"2B8E4E79",
    x"2B8E16ED",
    x"2B8DDF77",
    x"2B8DA816",
    x"2B8D70CC",
    x"2B8D3996",
    x"2B8D0277",
    x"2B8CCB6C",
    x"2B8C9478",
    x"2B8C5D98",
    x"2B8C26CF",
    x"2B8BF01A",
    x"2B8BB97B",
    x"2B8B82F1",
    x"2B8B4C7D",
    x"2B8B161D",
    x"2B8ADFD3",
    x"2B8AA99F",
    x"2B8A737F",
    x"2B8A3D74",
    x"2B8A077F",
    x"2B89D19E",
    x"2B899BD3",
    x"2B89661D",
    x"2B89307B",
    x"2B88FAEF",
    x"2B88C577",
    x"2B889014",
    x"2B885AC7",
    x"2B88258E",
    x"2B87F069",
    x"2B87BB5A",
    x"2B87865F",
    x"2B875179",
    x"2B871CA7",
    x"2B86E7EA",
    x"2B86B342",
    x"2B867EAE",
    x"2B864A2F",
    x"2B8615C4",
    x"2B85E16E",
    x"2B85AD2C",
    x"2B8578FF",
    x"2B8544E6",
    x"2B8510E1",
    x"2B84DCF0",
    x"2B84A914",
    x"2B84754C",
    x"2B844199",
    x"2B840DF9",
    x"2B83DA6E",
    x"2B83A6F6",
    x"2B837393",
    x"2B834044",
    x"2B830D09",
    x"2B82D9E2",
    x"2B82A6CF",
    x"2B8273D0",
    x"2B8240E4",
    x"2B820E0D",
    x"2B81DB49",
    x"2B81A89A",
    x"2B8175FE",
    x"2B814375",
    x"2B811101",
    x"2B80DEA0",
    x"2B80AC53",
    x"2B807A19",
    x"2B8047F4",
    x"2B8015E1",
    x"2B7FC7C5",
    x"2B7F63EE",
    x"2B7F003F",
    x"2B7E9CB6",
    x"2B7E3954",
    x"2B7DD619",
    x"2B7D7305",
    x"2B7D1017",
    x"2B7CAD50",
    x"2B7C4AB0",
    x"2B7BE836",
    x"2B7B85E3",
    x"2B7B23B5",
    x"2B7AC1AF",
    x"2B7A5FCE",
    x"2B79FE14",
    x"2B799C80",
    x"2B793B12",
    x"2B78D9C9",
    x"2B7878A7",
    x"2B7817AB",
    x"2B77B6D5",
    x"2B775624",
    x"2B76F59A",
    x"2B769534",
    x"2B7634F5",
    x"2B75D4DB",
    x"2B7574E7",
    x"2B751518",
    x"2B74B56E",
    x"2B7455EA",
    x"2B73F68B",
    x"2B739751",
    x"2B73383D",
    x"2B72D94D",
    x"2B727A83",
    x"2B721BDE",
    x"2B71BD5D",
    x"2B715F02",
    x"2B7100CB",
    x"2B70A2B9",
    x"2B7044CC",
    x"2B6FE703",
    x"2B6F895F",
    x"2B6F2BE0",
    x"2B6ECE85",
    x"2B6E714F",
    x"2B6E143C",
    x"2B6DB74F",
    x"2B6D5A85",
    x"2B6CFDE0",
    x"2B6CA15F",
    x"2B6C4502",
    x"2B6BE8C9",
    x"2B6B8CB4",
    x"2B6B30C3",
    x"2B6AD4F6",
    x"2B6A794D",
    x"2B6A1DC7",
    x"2B69C265",
    x"2B696727",
    x"2B690C0D",
    x"2B68B116",
    x"2B685642",
    x"2B67FB92",
    x"2B67A106",
    x"2B67469D",
    x"2B66EC57",
    x"2B669234",
    x"2B663834",
    x"2B65DE58",
    x"2B65849F",
    x"2B652B08",
    x"2B64D195",
    x"2B647845",
    x"2B641F17",
    x"2B63C60C",
    x"2B636D24",
    x"2B63145F",
    x"2B62BBBC",
    x"2B62633C",
    x"2B620ADF",
    x"2B61B2A4",
    x"2B615A8B",
    x"2B610295",
    x"2B60AAC1",
    x"2B605310",
    x"2B5FFB80",
    x"2B5FA413",
    x"2B5F4CC8",
    x"2B5EF59F",
    x"2B5E9E98",
    x"2B5E47B3",
    x"2B5DF0F0",
    x"2B5D9A4F",
    x"2B5D43D0",
    x"2B5CED72",
    x"2B5C9736",
    x"2B5C411C",
    x"2B5BEB23",
    x"2B5B954C",
    x"2B5B3F97",
    x"2B5AEA02",
    x"2B5A9490",
    x"2B5A3F3E",
    x"2B59EA0E",
    x"2B5994FF",
    x"2B594012",
    x"2B58EB45",
    x"2B58969A",
    x"2B584210",
    x"2B57EDA6",
    x"2B57995E",
    x"2B574537",
    x"2B56F130",
    x"2B569D4A",
    x"2B564985",
    x"2B55F5E1",
    x"2B55A25D",
    x"2B554EFA",
    x"2B54FBB7",
    x"2B54A895",
    x"2B545594",
    x"2B5402B2",
    x"2B53AFF1",
    x"2B535D51",
    x"2B530AD0",
    x"2B52B870",
    x"2B526630",
    x"2B521410",
    x"2B51C211",
    x"2B517031",
    x"2B511E71",
    x"2B50CCD1",
    x"2B507B51",
    x"2B5029F1",
    x"2B4FD8B0",
    x"2B4F878F",
    x"2B4F368E",
    x"2B4EE5AD",
    x"2B4E94EB",
    x"2B4E4448",
    x"2B4DF3C5",
    x"2B4DA362",
    x"2B4D531E",
    x"2B4D02F9",
    x"2B4CB2F3",
    x"2B4C630D",
    x"2B4C1346",
    x"2B4BC39E",
    x"2B4B7415",
    x"2B4B24AB",
    x"2B4AD561",
    x"2B4A8635",
    x"2B4A3728",
    x"2B49E83A",
    x"2B49996A",
    x"2B494ABA",
    x"2B48FC28",
    x"2B48ADB5",
    x"2B485F60",
    x"2B48112A",
    x"2B47C313",
    x"2B47751A",
    x"2B47273F",
    x"2B46D983",
    x"2B468BE5",
    x"2B463E66",
    x"2B45F104",
    x"2B45A3C1",
    x"2B45569D",
    x"2B450996",
    x"2B44BCAD",
    x"2B446FE2",
    x"2B442336",
    x"2B43D6A7",
    x"2B438A36",
    x"2B433DE3",
    x"2B42F1AE",
    x"2B42A596",
    x"2B42599C",
    x"2B420DC0",
    x"2B41C201",
    x"2B417660",
    x"2B412ADD",
    x"2B40DF77",
    x"2B40942E",
    x"2B404903",
    x"2B3FFDF5",
    x"2B3FB305",
    x"2B3F6831",
    x"2B3F1D7B",
    x"2B3ED2E2",
    x"2B3E8867",
    x"2B3E3E08",
    x"2B3DF3C6",
    x"2B3DA9A1",
    x"2B3D5F99",
    x"2B3D15AF",
    x"2B3CCBE1",
    x"2B3C822F",
    x"2B3C389B",
    x"2B3BEF23",
    x"2B3BA5C8",
    x"2B3B5C8A",
    x"2B3B1368",
    x"2B3ACA62",
    x"2B3A817A",
    x"2B3A38AD",
    x"2B39EFFD",
    x"2B39A76A",
    x"2B395EF2",
    x"2B391697",
    x"2B38CE59",
    x"2B388636",
    x"2B383E30",
    x"2B37F646",
    x"2B37AE77",
    x"2B3766C5",
    x"2B371F2F",
    x"2B36D7B5",
    x"2B369057",
    x"2B364914",
    x"2B3601EE",
    x"2B35BAE3",
    x"2B3573F4",
    x"2B352D20",
    x"2B34E668",
    x"2B349FCC",
    x"2B34594B",
    x"2B3412E6",
    x"2B33CC9D",
    x"2B33866E",
    x"2B33405C",
    x"2B32FA64",
    x"2B32B488",
    x"2B326EC7",
    x"2B322921",
    x"2B31E397",
    x"2B319E28",
    x"2B3158D3",
    x"2B31139A",
    x"2B30CE7C",
    x"2B308979",
    x"2B304491",
    x"2B2FFFC3",
    x"2B2FBB11",
    x"2B2F7679",
    x"2B2F31FC",
    x"2B2EED9A",
    x"2B2EA953",
    x"2B2E6526",
    x"2B2E2114",
    x"2B2DDD1C",
    x"2B2D993F",
    x"2B2D557C",
    x"2B2D11D4",
    x"2B2CCE46",
    x"2B2C8AD3",
    x"2B2C477A",
    x"2B2C043B",
    x"2B2BC116",
    x"2B2B7E0C",
    x"2B2B3B1C",
    x"2B2AF846",
    x"2B2AB58A",
    x"2B2A72E8",
    x"2B2A3060",
    x"2B29EDF2",
    x"2B29AB9E",
    x"2B296964",
    x"2B292744",
    x"2B28E53D",
    x"2B28A351",
    x"2B28617E",
    x"2B281FC5",
    x"2B27DE25",
    x"2B279C9F",
    x"2B275B33",
    x"2B2719E0",
    x"2B26D8A6",
    x"2B269787",
    x"2B265680",
    x"2B261593",
    x"2B25D4BF",
    x"2B259405",
    x"2B255364",
    x"2B2512DC",
    x"2B24D26D",
    x"2B249217",
    x"2B2451DB",
    x"2B2411B7",
    x"2B23D1AD",
    x"2B2391BB",
    x"2B2351E3",
    x"2B231223",
    x"2B22D27D",
    x"2B2292EF",
    x"2B22537A",
    x"2B22141E",
    x"2B21D4DA",
    x"2B2195AF",
    x"2B21569D",
    x"2B2117A4",
    x"2B20D8C3",
    x"2B2099FA",
    x"2B205B4A",
    x"2B201CB3",
    x"2B1FDE34",
    x"2B1F9FCD",
    x"2B1F617F",
    x"2B1F2349",
    x"2B1EE52C",
    x"2B1EA726",
    x"2B1E6939",
    x"2B1E2B64",
    x"2B1DEDA7",
    x"2B1DB002",
    x"2B1D7276",
    x"2B1D3501",
    x"2B1CF7A4",
    x"2B1CBA5F",
    x"2B1C7D33",
    x"2B1C401E",
    x"2B1C0320",
    x"2B1BC63B",
    x"2B1B896E",
    x"2B1B4CB8",
    x"2B1B101A",
    x"2B1AD393",
    x"2B1A9724",
    x"2B1A5ACD",
    x"2B1A1E8D",
    x"2B19E265",
    x"2B19A654",
    x"2B196A5B",
    x"2B192E79",
    x"2B18F2AF",
    x"2B18B6FC",
    x"2B187B60",
    x"2B183FDB",
    x"2B18046E",
    x"2B17C918",
    x"2B178DD9",
    x"2B1752B1",
    x"2B1717A0",
    x"2B16DCA7",
    x"2B16A1C4",
    x"2B1666F8",
    x"2B162C43",
    x"2B15F1A6",
    x"2B15B71F",
    x"2B157CAF",
    x"2B154255",
    x"2B150813",
    x"2B14CDE7",
    x"2B1493D2",
    x"2B1459D3",
    x"2B141FEC",
    x"2B13E61A",
    x"2B13AC60",
    x"2B1372BC",
    x"2B13392E",
    x"2B12FFB7",
    x"2B12C656",
    x"2B128D0C",
    x"2B1253D8",
    x"2B121ABB",
    x"2B11E1B3",
    x"2B11A8C2",
    x"2B116FE7",
    x"2B113723",
    x"2B10FE74",
    x"2B10C5DC",
    x"2B108D5A",
    x"2B1054EE",
    x"2B101C97",
    x"2B0FE457",
    x"2B0FAC2D",
    x"2B0F7419",
    x"2B0F3C1A",
    x"2B0F0432",
    x"2B0ECC5F",
    x"2B0E94A2",
    x"2B0E5CFB",
    x"2B0E2569",
    x"2B0DEDEE",
    x"2B0DB688",
    x"2B0D7F37",
    x"2B0D47FC",
    x"2B0D10D7",
    x"2B0CD9C7",
    x"2B0CA2CD",
    x"2B0C6BE8",
    x"2B0C3518",
    x"2B0BFE5E",
    x"2B0BC7BA",
    x"2B0B912A",
    x"2B0B5AB0",
    x"2B0B244B",
    x"2B0AEDFC",
    x"2B0AB7C1",
    x"2B0A819C",
    x"2B0A4B8C",
    x"2B0A1591",
    x"2B09DFAB",
    x"2B09A9DA",
    x"2B09741F",
    x"2B093E78",
    x"2B0908E6",
    x"2B08D369",
    x"2B089E01",
    x"2B0868AD",
    x"2B08336F",
    x"2B07FE45",
    x"2B07C930",
    x"2B079430",
    x"2B075F44",
    x"2B072A6D",
    x"2B06F5AB",
    x"2B06C0FE",
    x"2B068C64",
    x"2B0657E0",
    x"2B062370",
    x"2B05EF14",
    x"2B05BACD",
    x"2B05869A",
    x"2B05527C",
    x"2B051E72",
    x"2B04EA7C",
    x"2B04B69B",
    x"2B0482CD",
    x"2B044F14",
    x"2B041B70",
    x"2B03E7DF",
    x"2B03B462",
    x"2B0380FA",
    x"2B034DA6",
    x"2B031A65",
    x"2B02E739",
    x"2B02B421",
    x"2B02811C",
    x"2B024E2C",
    x"2B021B4F",
    x"2B01E886",
    x"2B01B5D2",
    x"2B018330",
    x"2B0150A3",
    x"2B011E29",
    x"2B00EBC3",
    x"2B00B971",
    x"2B008733",
    x"2B005508",
    x"2B0022F0",
    x"2AFFE1D8",
    x"2AFF7DF8",
    x"2AFF1A3E",
    x"2AFEB6AB",
    x"2AFE533F",
    x"2AFDEFFA",
    x"2AFD8CDC",
    x"2AFD29E4",
    x"2AFCC713",
    x"2AFC6469",
    x"2AFC01E5",
    x"2AFB9F87",
    x"2AFB3D50",
    x"2AFADB3F",
    x"2AFA7955",
    x"2AFA1790",
    x"2AF9B5F2",
    x"2AF9547A",
    x"2AF8F328",
    x"2AF891FC",
    x"2AF830F6",
    x"2AF7D016",
    x"2AF76F5C",
    x"2AF70EC7",
    x"2AF6AE58",
    x"2AF64E0F",
    x"2AF5EDEB",
    x"2AF58DED",
    x"2AF52E14",
    x"2AF4CE61",
    x"2AF46ED3",
    x"2AF40F6A",
    x"2AF3B027",
    x"2AF35109",
    x"2AF2F20F",
    x"2AF2933B",
    x"2AF2348C",
    x"2AF1D602",
    x"2AF1779D",
    x"2AF1195D",
    x"2AF0BB41",
    x"2AF05D4B",
    x"2AEFFF78",
    x"2AEFA1CB",
    x"2AEF4442",
    x"2AEEE6DE",
    x"2AEE899E",
    x"2AEE2C82",
    x"2AEDCF8B",
    x"2AED72B8",
    x"2AED1609",
    x"2AECB97F",
    x"2AEC5D18",
    x"2AEC00D6",
    x"2AEBA4B8",
    x"2AEB48BD",
    x"2AEAECE7",
    x"2AEA9134",
    x"2AEA35A5",
    x"2AE9DA3A",
    x"2AE97EF3",
    x"2AE923CF",
    x"2AE8C8CF",
    x"2AE86DF2",
    x"2AE81339",
    x"2AE7B8A3",
    x"2AE75E31",
    x"2AE703E1",
    x"2AE6A9B6",
    x"2AE64FAD",
    x"2AE5F5C7",
    x"2AE59C05",
    x"2AE54265",
    x"2AE4E8E9",
    x"2AE48F8F",
    x"2AE43659",
    x"2AE3DD45",
    x"2AE38454",
    x"2AE32B86",
    x"2AE2D2DA",
    x"2AE27A51",
    x"2AE221EA",
    x"2AE1C9A6",
    x"2AE17185",
    x"2AE11986",
    x"2AE0C1A9",
    x"2AE069EE",
    x"2AE01256",
    x"2ADFBAE0",
    x"2ADF638C",
    x"2ADF0C5A",
    x"2ADEB54A",
    x"2ADE5E5C",
    x"2ADE0791",
    x"2ADDB0E7",
    x"2ADD5A5E",
    x"2ADD03F8",
    x"2ADCADB3",
    x"2ADC5790",
    x"2ADC018F",
    x"2ADBABAF",
    x"2ADB55F1",
    x"2ADB0054",
    x"2ADAAAD8",
    x"2ADA557E",
    x"2ADA0046",
    x"2AD9AB2E",
    x"2AD95638",
    x"2AD90163",
    x"2AD8ACAF",
    x"2AD8581C",
    x"2AD803AA",
    x"2AD7AF59",
    x"2AD75B29",
    x"2AD7071A",
    x"2AD6B32B",
    x"2AD65F5E",
    x"2AD60BB1",
    x"2AD5B825",
    x"2AD564B9",
    x"2AD5116E",
    x"2AD4BE43",
    x"2AD46B39",
    x"2AD4184F",
    x"2AD3C586",
    x"2AD372DD",
    x"2AD32054",
    x"2AD2CDEC",
    x"2AD27BA4",
    x"2AD2297B",
    x"2AD1D773",
    x"2AD1858B",
    x"2AD133C3",
    x"2AD0E21A",
    x"2AD09092",
    x"2AD03F2A",
    x"2ACFEDE1",
    x"2ACF9CB8",
    x"2ACF4BAE",
    x"2ACEFAC5",
    x"2ACEA9FA",
    x"2ACE5950",
    x"2ACE08C5",
    x"2ACDB859",
    x"2ACD680D",
    x"2ACD17E0",
    x"2ACCC7D2",
    x"2ACC77E3",
    x"2ACC2814",
    x"2ACBD864",
    x"2ACB88D3",
    x"2ACB3961",
    x"2ACAEA0E",
    x"2ACA9ADA",
    x"2ACA4BC5",
    x"2AC9FCCF",
    x"2AC9ADF8",
    x"2AC95F3F",
    x"2AC910A5",
    x"2AC8C22A",
    x"2AC873CE",
    x"2AC82590",
    x"2AC7D770",
    x"2AC7896F",
    x"2AC73B8D",
    x"2AC6EDC9",
    x"2AC6A023",
    x"2AC6529C",
    x"2AC60533",
    x"2AC5B7E8",
    x"2AC56ABB",
    x"2AC51DAC",
    x"2AC4D0BC",
    x"2AC483E9",
    x"2AC43735",
    x"2AC3EA9E",
    x"2AC39E25",
    x"2AC351CA",
    x"2AC3058D",
    x"2AC2B96E",
    x"2AC26D6C",
    x"2AC22189",
    x"2AC1D5C2",
    x"2AC18A1A",
    x"2AC13E8E",
    x"2AC0F321",
    x"2AC0A7D0",
    x"2AC05C9E",
    x"2AC01188",
    x"2ABFC690",
    x"2ABF7BB5",
    x"2ABF30F7",
    x"2ABEE657",
    x"2ABE9BD3",
    x"2ABE516D",
    x"2ABE0724",
    x"2ABDBCF7",
    x"2ABD72E8",
    x"2ABD28F5",
    x"2ABCDF20",
    x"2ABC9567",
    x"2ABC4BCB",
    x"2ABC024C",
    x"2ABBB8E9",
    x"2ABB6FA3",
    x"2ABB267A",
    x"2ABADD6D",
    x"2ABA947D",
    x"2ABA4BA9",
    x"2ABA02F2",
    x"2AB9BA57",
    x"2AB971D8",
    x"2AB92976",
    x"2AB8E130",
    x"2AB89906",
    x"2AB850F8",
    x"2AB80907",
    x"2AB7C131",
    x"2AB77978",
    x"2AB731DA",
    x"2AB6EA59",
    x"2AB6A2F3",
    x"2AB65BAA",
    x"2AB6147C",
    x"2AB5CD6A",
    x"2AB58673",
    x"2AB53F99",
    x"2AB4F8DA",
    x"2AB4B236",
    x"2AB46BAE",
    x"2AB42542",
    x"2AB3DEF1",
    x"2AB398BC",
    x"2AB352A2",
    x"2AB30CA3",
    x"2AB2C6C0",
    x"2AB280F8",
    x"2AB23B4B",
    x"2AB1F5BA",
    x"2AB1B043",
    x"2AB16AE8",
    x"2AB125A8",
    x"2AB0E082",
    x"2AB09B78",
    x"2AB05689",
    x"2AB011B5",
    x"2AAFCCFB",
    x"2AAF885C",
    x"2AAF43D9",
    x"2AAEFF6F",
    x"2AAEBB21",
    x"2AAE76ED",
    x"2AAE32D4",
    x"2AADEED6",
    x"2AADAAF1",
    x"2AAD6728",
    x"2AAD2379",
    x"2AACDFE4",
    x"2AAC9C6A",
    x"2AAC590A",
    x"2AAC15C4",
    x"2AABD299",
    x"2AAB8F88",
    x"2AAB4C91",
    x"2AAB09B4",
    x"2AAAC6F1",
    x"2AAA8449",
    x"2AAA41BA",
    x"2AA9FF45",
    x"2AA9BCEA",
    x"2AA97AAA",
    x"2AA93883",
    x"2AA8F675",
    x"2AA8B482",
    x"2AA872A8",
    x"2AA830E8",
    x"2AA7EF42",
    x"2AA7ADB6",
    x"2AA76C42",
    x"2AA72AE9",
    x"2AA6E9A9",
    x"2AA6A882",
    x"2AA66775",
    x"2AA62682",
    x"2AA5E5A7",
    x"2AA5A4E6",
    x"2AA5643E",
    x"2AA523B0",
    x"2AA4E33A",
    x"2AA4A2DE",
    x"2AA4629B",
    x"2AA42271",
    x"2AA3E260",
    x"2AA3A268",
    x"2AA36289",
    x"2AA322C3",
    x"2AA2E316",
    x"2AA2A382",
    x"2AA26406",
    x"2AA224A4",
    x"2AA1E55A",
    x"2AA1A629",
    x"2AA16710",
    x"2AA12810",
    x"2AA0E929",
    x"2AA0AA5A",
    x"2AA06BA4",
    x"2AA02D06",
    x"2A9FEE80",
    x"2A9FB013",
    x"2A9F71BF",
    x"2A9F3383",
    x"2A9EF55F",
    x"2A9EB753",
    x"2A9E795F",
    x"2A9E3B84",
    x"2A9DFDC1",
    x"2A9DC016",
    x"2A9D8283",
    x"2A9D4508",
    x"2A9D07A5",
    x"2A9CCA5A",
    x"2A9C8D27",
    x"2A9C500C",
    x"2A9C1308",
    x"2A9BD61D",
    x"2A9B9949",
    x"2A9B5C8D",
    x"2A9B1FE9",
    x"2A9AE35C",
    x"2A9AA6E7",
    x"2A9A6A8A",
    x"2A9A2E44",
    x"2A99F215",
    x"2A99B5FF",
    x"2A9979FF",
    x"2A993E17",
    x"2A990247",
    x"2A98C68D",
    x"2A988AEC",
    x"2A984F61",
    x"2A9813ED",
    x"2A97D891",
    x"2A979D4C",
    x"2A97621E",
    x"2A972708",
    x"2A96EC08",
    x"2A96B11F",
    x"2A96764E",
    x"2A963B93",
    x"2A9600EF",
    x"2A95C662",
    x"2A958BEC",
    x"2A95518D",
    x"2A951744",
    x"2A94DD13",
    x"2A94A2F8",
    x"2A9468F3",
    x"2A942F06",
    x"2A93F52E",
    x"2A93BB6E",
    x"2A9381C4",
    x"2A934831",
    x"2A930EB4",
    x"2A92D54D",
    x"2A929BFD",
    x"2A9262C3",
    x"2A9229A0",
    x"2A91F093",
    x"2A91B79C",
    x"2A917EBB",
    x"2A9145F1",
    x"2A910D3D",
    x"2A90D49E",
    x"2A909C16",
    x"2A9063A4",
    x"2A902B49",
    x"2A8FF303",
    x"2A8FBAD3",
    x"2A8F82B9",
    x"2A8F4AB5",
    x"2A8F12C6",
    x"2A8EDAEE",
    x"2A8EA32B",
    x"2A8E6B7E",
    x"2A8E33E7",
    x"2A8DFC66",
    x"2A8DC4FA",
    x"2A8D8DA4",
    x"2A8D5663",
    x"2A8D1F38",
    x"2A8CE823",
    x"2A8CB123",
    x"2A8C7A39",
    x"2A8C4364",
    x"2A8C0CA4",
    x"2A8BD5FA",
    x"2A8B9F65",
    x"2A8B68E5",
    x"2A8B327B",
    x"2A8AFC26",
    x"2A8AC5E6",
    x"2A8A8FBB",
    x"2A8A59A6",
    x"2A8A23A5",
    x"2A89EDBA",
    x"2A89B7E3",
    x"2A898222",
    x"2A894C76",
    x"2A8916DE",
    x"2A88E15C",
    x"2A88ABEE",
    x"2A887695",
    x"2A884152",
    x"2A880C22",
    x"2A87D708",
    x"2A87A202",
    x"2A876D11",
    x"2A873835",
    x"2A87036E",
    x"2A86CEBA",
    x"2A869A1C",
    x"2A866592",
    x"2A86311D",
    x"2A85FCBC",
    x"2A85C86F",
    x"2A859437",
    x"2A856013",
    x"2A852C04",
    x"2A84F809",
    x"2A84C422",
    x"2A849050",
    x"2A845C91",
    x"2A8428E7",
    x"2A83F552",
    x"2A83C1D0",
    x"2A838E62",
    x"2A835B08",
    x"2A8327C3",
    x"2A82F491",
    x"2A82C174",
    x"2A828E6A",
    x"2A825B75",
    x"2A822893",
    x"2A81F5C5",
    x"2A81C30B",
    x"2A819065",
    x"2A815DD2",
    x"2A812B53",
    x"2A80F8E8",
    x"2A80C691",
    x"2A80944D",
    x"2A80621D",
    x"2A803000",
    x"2A7FFBEF",
    x"2A7F9804",
    x"2A7F3440",
    x"2A7ED0A3",
    x"2A7E6D2D",
    x"2A7E09DE",
    x"2A7DA6B5",
    x"2A7D43B3",
    x"2A7CE0D8",
    x"2A7C7E24",
    x"2A7C1B96",
    x"2A7BB92E",
    x"2A7B56ED",
    x"2A7AF4D2",
    x"2A7A92DE",
    x"2A7A310F",
    x"2A79CF67",
    x"2A796DE5",
    x"2A790C89",
    x"2A78AB54",
    x"2A784A44",
    x"2A77E95A",
    x"2A778895",
    x"2A7727F7",
    x"2A76C77E",
    x"2A76672B",
    x"2A7606FD",
    x"2A75A6F5",
    x"2A754713",
    x"2A74E756",
    x"2A7487BE",
    x"2A74284C",
    x"2A73C8FF",
    x"2A7369D7",
    x"2A730AD4",
    x"2A72ABF6",
    x"2A724D3E",
    x"2A71EEAA",
    x"2A71903B",
    x"2A7131F1",
    x"2A70D3CC",
    x"2A7075CC",
    x"2A7017F0",
    x"2A6FBA39",
    x"2A6F5CA7",
    x"2A6EFF39",
    x"2A6EA1EF",
    x"2A6E44CA",
    x"2A6DE7C9",
    x"2A6D8AED",
    x"2A6D2E35",
    x"2A6CD1A1",
    x"2A6C7531",
    x"2A6C18E5",
    x"2A6BBCBE",
    x"2A6B60BA",
    x"2A6B04DA",
    x"2A6AA91E",
    x"2A6A4D86",
    x"2A69F211",
    x"2A6996C1",
    x"2A693B94",
    x"2A68E08A",
    x"2A6885A4",
    x"2A682AE2",
    x"2A67D043",
    x"2A6775C7",
    x"2A671B6F",
    x"2A66C13A",
    x"2A666728",
    x"2A660D39",
    x"2A65B36D",
    x"2A6559C5",
    x"2A65003F",
    x"2A64A6DD",
    x"2A644D9D",
    x"2A63F480",
    x"2A639B86",
    x"2A6342AE",
    x"2A62E9FA",
    x"2A629168",
    x"2A6238F8",
    x"2A61E0AB",
    x"2A618881",
    x"2A613078",
    x"2A60D893",
    x"2A6080CF",
    x"2A60292E",
    x"2A5FD1AF",
    x"2A5F7A52",
    x"2A5F2317",
    x"2A5ECBFF",
    x"2A5E7508",
    x"2A5E1E33",
    x"2A5DC780",
    x"2A5D70EF",
    x"2A5D1A80",
    x"2A5CC433",
    x"2A5C6E07",
    x"2A5C17FD",
    x"2A5BC214",
    x"2A5B6C4D",
    x"2A5B16A7",
    x"2A5AC123",
    x"2A5A6BC1",
    x"2A5A167F",
    x"2A59C15F",
    x"2A596C60",
    x"2A591782",
    x"2A58C2C6",
    x"2A586E2A",
    x"2A5819B0",
    x"2A57C556",
    x"2A57711D",
    x"2A571D06",
    x"2A56C90F",
    x"2A567539",
    x"2A562183",
    x"2A55CDEE",
    x"2A557A7A",
    x"2A552727",
    x"2A54D3F4",
    x"2A5480E1",
    x"2A542DEF",
    x"2A53DB1D",
    x"2A53886C",
    x"2A5335DB",
    x"2A52E36A",
    x"2A529119",
    x"2A523EE8",
    x"2A51ECD8",
    x"2A519AE7",
    x"2A514917",
    x"2A50F766",
    x"2A50A5D5",
    x"2A505465",
    x"2A500313",
    x"2A4FB1E2",
    x"2A4F60D0",
    x"2A4F0FDE",
    x"2A4EBF0C",
    x"2A4E6E59",
    x"2A4E1DC6",
    x"2A4DCD52",
    x"2A4D7CFD",
    x"2A4D2CC8",
    x"2A4CDCB2",
    x"2A4C8CBC",
    x"2A4C3CE4",
    x"2A4BED2C",
    x"2A4B9D93",
    x"2A4B4E19",
    x"2A4AFEBE",
    x"2A4AAF82",
    x"2A4A6065",
    x"2A4A1167",
    x"2A49C287",
    x"2A4973C7",
    x"2A492525",
    x"2A48D6A2",
    x"2A48883D",
    x"2A4839F7",
    x"2A47EBD0",
    x"2A479DC7",
    x"2A474FDD",
    x"2A470211",
    x"2A46B463",
    x"2A4666D4",
    x"2A461963",
    x"2A45CC10",
    x"2A457EDB",
    x"2A4531C5",
    x"2A44E4CC",
    x"2A4497F2",
    x"2A444B36",
    x"2A43FE97",
    x"2A43B217",
    x"2A4365B4",
    x"2A43196F",
    x"2A42CD48",
    x"2A42813F",
    x"2A423553",
    x"2A41E985",
    x"2A419DD5",
    x"2A415242",
    x"2A4106CC",
    x"2A40BB74",
    x"2A40703A",
    x"2A40251D",
    x"2A3FDA1D",
    x"2A3F8F3A",
    x"2A3F4475",
    x"2A3EF9CD",
    x"2A3EAF42",
    x"2A3E64D4",
    x"2A3E1A83",
    x"2A3DD04F",
    x"2A3D8638",
    x"2A3D3C3E",
    x"2A3CF261",
    x"2A3CA8A1",
    x"2A3C5EFD",
    x"2A3C1577",
    x"2A3BCC0D",
    x"2A3B82BF",
    x"2A3B398F",
    x"2A3AF07A",
    x"2A3AA783",
    x"2A3A5EA7",
    x"2A3A15E9",
    x"2A39CD46",
    x"2A3984C0",
    x"2A393C57",
    x"2A38F409",
    x"2A38ABD8",
    x"2A3863C3",
    x"2A381BCA",
    x"2A37D3ED",
    x"2A378C2C",
    x"2A374488",
    x"2A36FCFF",
    x"2A36B592",
    x"2A366E41",
    x"2A36270C",
    x"2A35DFF2",
    x"2A3598F5",
    x"2A355213",
    x"2A350B4D",
    x"2A34C4A2",
    x"2A347E13",
    x"2A3437A0",
    x"2A33F148",
    x"2A33AB0B",
    x"2A3364EA",
    x"2A331EE4",
    x"2A32D8FA",
    x"2A32932B",
    x"2A324D77",
    x"2A3207DE",
    x"2A31C261",
    x"2A317CFE",
    x"2A3137B7",
    x"2A30F28B",
    x"2A30AD79",
    x"2A306883",
    x"2A3023A8",
    x"2A2FDEE7",
    x"2A2F9A42",
    x"2A2F55B7",
    x"2A2F1147",
    x"2A2ECCF1",
    x"2A2E88B7",
    x"2A2E4496",
    x"2A2E0091",
    x"2A2DBCA6",
    x"2A2D78D6",
    x"2A2D3520",
    x"2A2CF184",
    x"2A2CAE03",
    x"2A2C6A9C",
    x"2A2C2750",
    x"2A2BE41D",
    x"2A2BA105",
    x"2A2B5E08",
    x"2A2B1B24",
    x"2A2AD85A",
    x"2A2A95AB",
    x"2A2A5315",
    x"2A2A109A",
    x"2A29CE38",
    x"2A298BF1",
    x"2A2949C3",
    x"2A2907AF",
    x"2A28C5B5",
    x"2A2883D5",
    x"2A28420E",
    x"2A280061",
    x"2A27BECE",
    x"2A277D54",
    x"2A273BF4",
    x"2A26FAAD",
    x"2A26B980",
    x"2A26786C",
    x"2A263772",
    x"2A25F691",
    x"2A25B5C9",
    x"2A25751B",
    x"2A253486",
    x"2A24F40A",
    x"2A24B3A7",
    x"2A24735D",
    x"2A24332D",
    x"2A23F315",
    x"2A23B317",
    x"2A237332",
    x"2A233365",
    x"2A22F3B1",
    x"2A22B417",
    x"2A227495",
    x"2A22352C",
    x"2A21F5DB",
    x"2A21B6A3",
    x"2A217784",
    x"2A21387E",
    x"2A20F990",
    x"2A20BABB",
    x"2A207BFE",
    x"2A203D5A",
    x"2A1FFECE",
    x"2A1FC05B",
    x"2A1F8200",
    x"2A1F43BE",
    x"2A1F0593",
    x"2A1EC781",
    x"2A1E8987",
    x"2A1E4BA6",
    x"2A1E0DDC",
    x"2A1DD02B",
    x"2A1D9292",
    x"2A1D5510",
    x"2A1D17A7",
    x"2A1CDA56",
    x"2A1C9D1D",
    x"2A1C5FFB",
    x"2A1C22F2",
    x"2A1BE600",
    x"2A1BA926",
    x"2A1B6C64",
    x"2A1B2FB9",
    x"2A1AF326",
    x"2A1AB6AB",
    x"2A1A7A48",
    x"2A1A3DFC",
    x"2A1A01C7",
    x"2A19C5AA",
    x"2A1989A5",
    x"2A194DB7",
    x"2A1911E0",
    x"2A18D621",
    x"2A189A79",
    x"2A185EE8",
    x"2A18236F",
    x"2A17E80C",
    x"2A17ACC1",
    x"2A17718D",
    x"2A173671",
    x"2A16FB6B",
    x"2A16C07C",
    x"2A1685A4",
    x"2A164AE4",
    x"2A16103A",
    x"2A15D5A7",
    x"2A159B2B",
    x"2A1560C6",
    x"2A152677",
    x"2A14EC40",
    x"2A14B21F",
    x"2A147815",
    x"2A143E21",
    x"2A140444",
    x"2A13CA7E",
    x"2A1390CE",
    x"2A135734",
    x"2A131DB2",
    x"2A12E445",
    x"2A12AAEF",
    x"2A1271B0",
    x"2A123886",
    x"2A11FF74",
    x"2A11C677",
    x"2A118D90",
    x"2A1154C0",
    x"2A111C06",
    x"2A10E362",
    x"2A10AAD5",
    x"2A10725D",
    x"2A1039FB",
    x"2A1001B0",
    x"2A0FC97A",
    x"2A0F915A",
    x"2A0F5950",
    x"2A0F215C",
    x"2A0EE97E",
    x"2A0EB1B6",
    x"2A0E7A03",
    x"2A0E4267",
    x"2A0E0AE0",
    x"2A0DD36E",
    x"2A0D9C12",
    x"2A0D64CC",
    x"2A0D2D9C",
    x"2A0CF681",
    x"2A0CBF7B",
    x"2A0C888B",
    x"2A0C51B0",
    x"2A0C1AEB",
    x"2A0BE43B",
    x"2A0BADA1",
    x"2A0B771C",
    x"2A0B40AC",
    x"2A0B0A51",
    x"2A0AD40C",
    x"2A0A9DDB",
    x"2A0A67C0",
    x"2A0A31BA",
    x"2A09FBC9",
    x"2A09C5EE",
    x"2A099027",
    x"2A095A75",
    x"2A0924D8",
    x"2A08EF50",
    x"2A08B9DD",
    x"2A08847F",
    x"2A084F36",
    x"2A081A01",
    x"2A07E4E1",
    x"2A07AFD6",
    x"2A077AE0",
    x"2A0745FE",
    x"2A071131",
    x"2A06DC79",
    x"2A06A7D5",
    x"2A067346",
    x"2A063ECB",
    x"2A060A65",
    x"2A05D613",
    x"2A05A1D5",
    x"2A056DAC",
    x"2A053998",
    x"2A050597",
    x"2A04D1AB",
    x"2A049DD3",
    x"2A046A10",
    x"2A043661",
    x"2A0402C5",
    x"2A03CF3E",
    x"2A039BCC",
    x"2A03686D",
    x"2A033522",
    x"2A0301EB",
    x"2A02CEC8",
    x"2A029BBA",
    x"2A0268BF",
    x"2A0235D8",
    x"2A020305",
    x"2A01D045",
    x"2A019D9A",
    x"2A016B02",
    x"2A01387E",
    x"2A01060E",
    x"2A00D3B2",
    x"2A00A169",
    x"2A006F34",
    x"2A003D12",
    x"2A000B04",
    x"29FFB212",
    x"29FF4E44",
    x"29FEEA9D",
    x"29FE871D",
    x"29FE23C4",
    x"29FDC091",
    x"29FD5D85",
    x"29FCFAA0",
    x"29FC97E1",
    x"29FC3549",
    x"29FBD2D8",
    x"29FB708D",
    x"29FB0E68",
    x"29FAAC69",
    x"29FA4A91",
    x"29F9E8DF",
    x"29F98753",
    x"29F925ED",
    x"29F8C4AE",
    x"29F86394",
    x"29F802A0",
    x"29F7A1D2",
    x"29F74129",
    x"29F6E0A7",
    x"29F6804A",
    x"29F62012",
    x"29F5C001",
    x"29F56014",
    x"29F5004E",
    x"29F4A0AC",
    x"29F44130",
    x"29F3E1D9",
    x"29F382A8",
    x"29F3239B",
    x"29F2C4B4",
    x"29F265F1",
    x"29F20754",
    x"29F1A8DC",
    x"29F14A88",
    x"29F0EC59",
    x"29F08E50",
    x"29F0306A",
    x"29EFD2AA",
    x"29EF750E",
    x"29EF1796",
    x"29EEBA43",
    x"29EE5D15",
    x"29EE000A",
    x"29EDA325",
    x"29ED4663",
    x"29ECE9C6",
    x"29EC8D4C",
    x"29EC30F7",
    x"29EBD4C6",
    x"29EB78B9",
    x"29EB1CD0",
    x"29EAC10A",
    x"29EA6569",
    x"29EA09EB",
    x"29E9AE91",
    x"29E9535B",
    x"29E8F848",
    x"29E89D59",
    x"29E8428D",
    x"29E7E7E5",
    x"29E78D60",
    x"29E732FE",
    x"29E6D8C0",
    x"29E67EA5",
    x"29E624AD",
    x"29E5CAD8",
    x"29E57127",
    x"29E51798",
    x"29E4BE2C",
    x"29E464E3",
    x"29E40BBD",
    x"29E3B2BA",
    x"29E359DA",
    x"29E3011C",
    x"29E2A881",
    x"29E25008",
    x"29E1F7B2",
    x"29E19F7F",
    x"29E1476E",
    x"29E0EF7F",
    x"29E097B2",
    x"29E04008",
    x"29DFE880",
    x"29DF911B",
    x"29DF39D7",
    x"29DEE2B5",
    x"29DE8BB6",
    x"29DE34D8",
    x"29DDDE1D",
    x"29DD8783",
    x"29DD310B",
    x"29DCDAB4",
    x"29DC8480",
    x"29DC2E6D",
    x"29DBD87C",
    x"29DB82AC",
    x"29DB2CFD",
    x"29DAD771",
    x"29DA8205",
    x"29DA2CBB",
    x"29D9D792",
    x"29D9828B",
    x"29D92DA4",
    x"29D8D8DF",
    x"29D8843B",
    x"29D82FB8",
    x"29D7DB55",
    x"29D78714",
    x"29D732F4",
    x"29D6DEF4",
    x"29D68B16",
    x"29D63758",
    x"29D5E3BA",
    x"29D5903E",
    x"29D53CE2",
    x"29D4E9A6",
    x"29D4968B",
    x"29D44391",
    x"29D3F0B6",
    x"29D39DFC",
    x"29D34B63",
    x"29D2F8EA",
    x"29D2A690",
    x"29D25457",
    x"29D2023F",
    x"29D1B046",
    x"29D15E6D",
    x"29D10CB4",
    x"29D0BB1B",
    x"29D069A2",
    x"29D01848",
    x"29CFC70F",
    x"29CF75F5",
    x"29CF24FB",
    x"29CED420",
    x"29CE8365",
    x"29CE32C9",
    x"29CDE24D",
    x"29CD91F0",
    x"29CD41B3",
    x"29CCF195",
    x"29CCA196",
    x"29CC51B7",
    x"29CC01F6",
    x"29CBB255",
    x"29CB62D3",
    x"29CB1370",
    x"29CAC42C",
    x"29CA7507",
    x"29CA2600",
    x"29C9D719",
    x"29C98850",
    x"29C939A7",
    x"29C8EB1B",
    x"29C89CAF",
    x"29C84E61",
    x"29C80032",
    x"29C7B221",
    x"29C7642E",
    x"29C7165A",
    x"29C6C8A5",
    x"29C67B0E",
    x"29C62D95",
    x"29C5E03A",
    x"29C592FE",
    x"29C545DF",
    x"29C4F8DF",
    x"29C4ABFD",
    x"29C45F39",
    x"29C41292",
    x"29C3C60A",
    x"29C379A0",
    x"29C32D53",
    x"29C2E124",
    x"29C29513",
    x"29C24920",
    x"29C1FD4A",
    x"29C1B192",
    x"29C165F7",
    x"29C11A7A",
    x"29C0CF1B",
    x"29C083D8",
    x"29C038B4",
    x"29BFEDAC",
    x"29BFA2C2",
    x"29BF57F5",
    x"29BF0D45",
    x"29BEC2B2",
    x"29BE783D",
    x"29BE2DE5",
    x"29BDE3A9",
    x"29BD998B",
    x"29BD4F89",
    x"29BD05A5",
    x"29BCBBDD",
    x"29BC7232",
    x"29BC28A3",
    x"29BBDF32",
    x"29BB95DD",
    x"29BB4CA5",
    x"29BB0389",
    x"29BABA8A",
    x"29BA71A7",
    x"29BA28E1",
    x"29B9E038",
    x"29B997AA",
    x"29B94F39",
    x"29B906E4",
    x"29B8BEAC",
    x"29B8768F",
    x"29B82E8F",
    x"29B7E6AB",
    x"29B79EE3",
    x"29B75737",
    x"29B70FA7",
    x"29B6C832",
    x"29B680DA",
    x"29B6399E",
    x"29B5F27D",
    x"29B5AB78",
    x"29B5648F",
    x"29B51DC2",
    x"29B4D710",
    x"29B4907A",
    x"29B449FF",
    x"29B403A0",
    x"29B3BD5C",
    x"29B37734",
    x"29B33127",
    x"29B2EB36",
    x"29B2A55F",
    x"29B25FA4",
    x"29B21A05",
    x"29B1D480",
    x"29B18F17",
    x"29B149C8",
    x"29B10495",
    x"29B0BF7D",
    x"29B07A7F",
    x"29B0359D",
    x"29AFF0D5",
    x"29AFAC29",
    x"29AF6797",
    x"29AF2320",
    x"29AEDEC3",
    x"29AE9A82",
    x"29AE565B",
    x"29AE124E",
    x"29ADCE5C",
    x"29AD8A85",
    x"29AD46C8",
    x"29AD0326",
    x"29ACBF9E",
    x"29AC7C30",
    x"29AC38DD",
    x"29ABF5A4",
    x"29ABB285",
    x"29AB6F80",
    x"29AB2C96",
    x"29AAE9C5",
    x"29AAA70F",
    x"29AA6473",
    x"29AA21F0",
    x"29A9DF88",
    x"29A99D3A",
    x"29A95B05",
    x"29A918EB",
    x"29A8D6EA",
    x"29A89503",
    x"29A85335",
    x"29A81182",
    x"29A7CFE8",
    x"29A78E67",
    x"29A74D00",
    x"29A70BB3",
    x"29A6CA7F",
    x"29A68965",
    x"29A64864",
    x"29A6077C",
    x"29A5C6AE",
    x"29A585F9",
    x"29A5455D",
    x"29A504DB",
    x"29A4C472",
    x"29A48421",
    x"29A443EA",
    x"29A403CC",
    x"29A3C3C7",
    x"29A383DB",
    x"29A34408",
    x"29A3044E",
    x"29A2C4AD",
    x"29A28525",
    x"29A245B5",
    x"29A2065E",
    x"29A1C720",
    x"29A187FB",
    x"29A148EE",
    x"29A109FA",
    x"29A0CB1E",
    x"29A08C5B",
    x"29A04DB0",
    x"29A00F1E",
    x"299FD0A4",
    x"299F9243",
    x"299F53FA",
    x"299F15C9",
    x"299ED7B1",
    x"299E99B1",
    x"299E5BC9",
    x"299E1DF9",
    x"299DE042",
    x"299DA2A2",
    x"299D651B",
    x"299D27AB",
    x"299CEA54",
    x"299CAD14",
    x"299C6FEC",
    x"299C32DC",
    x"299BF5E5",
    x"299BB904",
    x"299B7C3C",
    x"299B3F8B",
    x"299B02F2",
    x"299AC671",
    x"299A8A07",
    x"299A4DB5",
    x"299A117B",
    x"2999D557",
    x"2999994C",
    x"29995D58",
    x"2999217B",
    x"2998E5B6",
    x"2998AA07",
    x"29986E71",
    x"299832F1",
    x"2997F789",
    x"2997BC38",
    x"299780FE",
    x"299745DB",
    x"29970ACF",
    x"2996CFDB",
    x"299694FD",
    x"29965A36",
    x"29961F86",
    x"2995E4ED",
    x"2995AA6B",
    x"29957000",
    x"299535AC",
    x"2994FB6E",
    x"2994C148",
    x"29948737",
    x"29944D3E",
    x"2994135B",
    x"2993D98F",
    x"29939FD9",
    x"2993663A",
    x"29932CB1",
    x"2992F33F",
    x"2992B9E3",
    x"2992809E",
    x"2992476F",
    x"29920E56",
    x"2991D553",
    x"29919C67",
    x"29916391",
    x"29912AD1",
    x"2990F228",
    x"2990B994",
    x"29908117",
    x"299048AF",
    x"2990105E",
    x"298FD823",
    x"298F9FFD",
    x"298F67EE",
    x"298F2FF4",
    x"298EF810",
    x"298EC042",
    x"298E888A",
    x"298E50E7",
    x"298E195B",
    x"298DE1E4",
    x"298DAA82",
    x"298D7336",
    x"298D3C00",
    x"298D04DF",
    x"298CCDD4",
    x"298C96DF",
    x"298C5FFE",
    x"298C2934",
    x"298BF27E",
    x"298BBBDE",
    x"298B8553",
    x"298B4EDE",
    x"298B187E",
    x"298AE233",
    x"298AABFD",
    x"298A75DC",
    x"298A3FD1",
    x"298A09DB",
    x"2989D3F9",
    x"29899E2D",
    x"29896876",
    x"298932D3",
    x"2988FD46",
    x"2988C7CE",
    x"2988926A",
    x"29885D1B",
    x"298827E1",
    x"2987F2BC",
    x"2987BDAB",
    x"298788B0",
    x"298753C9",
    x"29871EF6",
    x"2986EA39",
    x"2986B58F",
    x"298680FB",
    x"29864C7B",
    x"2986180F",
    x"2985E3B8",
    x"2985AF75",
    x"29857B47",
    x"2985472D",
    x"29851327",
    x"2984DF36",
    x"2984AB59",
    x"29847790",
    x"298443DB",
    x"2984103B",
    x"2983DCAF",
    x"2983A936",
    x"298375D2",
    x"29834282",
    x"29830F46",
    x"2982DC1E",
    x"2982A90A",
    x"2982760A",
    x"2982431E",
    x"29821046",
    x"2981DD81",
    x"2981AAD1",
    x"29817834",
    x"298145AB",
    x"29811336",
    x"2980E0D4",
    x"2980AE86",
    x"29807C4B",
    x"29804A25",
    x"29801812",
    x"297FCC24",
    x"297F684C",
    x"297F049A",
    x"297EA110",
    x"297E3DAC",
    x"297DDA70",
    x"297D775A",
    x"297D146B",
    x"297CB1A2",
    x"297C4F00",
    x"297BEC84",
    x"297B8A2F",
    x"297B2800",
    x"297AC5F8",
    x"297A6415",
    x"297A0259",
    x"2979A0C4",
    x"29793F54",
    x"2978DE0A",
    x"29787CE6",
    x"29781BE9",
    x"2977BB11",
    x"29775A5E",
    x"2976F9D2",
    x"2976996B",
    x"2976392A",
    x"2975D90E",
    x"29757918",
    x"29751948",
    x"2974B99D",
    x"29745A17",
    x"2973FAB6",
    x"29739B7B",
    x"29733C65",
    x"2972DD74",
    x"29727EA8",
    x"29722001",
    x"2971C17F",
    x"29716322",
    x"297104E9",
    x"2970A6D6",
    x"297048E7",
    x"296FEB1D",
    x"296F8D77",
    x"296F2FF6",
    x"296ED29A",
    x"296E7562",
    x"296E184E",
    x"296DBB5F",
    x"296D5E94",
    x"296D01ED",
    x"296CA56A",
    x"296C490C",
    x"296BECD1",
    x"296B90BA",
    x"296B34C8",
    x"296AD8F9",
    x"296A7D4E",
    x"296A21C7",
    x"2969C664",
    x"29696B24",
    x"29691008",
    x"2968B510",
    x"29685A3B",
    x"2967FF89",
    x"2967A4FB",
    x"29674A90",
    x"2966F049",
    x"29669625",
    x"29663C24",
    x"2965E246",
    x"2965888B",
    x"29652EF3",
    x"2964D57E",
    x"29647C2C",
    x"296422FD",
    x"2963C9F1",
    x"29637107",
    x"29631840",
    x"2962BF9C",
    x"2962671B",
    x"29620EBC",
    x"2961B67F",
    x"29615E65",
    x"2961066D",
    x"2960AE98",
    x"296056E5",
    x"295FFF54",
    x"295FA7E6",
    x"295F5099",
    x"295EF96F",
    x"295EA266",
    x"295E4B80",
    x"295DF4BB",
    x"295D9E18",
    x"295D4798",
    x"295CF138",
    x"295C9AFB",
    x"295C44DF",
    x"295BEEE5",
    x"295B990D",
    x"295B4356",
    x"295AEDC0",
    x"295A984C",
    x"295A42F9",
    x"2959EDC8",
    x"295998B7",
    x"295943C8",
    x"2958EEFA",
    x"29589A4E",
    x"295845C2",
    x"2957F157",
    x"29579D0D",
    x"295748E4",
    x"2956F4DC",
    x"2956A0F5",
    x"29564D2E",
    x"2955F989",
    x"2955A604",
    x"2955529F",
    x"2954FF5B",
    x"2954AC37",
    x"29545934",
    x"29540652",
    x"2953B38F",
    x"295360ED",
    x"29530E6C",
    x"2952BC0A",
    x"295269C9",
    x"295217A8",
    x"2951C5A6",
    x"295173C5",
    x"29512204",
    x"2950D062",
    x"29507EE1",
    x"29502D7F",
    x"294FDC3D",
    x"294F8B1B",
    x"294F3A19",
    x"294EE936",
    x"294E9873",
    x"294E47CF",
    x"294DF74A",
    x"294DA6E6",
    x"294D56A0",
    x"294D067A",
    x"294CB673",
    x"294C668B",
    x"294C16C3",
    x"294BC719",
    x"294B778F",
    x"294B2824",
    x"294AD8D8",
    x"294A89AB",
    x"294A3A9C",
    x"2949EBAD",
    x"29499CDC",
    x"29494E2A",
    x"2948FF97",
    x"2948B123",
    x"294862CD",
    x"29481495",
    x"2947C67D",
    x"29477882",
    x"29472AA6",
    x"2946DCE9",
    x"29468F4A",
    x"294641C9",
    x"2945F466",
    x"2945A722",
    x"294559FC",
    x"29450CF4",
    x"2944C00A",
    x"2944733E",
    x"29442690",
    x"2943DA00",
    x"29438D8D",
    x"29434139",
    x"2942F502",
    x"2942A8EA",
    x"29425CEE",
    x"29421111",
    x"2941C551",
    x"294179AF",
    x"29412E2A",
    x"2940E2C3",
    x"29409779",
    x"29404C4C",
    x"2940013D",
    x"293FB64B",
    x"293F6B77",
    x"293F20BF",
    x"293ED625",
    x"293E8BA8",
    x"293E4148",
    x"293DF705",
    x"293DACDF",
    x"293D62D6",
    x"293D18EA",
    x"293CCF1A",
    x"293C8568",
    x"293C3BD2",
    x"293BF259",
    x"293BA8FD",
    x"293B5FBD",
    x"293B169A",
    x"293ACD93",
    x"293A84A9",
    x"293A3BDC",
    x"2939F32B",
    x"2939AA96",
    x"2939621D",
    x"293919C1",
    x"2938D181",
    x"2938895D",
    x"29384156",
    x"2937F96A",
    x"2937B19B",
    x"293769E8",
    x"29372250",
    x"2936DAD5",
    x"29369375",
    x"29364C32",
    x"2936050A",
    x"2935BDFE",
    x"2935770D",
    x"29353039",
    x"2934E980",
    x"2934A2E2",
    x"29345C60",
    x"293415FA",
    x"2933CFAF",
    x"29338980",
    x"2933436C",
    x"2932FD73",
    x"2932B796",
    x"293271D4",
    x"29322C2D",
    x"2931E6A1",
    x"2931A131",
    x"29315BDB",
    x"293116A1",
    x"2930D181",
    x"29308C7D",
    x"29304794",
    x"293002C5",
    x"292FBE12",
    x"292F7979",
    x"292F34FB",
    x"292EF097",
    x"292EAC4F",
    x"292E6821",
    x"292E240D",
    x"292DE014",
    x"292D9C36",
    x"292D5872",
    x"292D14C9",
    x"292CD13A",
    x"292C8DC6",
    x"292C4A6B",
    x"292C072B",
    x"292BC406",
    x"292B80FA",
    x"292B3E09",
    x"292AFB32",
    x"292AB875",
    x"292A75D2",
    x"292A3349",
    x"2929F0DA",
    x"2929AE85",
    x"29296C49",
    x"29292A28",
    x"2928E820",
    x"2928A633",
    x"2928645E",
    x"292822A4",
    x"2927E103",
    x"29279F7C",
    x"29275E0F",
    x"29271CBB",
    x"2926DB80",
    x"29269A5F",
    x"29265958",
    x"2926186A",
    x"2925D795",
    x"292596D9",
    x"29255637",
    x"292515AE",
    x"2924D53E",
    x"292494E7",
    x"292454A9",
    x"29241485",
    x"2923D479",
    x"29239487",
    x"292354AD",
    x"292314ED",
    x"2922D545",
    x"292295B6",
    x"29225640",
    x"292216E3",
    x"2921D79E",
    x"29219872",
    x"2921595F",
    x"29211A64",
    x"2920DB82",
    x"29209CB9",
    x"29205E08",
    x"29201F6F",
    x"291FE0EF",
    x"291FA288",
    x"291F6438",
    x"291F2601",
    x"291EE7E3",
    x"291EA9DC",
    x"291E6BEE",
    x"291E2E18",
    x"291DF05A",
    x"291DB2B4",
    x"291D7526",
    x"291D37B1",
    x"291CFA53",
    x"291CBD0D",
    x"291C7FDF",
    x"291C42C9",
    x"291C05CB",
    x"291BC8E5",
    x"291B8C16",
    x"291B4F5F",
    x"291B12C0",
    x"291AD638",
    x"291A99C9",
    x"291A5D70",
    x"291A2130",
    x"2919E506",
    x"2919A8F5",
    x"29196CFA",
    x"29193117",
    x"2918F54C",
    x"2918B998",
    x"29187DFB",
    x"29184275",
    x"29180707",
    x"2917CBB0",
    x"29179070",
    x"29175547",
    x"29171A35",
    x"2916DF3B",
    x"2916A457",
    x"2916698A",
    x"29162ED4",
    x"2915F436",
    x"2915B9AE",
    x"29157F3C",
    x"291544E2",
    x"29150A9F",
    x"2914D072",
    x"2914965C",
    x"29145C5C",
    x"29142274",
    x"2913E8A1",
    x"2913AEE6",
    x"29137541",
    x"29133BB2",
    x"2913023A",
    x"2912C8D8",
    x"29128F8D",
    x"29125658",
    x"29121D3A",
    x"2911E431",
    x"2911AB3F",
    x"29117264",
    x"2911399E",
    x"291100EF",
    x"2910C855",
    x"29108FD2",
    x"29105765",
    x"29101F0E",
    x"290FE6CD",
    x"290FAEA2",
    x"290F768C",
    x"290F3E8D",
    x"290F06A3",
    x"290ECED0",
    x"290E9712",
    x"290E5F6A",
    x"290E27D7",
    x"290DF05B",
    x"290DB8F3",
    x"290D81A2",
    x"290D4A66",
    x"290D1340",
    x"290CDC2F",
    x"290CA534",
    x"290C6E4E",
    x"290C377E",
    x"290C00C3",
    x"290BCA1D",
    x"290B938D",
    x"290B5D12",
    x"290B26AC",
    x"290AF05C",
    x"290ABA20",
    x"290A83FA",
    x"290A4DE9",
    x"290A17ED",
    x"2909E206",
    x"2909AC35",
    x"29097678",
    x"290940D0",
    x"29090B3D",
    x"2908D5BF",
    x"2908A056",
    x"29086B02",
    x"290835C3",
    x"29080098",
    x"2907CB82",
    x"29079681",
    x"29076195",
    x"29072CBD",
    x"2906F7FA",
    x"2906C34B",
    x"29068EB1",
    x"29065A2C",
    x"290625BB",
    x"2905F15E",
    x"2905BD16",
    x"290588E2",
    x"290554C3",
    x"290520B8",
    x"2904ECC1",
    x"2904B8DF",
    x"29048511",
    x"29045157",
    x"29041DB1",
    x"2903EA20",
    x"2903B6A3",
    x"29038339",
    x"29034FE4",
    x"29031CA3",
    x"2902E976",
    x"2902B65C",
    x"29028357",
    x"29025066",
    x"29021D88",
    x"2901EABF",
    x"2901B809",
    x"29018567",
    x"290152D9",
    x"2901205E",
    x"2900EDF7",
    x"2900BBA4",
    x"29008965",
    x"29005739",
    x"29002521",
    x"28FFE638",
    x"28FF8255",
    x"28FF1E9A",
    x"28FEBB06",
    x"28FE5798",
    x"28FDF451",
    x"28FD9131",
    x"28FD2E38",
    x"28FCCB65",
    x"28FC68B9",
    x"28FC0633",
    x"28FBA3D4",
    x"28FB419B",
    x"28FADF89",
    x"28FA7D9C",
    x"28FA1BD6",
    x"28F9BA37",
    x"28F958BD",
    x"28F8F769",
    x"28F8963C",
    x"28F83534",
    x"28F7D452",
    x"28F77396",
    x"28F71300",
    x"28F6B28F",
    x"28F65244",
    x"28F5F21F",
    x"28F5921F",
    x"28F53245",
    x"28F4D290",
    x"28F47300",
    x"28F41396",
    x"28F3B451",
    x"28F35531",
    x"28F2F636",
    x"28F29761",
    x"28F238B0",
    x"28F1DA24",
    x"28F17BBE",
    x"28F11D7C",
    x"28F0BF5E",
    x"28F06166",
    x"28F00392",
    x"28EFA5E3",
    x"28EF4859",
    x"28EEEAF3",
    x"28EE8DB1",
    x"28EE3094",
    x"28EDD39B",
    x"28ED76C7",
    x"28ED1A16",
    x"28ECBD8A",
    x"28EC6122",
    x"28EC04DE",
    x"28EBA8BE",
    x"28EB4CC3",
    x"28EAF0EA",
    x"28EA9536",
    x"28EA39A6",
    x"28E9DE39",
    x"28E982F0",
    x"28E927CB",
    x"28E8CCC9",
    x"28E871EB",
    x"28E81730",
    x"28E7BC99",
    x"28E76225",
    x"28E707D4",
    x"28E6ADA7",
    x"28E6539C",
    x"28E5F9B5",
    x"28E59FF1",
    x"28E54650",
    x"28E4ECD2",
    x"28E49377",
    x"28E43A3F",
    x"28E3E12A",
    x"28E38837",
    x"28E32F67",
    x"28E2D6BA",
    x"28E27E30",
    x"28E225C8",
    x"28E1CD82",
    x"28E1755F",
    x"28E11D5E",
    x"28E0C580",
    x"28E06DC4",
    x"28E0162A",
    x"28DFBEB3",
    x"28DF675D",
    x"28DF102A",
    x"28DEB919",
    x"28DE6229",
    x"28DE0B5C",
    x"28DDB4B0",
    x"28DD5E27",
    x"28DD07BF",
    x"28DCB179",
    x"28DC5B54",
    x"28DC0551",
    x"28DBAF70",
    x"28DB59B0",
    x"28DB0412",
    x"28DAAE95",
    x"28DA5939",
    x"28DA03FF",
    x"28D9AEE6",
    x"28D959EF",
    x"28D90518",
    x"28D8B063",
    x"28D85BCE",
    x"28D8075B",
    x"28D7B308",
    x"28D75ED7",
    x"28D70AC6",
    x"28D6B6D7",
    x"28D66308",
    x"28D60F59",
    x"28D5BBCB",
    x"28D5685E",
    x"28D51512",
    x"28D4C1E6",
    x"28D46EDA",
    x"28D41BEF",
    x"28D3C925",
    x"28D3767A",
    x"28D323F0",
    x"28D2D186",
    x"28D27F3C",
    x"28D22D13",
    x"28D1DB09",
    x"28D18920",
    x"28D13756",
    x"28D0E5AC",
    x"28D09422",
    x"28D042B9",
    x"28CFF16E",
    x"28CFA044",
    x"28CF4F39",
    x"28CEFE4E",
    x"28CEAD82",
    x"28CE5CD6",
    x"28CE0C4A",
    x"28CDBBDD",
    x"28CD6B8F",
    x"28CD1B61",
    x"28CCCB52",
    x"28CC7B62",
    x"28CC2B91",
    x"28CBDBE0",
    x"28CB8C4E",
    x"28CB3CDA",
    x"28CAED86",
    x"28CA9E51",
    x"28CA4F3A",
    x"28CA0043",
    x"28C9B16A",
    x"28C962B0",
    x"28C91415",
    x"28C8C598",
    x"28C8773B",
    x"28C828FB",
    x"28C7DADA",
    x"28C78CD8",
    x"28C73EF4",
    x"28C6F12F",
    x"28C6A388",
    x"28C655FF",
    x"28C60895",
    x"28C5BB49",
    x"28C56E1A",
    x"28C5210B",
    x"28C4D419",
    x"28C48745",
    x"28C43A8F",
    x"28C3EDF7",
    x"28C3A17D",
    x"28C35521",
    x"28C308E2",
    x"28C2BCC2",
    x"28C270BF",
    x"28C224DA",
    x"28C1D912",
    x"28C18D68",
    x"28C141DC",
    x"28C0F66D",
    x"28C0AB1B",
    x"28C05FE7",
    x"28C014D0",
    x"28BFC9D7",
    x"28BF7EFB",
    x"28BF343C",
    x"28BEE99A",
    x"28BE9F15",
    x"28BE54AD",
    x"28BE0A63",
    x"28BDC035",
    x"28BD7625",
    x"28BD2C31",
    x"28BCE25A",
    x"28BC98A0",
    x"28BC4F03",
    x"28BC0582",
    x"28BBBC1F",
    x"28BB72D7",
    x"28BB29AD",
    x"28BAE09F",
    x"28BA97AD",
    x"28BA4ED8",
    x"28BA0620",
    x"28B9BD84",
    x"28B97504",
    x"28B92CA0",
    x"28B8E459",
    x"28B89C2E",
    x"28B8541F",
    x"28B80C2C",
    x"28B7C455",
    x"28B77C9B",
    x"28B734FC",
    x"28B6ED79",
    x"28B6A612",
    x"28B65EC7",
    x"28B61798",
    x"28B5D085",
    x"28B5898D",
    x"28B542B1",
    x"28B4FBF1",
    x"28B4B54D",
    x"28B46EC4",
    x"28B42856",
    x"28B3E204",
    x"28B39BCD",
    x"28B355B2",
    x"28B30FB3",
    x"28B2C9CE",
    x"28B28405",
    x"28B23E57",
    x"28B1F8C4",
    x"28B1B34D",
    x"28B16DF0",
    x"28B128AF",
    x"28B0E388",
    x"28B09E7D",
    x"28B0598C",
    x"28B014B7",
    x"28AFCFFC",
    x"28AF8B5C",
    x"28AF46D7",
    x"28AF026D",
    x"28AEBE1D",
    x"28AE79E8",
    x"28AE35CE",
    x"28ADF1CE",
    x"28ADADE9",
    x"28AD6A1F",
    x"28AD266E",
    x"28ACE2D9",
    x"28AC9F5D",
    x"28AC5BFC",
    x"28AC18B5",
    x"28ABD589",
    x"28AB9276",
    x"28AB4F7E",
    x"28AB0CA0",
    x"28AAC9DC",
    x"28AA8733",
    x"28AA44A3",
    x"28AA022D",
    x"28A9BFD1",
    x"28A97D8F",
    x"28A93B67",
    x"28A8F959",
    x"28A8B764",
    x"28A87589",
    x"28A833C8",
    x"28A7F221",
    x"28A7B093",
    x"28A76F1F",
    x"28A72DC4",
    x"28A6EC83",
    x"28A6AB5B",
    x"28A66A4D",
    x"28A62958",
    x"28A5E87D",
    x"28A5A7BB",
    x"28A56712",
    x"28A52682",
    x"28A4E60C",
    x"28A4A5AE",
    x"28A4656A",
    x"28A4253F",
    x"28A3E52D",
    x"28A3A534",
    x"28A36554",
    x"28A3258D",
    x"28A2E5DF",
    x"28A2A649",
    x"28A266CD",
    x"28A22769",
    x"28A1E81E",
    x"28A1A8EC",
    x"28A169D2",
    x"28A12AD1",
    x"28A0EBE9",
    x"28A0AD19",
    x"28A06E61",
    x"28A02FC2",
    x"289FF13C",
    x"289FB2CE",
    x"289F7478",
    x"289F363B",
    x"289EF816",
    x"289EBA09",
    x"289E7C15",
    x"289E3E38",
    x"289E0074",
    x"289DC2C8",
    x"289D8534",
    x"289D47B8",
    x"289D0A54",
    x"289CCD08",
    x"289C8FD4",
    x"289C52B7",
    x"289C15B3",
    x"289BD8C6",
    x"289B9BF2",
    x"289B5F35",
    x"289B228F",
    x"289AE601",
    x"289AA98B",
    x"289A6D2D",
    x"289A30E6",
    x"2899F4B7",
    x"2899B89F",
    x"28997C9F",
    x"289940B6",
    x"289904E4",
    x"2898C92A",
    x"28988D87",
    x"289851FB",
    x"28981687",
    x"2897DB2A",
    x"28979FE4",
    x"289764B5",
    x"2897299D",
    x"2896EE9C",
    x"2896B3B2",
    x"289678E0",
    x"28963E24",
    x"2896037F",
    x"2895C8F1",
    x"28958E7A",
    x"2895541A",
    x"289519D0",
    x"2894DF9E",
    x"2894A582",
    x"28946B7C",
    x"2894318E",
    x"2893F7B6",
    x"2893BDF4",
    x"28938449",
    x"28934AB5",
    x"28931137",
    x"2892D7CF",
    x"28929E7E",
    x"28926544",
    x"28922C1F",
    x"2891F311",
    x"2891BA19",
    x"28918138",
    x"2891486C",
    x"28910FB7",
    x"2890D718",
    x"28909E8F",
    x"2890661C",
    x"28902DBF",
    x"288FF578",
    x"288FBD47",
    x"288F852C",
    x"288F4D27",
    x"288F1538",
    x"288EDD5F",
    x"288EA59B",
    x"288E6DED",
    x"288E3655",
    x"288DFED3",
    x"288DC766",
    x"288D900F",
    x"288D58CE",
    x"288D21A2",
    x"288CEA8B",
    x"288CB38B",
    x"288C7C9F",
    x"288C45C9",
    x"288C0F09",
    x"288BD85D",
    x"288BA1C8",
    x"288B6B47",
    x"288B34DC",
    x"288AFE86",
    x"288AC845",
    x"288A9219",
    x"288A5C03",
    x"288A2601",
    x"2889F015",
    x"2889BA3E",
    x"2889847C",
    x"28894ECE",
    x"28891936",
    x"2888E3B3",
    x"2888AE44",
    x"288878EA",
    x"288843A6",
    x"28880E76",
    x"2887D95A",
    x"2887A454",
    x"28876F62",
    x"28873A85",
    x"288705BC",
    x"2886D108",
    x"28869C69",
    x"288667DE",
    x"28863368",
    x"2885FF06",
    x"2885CAB8",
    x"2885967F",
    x"2885625B",
    x"28852E4B",
    x"2884FA4F",
    x"2884C667",
    x"28849294",
    x"28845ED5",
    x"28842B2A",
    x"2883F793",
    x"2883C410",
    x"288390A2",
    x"28835D47",
    x"28832A01",
    x"2882F6CE",
    x"2882C3B0",
    x"288290A5",
    x"28825DAF",
    x"28822ACC",
    x"2881F7FD",
    x"2881C542",
    x"2881929B",
    x"28816008",
    x"28812D88",
    x"2880FB1C",
    x"2880C8C4",
    x"2880967F",
    x"2880644E",
    x"28803231",
    x"28800027",
    x"287F9C62",
    x"287F389C",
    x"287ED4FE",
    x"287E7186",
    x"287E0E35",
    x"287DAB0B",
    x"287D4807",
    x"287CE52B",
    x"287C8274",
    x"287C1FE5",
    x"287BBD7B",
    x"287B5B39",
    x"287AF91C",
    x"287A9726",
    x"287A3556",
    x"2879D3AC",
    x"28797229",
    x"287910CB",
    x"2878AF93",
    x"28784E82",
    x"2877ED96",
    x"28778CD0",
    x"28772C30",
    x"2876CBB6",
    x"28766B61",
    x"28760B32",
    x"2875AB28",
    x"28754B44",
    x"2874EB85",
    x"28748BEC",
    x"28742C78",
    x"2873CD29",
    x"28736E00",
    x"28730EFB",
    x"2872B01C",
    x"28725162",
    x"2871F2CC",
    x"2871945C",
    x"28713610",
    x"2870D7EA",
    x"287079E8",
    x"28701C0A",
    x"286FBE52",
    x"286F60BE",
    x"286F034E",
    x"286EA603",
    x"286E48DC",
    x"286DEBDA",
    x"286D8EFC",
    x"286D3242",
    x"286CD5AD",
    x"286C793B",
    x"286C1CEE",
    x"286BC0C5",
    x"286B64C0",
    x"286B08DE",
    x"286AAD21",
    x"286A5187",
    x"2869F611",
    x"28699ABF",
    x"28693F90",
    x"2868E485",
    x"2868899D",
    x"28682ED9",
    x"2867D439",
    x"286779BC",
    x"28671F62",
    x"2866C52B",
    x"28666B18",
    x"28661127",
    x"2865B75A",
    x"28655DB0",
    x"28650429",
    x"2864AAC5",
    x"28645184",
    x"2863F865",
    x"28639F6A",
    x"28634691",
    x"2862EDDA",
    x"28629547",
    x"28623CD6",
    x"2861E487",
    x"28618C5B",
    x"28613452",
    x"2860DC6A",
    x"286084A5",
    x"28602D03",
    x"285FD582",
    x"285F7E24",
    x"285F26E8",
    x"285ECFCD",
    x"285E78D5",
    x"285E21FF",
    x"285DCB4B",
    x"285D74B8",
    x"285D1E47",
    x"285CC7F8",
    x"285C71CB",
    x"285C1BC0",
    x"285BC5D5",
    x"285B700D",
    x"285B1A66",
    x"285AC4E0",
    x"285A6F7C",
    x"285A1A39",
    x"2859C518",
    x"28597017",
    x"28591B38",
    x"2858C67A",
    x"285871DD",
    x"28581D61",
    x"2857C906",
    x"285774CC",
    x"285720B3",
    x"2856CCBA",
    x"285678E3",
    x"2856252C",
    x"2855D196",
    x"28557E20",
    x"28552ACB",
    x"2854D797",
    x"28548483",
    x"2854318F",
    x"2853DEBC",
    x"28538C09",
    x"28533977",
    x"2852E704",
    x"285294B2",
    x"28524280",
    x"2851F06E",
    x"28519E7C",
    x"28514CAA",
    x"2850FAF8",
    x"2850A966",
    x"285057F4",
    x"285006A1",
    x"284FB56F",
    x"284F645C",
    x"284F1368",
    x"284EC294",
    x"284E71E0",
    x"284E214C",
    x"284DD0D6",
    x"284D8080",
    x"284D304A",
    x"284CE033",
    x"284C903B",
    x"284C4062",
    x"284BF0A8",
    x"284BA10E",
    x"284B5192",
    x"284B0236",
    x"284AB2F9",
    x"284A63DA",
    x"284A14DB",
    x"2849C5FA",
    x"28497738",
    x"28492895",
    x"2848DA10",
    x"28488BAA",
    x"28483D63",
    x"2847EF3A",
    x"2847A130",
    x"28475345",
    x"28470577",
    x"2846B7C8",
    x"28466A38",
    x"28461CC5",
    x"2845CF71",
    x"2845823B",
    x"28453523",
    x"2844E82A",
    x"28449B4E",
    x"28444E90",
    x"284401F1",
    x"2843B56F",
    x"2843690B",
    x"28431CC5",
    x"2842D09C",
    x"28428492",
    x"284238A5",
    x"2841ECD5",
    x"2841A124",
    x"28415590",
    x"28410A19",
    x"2840BEC0",
    x"28407384",
    x"28402865",
    x"283FDD64",
    x"283F9280",
    x"283F47BA",
    x"283EFD10",
    x"283EB284",
    x"283E6815",
    x"283E1DC3",
    x"283DD38E",
    x"283D8975",
    x"283D3F7A",
    x"283CF59C",
    x"283CABDA",
    x"283C6236",
    x"283C18AE",
    x"283BCF42",
    x"283B85F4",
    x"283B3CC2",
    x"283AF3AC",
    x"283AAAB3",
    x"283A61D7",
    x"283A1917",
    x"2839D073",
    x"283987EC",
    x"28393F81",
    x"2838F732",
    x"2838AF00",
    x"283866EA",
    x"28381EEF",
    x"2837D711",
    x"28378F4F",
    x"283747A9",
    x"2837001F",
    x"2836B8B1",
    x"2836715F",
    x"28362A29",
    x"2835E30E",
    x"28359C0F",
    x"2835552C",
    x"28350E65",
    x"2834C7B9",
    x"28348129",
    x"28343AB4",
    x"2833F45B",
    x"2833AE1D",
    x"283367FB",
    x"283321F4",
    x"2832DC08",
    x"28329638",
    x"28325083",
    x"28320AE9",
    x"2831C56A",
    x"28318007",
    x"28313ABE",
    x"2830F591",
    x"2830B07E",
    x"28306B87",
    x"283026AA",
    x"282FE1E9",
    x"282F9D42",
    x"282F58B6",
    x"282F1445",
    x"282ECFEE",
    x"282E8BB2",
    x"282E4791",
    x"282E038A",
    x"282DBF9E",
    x"282D7BCC",
    x"282D3815",
    x"282CF479",
    x"282CB0F6",
    x"282C6D8E",
    x"282C2A41",
    x"282BE70D",
    x"282BA3F4",
    x"282B60F5",
    x"282B1E10",
    x"282ADB46",
    x"282A9895",
    x"282A55FF",
    x"282A1382",
    x"2829D11F",
    x"28298ED7",
    x"28294CA8",
    x"28290A93",
    x"2828C897",
    x"282886B6",
    x"282844EE",
    x"28280340",
    x"2827C1AC",
    x"28278031",
    x"28273ECF",
    x"2826FD88",
    x"2826BC59",
    x"28267B44",
    x"28263A49",
    x"2825F967",
    x"2825B89E",
    x"282577EF",
    x"28253758",
    x"2824F6DB",
    x"2824B678",
    x"2824762D",
    x"282435FB",
    x"2823F5E3",
    x"2823B5E3",
    x"282375FD",
    x"2823362F",
    x"2822F67A",
    x"2822B6DE",
    x"2822775B",
    x"282237F1",
    x"2821F8A0",
    x"2821B967",
    x"28217A47",
    x"28213B3F",
    x"2820FC50",
    x"2820BD7A",
    x"28207EBC",
    x"28204017",
    x"2820018A",
    x"281FC316",
    x"281F84BA",
    x"281F4676",
    x"281F084B",
    x"281ECA38",
    x"281E8C3D",
    x"281E4E5A",
    x"281E1090",
    x"281DD2DD",
    x"281D9543",
    x"281D57C1",
    x"281D1A56",
    x"281CDD04",
    x"281C9FCA",
    x"281C62A7",
    x"281C259D",
    x"281BE8AA",
    x"281BABCF",
    x"281B6F0C",
    x"281B3260",
    x"281AF5CC",
    x"281AB950",
    x"281A7CEB",
    x"281A409E",
    x"281A0469",
    x"2819C84B",
    x"28198C44",
    x"28195055",
    x"2819147E",
    x"2818D8BD",
    x"28189D14",
    x"28186183",
    x"28182608",
    x"2817EAA5",
    x"2817AF59",
    x"28177424",
    x"28173906",
    x"2816FDFF",
    x"2816C310",
    x"28168837",
    x"28164D75",
    x"281612CA",
    x"2815D836",
    x"28159DB9",
    x"28156353",
    x"28152904",
    x"2814EECB",
    x"2814B4A9",
    x"28147A9E",
    x"281440A9",
    x"281406CB",
    x"2813CD04",
    x"28139353",
    x"281359B9",
    x"28132035",
    x"2812E6C8",
    x"2812AD71",
    x"28127430",
    x"28123B06",
    x"281201F2",
    x"2811C8F5",
    x"2811900D",
    x"2811573C",
    x"28111E81",
    x"2810E5DC",
    x"2810AD4D",
    x"281074D5",
    x"28103C72",
    x"28100426",
    x"280FCBEF",
    x"280F93CE",
    x"280F5BC3",
    x"280F23CF",
    x"280EEBEF",
    x"280EB426",
    x"280E7C73",
    x"280E44D5",
    x"280E0D4D",
    x"280DD5DB",
    x"280D9E7E",
    x"280D6737",
    x"280D3005",
    x"280CF8E9",
    x"280CC1E3",
    x"280C8AF2",
    x"280C5416",
    x"280C1D50",
    x"280BE69F",
    x"280BB004",
    x"280B797E",
    x"280B430D",
    x"280B0CB1",
    x"280AD66B",
    x"280AA03A",
    x"280A6A1E",
    x"280A3417",
    x"2809FE25",
    x"2809C848",
    x"28099281",
    x"28095CCE",
    x"28092730",
    x"2808F1A7",
    x"2808BC33",
    x"280886D4",
    x"2808518A",
    x"28081C54",
    x"2807E734",
    x"2807B228",
    x"28077D31",
    x"2807484E",
    x"28071380",
    x"2806DEC7",
    x"2806AA22",
    x"28067592",
    x"28064116",
    x"28060CAF",
    x"2805D85C",
    x"2805A41E",
    x"28056FF4",
    x"28053BDE",
    x"280507DD",
    x"2804D3F0",
    x"2804A018",
    x"28046C53",
    x"280438A3",
    x"28040507",
    x"2803D17F",
    x"28039E0B",
    x"28036AAC",
    x"28033760",
    x"28030428",
    x"2802D105",
    x"28029DF5",
    x"28026AF9",
    x"28023811",
    x"2802053D",
    x"2801D27D",
    x"28019FD1",
    x"28016D38",
    x"28013AB4",
    x"28010843",
    x"2800D5E5",
    x"2800A39B",
    x"28007165",
    x"28003F43",
    x"28000D34",
    x"27FFB671",
    x"27FF52A1",
    x"27FEEEF8",
    x"27FE8B77",
    x"27FE281C",
    x"27FDC4E7",
    x"27FD61DA",
    x"27FCFEF3",
    x"27FC9C32",
    x"27FC3999",
    x"27FBD725",
    x"27FB74D9",
    x"27FB12B2",
    x"27FAB0B2",
    x"27FA4ED8",
    x"27F9ED24",
    x"27F98B97",
    x"27F92A2F",
    x"27F8C8EE",
    x"27F867D2",
    x"27F806DD",
    x"27F7A60D",
    x"27F74563",
    x"27F6E4DF",
    x"27F68480",
    x"27F62447",
    x"27F5C434",
    x"27F56446",
    x"27F5047D",
    x"27F4A4DA",
    x"27F4455D",
    x"27F3E604",
    x"27F386D1",
    x"27F327C3",
    x"27F2C8DA",
    x"27F26A16",
    x"27F20B77",
    x"27F1ACFD",
    x"27F14EA8",
    x"27F0F077",
    x"27F0926C",
    x"27F03485",
    x"27EFD6C3",
    x"27EF7925",
    x"27EF1BAC",
    x"27EEBE58",
    x"27EE6127",
    x"27EE041C",
    x"27EDA734",
    x"27ED4A71",
    x"27ECEDD2",
    x"27EC9157",
    x"27EC3500",
    x"27EBD8CE",
    x"27EB7CBF",
    x"27EB20D4",
    x"27EAC50D",
    x"27EA696A",
    x"27EA0DEB",
    x"27E9B28F",
    x"27E95757",
    x"27E8FC43",
    x"27E8A152",
    x"27E84685",
    x"27E7EBDB",
    x"27E79155",
    x"27E736F2",
    x"27E6DCB2",
    x"27E68295",
    x"27E6289C",
    x"27E5CEC6",
    x"27E57512",
    x"27E51B82",
    x"27E4C215",
    x"27E468CA",
    x"27E40FA3",
    x"27E3B69E",
    x"27E35DBC",
    x"27E304FD",
    x"27E2AC60",
    x"27E253E6",
    x"27E1FB8F",
    x"27E1A35A",
    x"27E14B47",
    x"27E0F357",
    x"27E09B89",
    x"27E043DD",
    x"27DFEC54",
    x"27DF94ED",
    x"27DF3DA8",
    x"27DEE685",
    x"27DE8F83",
    x"27DE38A4",
    x"27DDE1E7",
    x"27DD8B4C",
    x"27DD34D2",
    x"27DCDE7B",
    x"27DC8845",
    x"27DC3230",
    x"27DBDC3D",
    x"27DB866C",
    x"27DB30BC",
    x"27DADB2E",
    x"27DA85C1",
    x"27DA3075",
    x"27D9DB4B",
    x"27D98642",
    x"27D9315A",
    x"27D8DC94",
    x"27D887EE",
    x"27D83369",
    x"27D7DF06",
    x"27D78AC3",
    x"27D736A1",
    x"27D6E2A0",
    x"27D68EC0",
    x"27D63B01",
    x"27D5E762",
    x"27D593E4",
    x"27D54087",
    x"27D4ED4A",
    x"27D49A2D",
    x"27D44731",
    x"27D3F456",
    x"27D3A19A",
    x"27D34EFF",
    x"27D2FC85",
    x"27D2AA2A",
    x"27D257F0",
    x"27D205D5",
    x"27D1B3DB",
    x"27D16201",
    x"27D11046",
    x"27D0BEAC",
    x"27D06D31",
    x"27D01BD7",
    x"27CFCA9C",
    x"27CF7980",
    x"27CF2885",
    x"27CED7A9",
    x"27CE86EC",
    x"27CE364F",
    x"27CDE5D2",
    x"27CD9574",
    x"27CD4535",
    x"27CCF516",
    x"27CCA515",
    x"27CC5535",
    x"27CC0573",
    x"27CBB5D0",
    x"27CB664D",
    x"27CB16E8",
    x"27CAC7A3",
    x"27CA787C",
    x"27CA2975",
    x"27C9DA8C",
    x"27C98BC2",
    x"27C93D17",
    x"27C8EE8A",
    x"27C8A01C",
    x"27C851CD",
    x"27C8039D",
    x"27C7B58A",
    x"27C76797",
    x"27C719C1",
    x"27C6CC0B",
    x"27C67E72",
    x"27C630F8",
    x"27C5E39C",
    x"27C5965E",
    x"27C5493E",
    x"27C4FC3D",
    x"27C4AF59",
    x"27C46294",
    x"27C415EC",
    x"27C3C963",
    x"27C37CF7",
    x"27C330A9",
    x"27C2E479",
    x"27C29866",
    x"27C24C72",
    x"27C2009B",
    x"27C1B4E1",
    x"27C16945",
    x"27C11DC7",
    x"27C0D266",
    x"27C08723",
    x"27C03BFC",
    x"27BFF0F4",
    x"27BFA608",
    x"27BF5B3A",
    x"27BF1089",
    x"27BEC5F5",
    x"27BE7B7E",
    x"27BE3125",
    x"27BDE6E8",
    x"27BD9CC8",
    x"27BD52C5",
    x"27BD08DF",
    x"27BCBF16",
    x"27BC756A",
    x"27BC2BDB",
    x"27BBE268",
    x"27BB9912",
    x"27BB4FD8",
    x"27BB06BB",
    x"27BABDBB",
    x"27BA74D7",
    x"27BA2C10",
    x"27B9E365",
    x"27B99AD6",
    x"27B95264",
    x"27B90A0E",
    x"27B8C1D4",
    x"27B879B6",
    x"27B831B5",
    x"27B7E9CF",
    x"27B7A206",
    x"27B75A59",
    x"27B712C7",
    x"27B6CB52",
    x"27B683F9",
    x"27B63CBB",
    x"27B5F599",
    x"27B5AE93",
    x"27B567A9",
    x"27B520DA",
    x"27B4DA27",
    x"27B49390",
    x"27B44D14",
    x"27B406B3",
    x"27B3C06E",
    x"27B37A45",
    x"27B33437",
    x"27B2EE44",
    x"27B2A86D",
    x"27B262B1",
    x"27B21D10",
    x"27B1D78A",
    x"27B1921F",
    x"27B14CD0",
    x"27B1079B",
    x"27B0C282",
    x"27B07D83",
    x"27B038A0",
    x"27AFF3D7",
    x"27AFAF29",
    x"27AF6A96",
    x"27AF261E",
    x"27AEE1C0",
    x"27AE9D7E",
    x"27AE5955",
    x"27AE1548",
    x"27ADD155",
    x"27AD8D7C",
    x"27AD49BE",
    x"27AD061B",
    x"27ACC291",
    x"27AC7F23",
    x"27AC3BCE",
    x"27ABF894",
    x"27ABB574",
    x"27AB726E",
    x"27AB2F82",
    x"27AAECB1",
    x"27AAA9F9",
    x"27AA675C",
    x"27AA24D9",
    x"27A9E26F",
    x"27A9A020",
    x"27A95DEA",
    x"27A91BCE",
    x"27A8D9CC",
    x"27A897E4",
    x"27A85616",
    x"27A81461",
    x"27A7D2C6",
    x"27A79144",
    x"27A74FDC",
    x"27A70E8E",
    x"27A6CD59",
    x"27A68C3D",
    x"27A64B3B",
    x"27A60A53",
    x"27A5C983",
    x"27A588CD",
    x"27A54830",
    x"27A507AD",
    x"27A4C742",
    x"27A486F1",
    x"27A446B9",
    x"27A4069A",
    x"27A3C694",
    x"27A386A7",
    x"27A346D3",
    x"27A30717",
    x"27A2C775",
    x"27A287EC",
    x"27A2487B",
    x"27A20923",
    x"27A1C9E4",
    x"27A18ABD",
    x"27A14BAF",
    x"27A10CBA",
    x"27A0CDDD",
    x"27A08F19",
    x"27A0506E",
    x"27A011DA",
    x"279FD360",
    x"279F94FD",
    x"279F56B3",
    x"279F1881",
    x"279EDA68",
    x"279E9C67",
    x"279E5E7E",
    x"279E20AD",
    x"279DE2F4",
    x"279DA554",
    x"279D67CB",
    x"279D2A5B",
    x"279CED02",
    x"279CAFC1",
    x"279C7299",
    x"279C3588",
    x"279BF88F",
    x"279BBBAE",
    x"279B7EE4",
    x"279B4232",
    x"279B0598",
    x"279AC916",
    x"279A8CAB",
    x"279A5058",
    x"279A141D",
    x"2799D7F8",
    x"27999BEC",
    x"27995FF7",
    x"27992419",
    x"2798E852",
    x"2798ACA3",
    x"2798710C",
    x"2798358B",
    x"2797FA22",
    x"2797BED0",
    x"27978395",
    x"27974871",
    x"27970D64",
    x"2796D26E",
    x"27969790",
    x"27965CC8",
    x"27962217",
    x"2795E77D",
    x"2795ACFA",
    x"2795728E",
    x"27953839",
    x"2794FDFA",
    x"2794C3D2",
    x"279489C1",
    x"27944FC7",
    x"279415E3",
    x"2793DC16",
    x"2793A25F",
    x"279368BF",
    x"27932F35",
    x"2792F5C2",
    x"2792BC65",
    x"2792831F",
    x"279249EF",
    x"279210D5",
    x"2791D7D1",
    x"27919EE4",
    x"2791660D",
    x"27912D4C",
    x"2790F4A2",
    x"2790BC0D",
    x"2790838F",
    x"27904B27",
    x"279012D4",
    x"278FDA98",
    x"278FA271",
    x"278F6A61",
    x"278F3266",
    x"278EFA82",
    x"278EC2B3",
    x"278E8AF9",
    x"278E5356",
    x"278E1BC8",
    x"278DE450",
    x"278DACEE",
    x"278D75A1",
    x"278D3E6A",
    x"278D0748",
    x"278CD03C",
    x"278C9946",
    x"278C6265",
    x"278C2B99",
    x"278BF4E2",
    x"278BBE41",
    x"278B87B6",
    x"278B513F",
    x"278B1ADE",
    x"278AE492",
    x"278AAE5C",
    x"278A783A",
    x"278A422E",
    x"278A0C36",
    x"2789D654",
    x"2789A087",
    x"27896ACF",
    x"2789352C",
    x"2788FF9D",
    x"2788CA24",
    x"278894BF",
    x"27885F70",
    x"27882A35",
    x"2787F50F",
    x"2787BFFD",
    x"27878B01",
    x"27875619",
    x"27872145",
    x"2786EC87",
    x"2786B7DD",
    x"27868347",
    x"27864EC6",
    x"27861A5A",
    x"2785E601",
    x"2785B1BE",
    x"27857D8F",
    x"27854974",
    x"2785156D",
    x"2784E17B",
    x"2784AD9D",
    x"278479D3",
    x"2784461E",
    x"2784127D",
    x"2783DEEF",
    x"2783AB76",
    x"27837811",
    x"278344C1",
    x"27831184",
    x"2782DE5B",
    x"2782AB46",
    x"27827845",
    x"27824558",
    x"2782127F",
    x"2781DFBA",
    x"2781AD08",
    x"27817A6A",
    x"278147E0",
    x"2781156A",
    x"2780E308",
    x"2780B0B9",
    x"27807E7E",
    x"27804C56",
    x"27801A42",
    x"277FD083",
    x"277F6CA9",
    x"277F08F6",
    x"277EA56A",
    x"277E4205",
    x"277DDEC6",
    x"277D7BAF",
    x"277D18BE",
    x"277CB5F3",
    x"277C534F",
    x"277BF0D2",
    x"277B8E7B",
    x"277B2C4B",
    x"277ACA41",
    x"277A685D",
    x"277A069F",
    x"2779A508",
    x"27794396",
    x"2778E24B",
    x"27788125",
    x"27782026",
    x"2777BF4C",
    x"27775E98",
    x"2776FE0A",
    x"27769DA2",
    x"27763D5F",
    x"2775DD42",
    x"27757D4A",
    x"27751D78",
    x"2774BDCB",
    x"27745E44",
    x"2773FEE2",
    x"27739FA5",
    x"2773408D",
    x"2772E19A",
    x"277282CD",
    x"27722424",
    x"2771C5A0",
    x"27716742",
    x"27710908",
    x"2770AAF2",
    x"27704D02",
    x"276FEF36",
    x"276F918F",
    x"276F340D",
    x"276ED6AE",
    x"276E7975",
    x"276E1C60",
    x"276DBF6F",
    x"276D62A2",
    x"276D05FA",
    x"276CA975",
    x"276C4D15",
    x"276BF0D9",
    x"276B94C1",
    x"276B38CD",
    x"276ADCFD",
    x"276A8150",
    x"276A25C8",
    x"2769CA63",
    x"27696F21",
    x"27691404",
    x"2768B90A",
    x"27685E33",
    x"27680380",
    x"2767A8F0",
    x"27674E84",
    x"2766F43B",
    x"27669A15",
    x"27664013",
    x"2765E633",
    x"27658C77",
    x"276532DD",
    x"2764D967",
    x"27648014",
    x"276426E3",
    x"2763CDD5",
    x"276374EA",
    x"27631C22",
    x"2762C37C",
    x"27626AF9",
    x"27621299",
    x"2761BA5B",
    x"2761623F",
    x"27610A46",
    x"2760B26F",
    x"27605ABA",
    x"27600328",
    x"275FABB8",
    x"275F546A",
    x"275EFD3E",
    x"275EA634",
    x"275E4F4C",
    x"275DF886",
    x"275DA1E2",
    x"275D4B60",
    x"275CF4FF",
    x"275C9EC0",
    x"275C48A3",
    x"275BF2A7",
    x"275B9CCD",
    x"275B4715",
    x"275AF17E",
    x"275A9C08",
    x"275A46B4",
    x"2759F181",
    x"27599C6F",
    x"2759477F",
    x"2758F2AF",
    x"27589E01",
    x"27584974",
    x"2757F508",
    x"2757A0BC",
    x"27574C92",
    x"2756F889",
    x"2756A4A0",
    x"275650D8",
    x"2755FD31",
    x"2755A9AA",
    x"27555644",
    x"275502FF",
    x"2754AFDA",
    x"27545CD5",
    x"275409F1",
    x"2753B72E",
    x"2753648A",
    x"27531207",
    x"2752BFA4",
    x"27526D61",
    x"27521B3F",
    x"2751C93C",
    x"27517759",
    x"27512597",
    x"2750D3F4",
    x"27508271",
    x"2750310E",
    x"274FDFCB",
    x"274F8EA7",
    x"274F3DA3",
    x"274EECBF",
    x"274E9BFA",
    x"274E4B55",
    x"274DFACF",
    x"274DAA69",
    x"274D5A22",
    x"274D09FB",
    x"274CB9F2",
    x"274C6A09",
    x"274C1A40",
    x"274BCA95",
    x"274B7B09",
    x"274B2B9D",
    x"274ADC4F",
    x"274A8D21",
    x"274A3E11",
    x"2749EF20",
    x"2749A04E",
    x"2749519B",
    x"27490306",
    x"2748B491",
    x"27486639",
    x"27481801",
    x"2747C9E7",
    x"27477BEB",
    x"27472E0E",
    x"2746E04F",
    x"274692AE",
    x"2746452C",
    x"2745F7C8",
    x"2745AA83",
    x"27455D5B",
    x"27451052",
    x"2744C366",
    x"27447699",
    x"274429EA",
    x"2743DD58",
    x"274390E5",
    x"2743448F",
    x"2742F857",
    x"2742AC3D",
    x"27426041",
    x"27421462",
    x"2741C8A1",
    x"27417CFD",
    x"27413177",
    x"2740E60E",
    x"27409AC3",
    x"27404F96",
    x"27400485",
    x"273FB992",
    x"273F6EBC",
    x"273F2403",
    x"273ED968",
    x"273E8EEA",
    x"273E4488",
    x"273DFA44",
    x"273DB01D",
    x"273D6612",
    x"273D1C25",
    x"273CD254",
    x"273C88A1",
    x"273C3F0A",
    x"273BF58F",
    x"273BAC32",
    x"273B62F1",
    x"273B19CD",
    x"273AD0C5",
    x"273A87D9",
    x"273A3F0B",
    x"2739F658",
    x"2739ADC2",
    x"27396548",
    x"27391CEB",
    x"2738D4AA",
    x"27388C85",
    x"2738447C",
    x"2737FC8F",
    x"2737B4BF",
    x"27376D0A",
    x"27372571",
    x"2736DDF5",
    x"27369694",
    x"27364F4F",
    x"27360826",
    x"2735C119",
    x"27357A27",
    x"27353351",
    x"2734EC97",
    x"2734A5F8",
    x"27345F75",
    x"2734190E",
    x"2733D2C2",
    x"27338C91",
    x"2733467C",
    x"27330082",
    x"2732BAA4",
    x"273274E0",
    x"27322F38",
    x"2731E9AB",
    x"2731A43A",
    x"27315EE3",
    x"273119A8",
    x"2730D487",
    x"27308F81",
    x"27304A97",
    x"273005C7",
    x"272FC112",
    x"272F7C78",
    x"272F37F9",
    x"272EF395",
    x"272EAF4B",
    x"272E6B1C",
    x"272E2707",
    x"272DE30D",
    x"272D9F2E",
    x"272D5B69",
    x"272D17BE",
    x"272CD42E",
    x"272C90B8",
    x"272C4D5D",
    x"272C0A1C",
    x"272BC6F5",
    x"272B83E9",
    x"272B40F6",
    x"272AFE1E",
    x"272ABB60",
    x"272A78BB",
    x"272A3631",
    x"2729F3C1",
    x"2729B16B",
    x"27296F2E",
    x"27292D0C",
    x"2728EB03",
    x"2728A914",
    x"2728673F",
    x"27282584",
    x"2727E3E2",
    x"2727A25A",
    x"272760EB",
    x"27271F96",
    x"2726DE5A",
    x"27269D38",
    x"27265C2F",
    x"27261B40",
    x"2725DA6A",
    x"272599AD",
    x"2725590A",
    x"27251880",
    x"2724D80F",
    x"272497B7",
    x"27245778",
    x"27241753",
    x"2723D746",
    x"27239753",
    x"27235778",
    x"272317B6",
    x"2722D80D",
    x"2722987D",
    x"27225906",
    x"272219A8",
    x"2721DA62",
    x"27219B35",
    x"27215C21",
    x"27211D25",
    x"2720DE42",
    x"27209F78",
    x"272060C6",
    x"2720222C",
    x"271FE3AB",
    x"271FA542",
    x"271F66F2",
    x"271F28BA",
    x"271EEA9A",
    x"271EAC92",
    x"271E6EA3",
    x"271E30CC",
    x"271DF30D",
    x"271DB566",
    x"271D77D7",
    x"271D3A60",
    x"271CFD02",
    x"271CBFBB",
    x"271C828C",
    x"271C4575",
    x"271C0875",
    x"271BCB8E",
    x"271B8EBE",
    x"271B5207",
    x"271B1566",
    x"271AD8DE",
    x"271A9C6D",
    x"271A6014",
    x"271A23D2",
    x"2719E7A8",
    x"2719AB95",
    x"27196F9A",
    x"271933B6",
    x"2718F7E9",
    x"2718BC34",
    x"27188096",
    x"2718450F",
    x"271809A0",
    x"2717CE48",
    x"27179307",
    x"271757DD",
    x"27171CCA",
    x"2716E1CF",
    x"2716A6EA",
    x"27166C1C",
    x"27163165",
    x"2715F6C6",
    x"2715BC3D",
    x"271581CA",
    x"2715476F",
    x"27150D2B",
    x"2714D2FD",
    x"271498E6",
    x"27145EE5",
    x"271424FC",
    x"2713EB29",
    x"2713B16C",
    x"271377C6",
    x"27133E36",
    x"271304BD",
    x"2712CB5B",
    x"2712920E",
    x"271258D9",
    x"27121FB9",
    x"2711E6B0",
    x"2711ADBD",
    x"271174E0",
    x"27113C19",
    x"27110369",
    x"2710CACF",
    x"2710924B",
    x"271059DC",
    x"27102184",
    x"270FE942",
    x"270FB116",
    x"270F7900",
    x"270F4100",
    x"270F0915",
    x"270ED140",
    x"270E9982",
    x"270E61D9",
    x"270E2A45",
    x"270DF2C7",
    x"270DBB5F",
    x"270D840D",
    x"270D4CD0",
    x"270D15A9",
    x"270CDE97",
    x"270CA79B",
    x"270C70B4",
    x"270C39E3",
    x"270C0327",
    x"270BCC81",
    x"270B95EF",
    x"270B5F73",
    x"270B290D",
    x"270AF2BB",
    x"270ABC7F",
    x"270A8658",
    x"270A5046",
    x"270A1A49",
    x"2709E462",
    x"2709AE8F",
    x"270978D1",
    x"27094329",
    x"27090D95",
    x"2708D816",
    x"2708A2AC",
    x"27086D57",
    x"27083817",
    x"270802EB",
    x"2707CDD4",
    x"270798D2",
    x"270763E5",
    x"27072F0C",
    x"2706FA48",
    x"2706C599",
    x"270690FE",
    x"27065C77",
    x"27062805",
    x"2705F3A8",
    x"2705BF5F",
    x"27058B2B",
    x"2705570A",
    x"270522FE",
    x"2704EF07",
    x"2704BB24",
    x"27048755",
    x"2704539A",
    x"27041FF3",
    x"2703EC61",
    x"2703B8E3",
    x"27038579",
    x"27035222",
    x"27031EE0",
    x"2702EBB2",
    x"2702B898",
    x"27028592",
    x"270252A0",
    x"27021FC2",
    x"2701ECF7",
    x"2701BA40",
    x"2701879E",
    x"2701550E",
    x"27012293",
    x"2700F02B",
    x"2700BDD7",
    x"27008B97",
    x"2700596A",
    x"27002751",
    x"26FFEA97",
    x"26FF86B3",
    x"26FF22F6",
    x"26FEBF60",
    x"26FE5BF1",
    x"26FDF8A8",
    x"26FD9586",
    x"26FD328B",
    x"26FCCFB7",
    x"26FC6D09",
    x"26FC0A82",
    x"26FBA821",
    x"26FB45E6",
    x"26FAE3D2",
    x"26FA81E4",
    x"26FA201D",
    x"26F9BE7B",
    x"26F95D00",
    x"26F8FBAA",
    x"26F89A7B",
    x"26F83972",
    x"26F7D88E",
    x"26F777D0",
    x"26F71739",
    x"26F6B6C6",
    x"26F6567A",
    x"26F5F653",
    x"26F59651",
    x"26F53675",
    x"26F4D6BF",
    x"26F4772E",
    x"26F417C2",
    x"26F3B87B",
    x"26F35959",
    x"26F2FA5D",
    x"26F29B86",
    x"26F23CD4",
    x"26F1DE46",
    x"26F17FDE",
    x"26F1219A",
    x"26F0C37C",
    x"26F06582",
    x"26F007AC",
    x"26EFA9FC",
    x"26EF4C70",
    x"26EEEF08",
    x"26EE91C5",
    x"26EE34A6",
    x"26EDD7AC",
    x"26ED7AD5",
    x"26ED1E24",
    x"26ECC196",
    x"26EC652C",
    x"26EC08E7",
    x"26EBACC5",
    x"26EB50C8",
    x"26EAF4EE",
    x"26EA9938",
    x"26EA3DA7",
    x"26E9E238",
    x"26E986EE",
    x"26E92BC7",
    x"26E8D0C4",
    x"26E875E4",
    x"26E81B27",
    x"26E7C08F",
    x"26E76619",
    x"26E70BC7",
    x"26E6B198",
    x"26E6578C",
    x"26E5FDA3",
    x"26E5A3DE",
    x"26E54A3B",
    x"26E4F0BC",
    x"26E4975F",
    x"26E43E26",
    x"26E3E50F",
    x"26E38C1B",
    x"26E33349",
    x"26E2DA9A",
    x"26E2820E",
    x"26E229A5",
    x"26E1D15E",
    x"26E17939",
    x"26E12137",
    x"26E0C957",
    x"26E0719A",
    x"26E019FF",
    x"26DFC285",
    x"26DF6B2F",
    x"26DF13FA",
    x"26DEBCE7",
    x"26DE65F6",
    x"26DE0F27",
    x"26DDB87A",
    x"26DD61EF",
    x"26DD0B86",
    x"26DCB53E",
    x"26DC5F18",
    x"26DC0914",
    x"26DBB331",
    x"26DB5D70",
    x"26DB07D0",
    x"26DAB252",
    x"26DA5CF5",
    x"26DA07B9",
    x"26D9B29F",
    x"26D95DA5",
    x"26D908CD",
    x"26D8B417",
    x"26D85F81",
    x"26D80B0C",
    x"26D7B6B8",
    x"26D76285",
    x"26D70E73",
    x"26D6BA82",
    x"26D666B1",
    x"26D61302",
    x"26D5BF73",
    x"26D56C04",
    x"26D518B6",
    x"26D4C589",
    x"26D4727C",
    x"26D41F8F",
    x"26D3CCC3",
    x"26D37A17",
    x"26D3278C",
    x"26D2D520",
    x"26D282D5",
    x"26D230AA",
    x"26D1DE9F",
    x"26D18CB4",
    x"26D13AE9",
    x"26D0E93E",
    x"26D097B3",
    x"26D04648",
    x"26CFF4FC",
    x"26CFA3D0",
    x"26CF52C4",
    x"26CF01D8",
    x"26CEB10B",
    x"26CE605D",
    x"26CE0FCF",
    x"26CDBF61",
    x"26CD6F12",
    x"26CD1EE2",
    x"26CCCED2",
    x"26CC7EE0",
    x"26CC2F0E",
    x"26CBDF5C",
    x"26CB8FC8",
    x"26CB4053",
    x"26CAF0FE",
    x"26CAA1C7",
    x"26CA52AF",
    x"26CA03B6",
    x"26C9B4DC",
    x"26C96621",
    x"26C91785",
    x"26C8C907",
    x"26C87AA7",
    x"26C82C67",
    x"26C7DE45",
    x"26C79041",
    x"26C7425C",
    x"26C6F495",
    x"26C6A6ED",
    x"26C65963",
    x"26C60BF7",
    x"26C5BEAA",
    x"26C5717A",
    x"26C52469",
    x"26C4D776",
    x"26C48AA1",
    x"26C43DE9",
    x"26C3F150",
    x"26C3A4D5",
    x"26C35877",
    x"26C30C38",
    x"26C2C016",
    x"26C27412",
    x"26C2282B",
    x"26C1DC62",
    x"26C190B7",
    x"26C14529",
    x"26C0F9B9",
    x"26C0AE66",
    x"26C06331",
    x"26C01819",
    x"26BFCD1E",
    x"26BF8240",
    x"26BF3780",
    x"26BEECDD",
    x"26BEA257",
    x"26BE57EE",
    x"26BE0DA2",
    x"26BDC373",
    x"26BD7962",
    x"26BD2F6D",
    x"26BCE594",
    x"26BC9BD9",
    x"26BC523B",
    x"26BC08B9",
    x"26BBBF54",
    x"26BB760B",
    x"26BB2CE0",
    x"26BAE3D0",
    x"26BA9ADE",
    x"26BA5207",
    x"26BA094E",
    x"26B9C0B0",
    x"26B9782F",
    x"26B92FCA",
    x"26B8E782",
    x"26B89F55",
    x"26B85745",
    x"26B80F51",
    x"26B7C779",
    x"26B77FBD",
    x"26B7381D",
    x"26B6F099",
    x"26B6A931",
    x"26B661E5",
    x"26B61AB5",
    x"26B5D3A0",
    x"26B58CA8",
    x"26B545CA",
    x"26B4FF09",
    x"26B4B863",
    x"26B471D9",
    x"26B42B6A",
    x"26B3E517",
    x"26B39EDF",
    x"26B358C3",
    x"26B312C2",
    x"26B2CCDC",
    x"26B28712",
    x"26B24163",
    x"26B1FBCF",
    x"26B1B656",
    x"26B170F8",
    x"26B12BB6",
    x"26B0E68E",
    x"26B0A181",
    x"26B05C90",
    x"26B017B9",
    x"26AFD2FD",
    x"26AF8E5C",
    x"26AF49D6",
    x"26AF056B",
    x"26AEC11A",
    x"26AE7CE4",
    x"26AE38C8",
    x"26ADF4C7",
    x"26ADB0E1",
    x"26AD6D15",
    x"26AD2964",
    x"26ACE5CD",
    x"26ACA250",
    x"26AC5EEE",
    x"26AC1BA6",
    x"26ABD878",
    x"26AB9565",
    x"26AB526C",
    x"26AB0F8D",
    x"26AACCC7",
    x"26AA8A1D",
    x"26AA478C",
    x"26AA0515",
    x"26A9C2B8",
    x"26A98074",
    x"26A93E4B",
    x"26A8FC3C",
    x"26A8BA46",
    x"26A8786A",
    x"26A836A8",
    x"26A7F500",
    x"26A7B371",
    x"26A771FB",
    x"26A730A0",
    x"26A6EF5D",
    x"26A6AE35",
    x"26A66D25",
    x"26A62C2F",
    x"26A5EB53",
    x"26A5AA8F",
    x"26A569E5",
    x"26A52955",
    x"26A4E8DD",
    x"26A4A87F",
    x"26A46839",
    x"26A4280D",
    x"26A3E7FA",
    x"26A3A800",
    x"26A3681F",
    x"26A32857",
    x"26A2E8A7",
    x"26A2A911",
    x"26A26993",
    x"26A22A2E",
    x"26A1EAE2",
    x"26A1ABAF",
    x"26A16C94",
    x"26A12D92",
    x"26A0EEA9",
    x"26A0AFD8",
    x"26A0711F",
    x"26A0327F",
    x"269FF3F8",
    x"269FB589",
    x"269F7732",
    x"269F38F3",
    x"269EFACD",
    x"269EBCC0",
    x"269E7ECA",
    x"269E40EC",
    x"269E0327",
    x"269DC57A",
    x"269D87E5",
    x"269D4A68",
    x"269D0D03",
    x"269CCFB6",
    x"269C9280",
    x"269C5563",
    x"269C185E",
    x"269BDB70",
    x"269B9E9A",
    x"269B61DC",
    x"269B2536",
    x"269AE8A7",
    x"269AAC30",
    x"269A6FD1",
    x"269A3389",
    x"2699F758",
    x"2699BB3F",
    x"26997F3E",
    x"26994354",
    x"26990781",
    x"2698CBC6",
    x"26989022",
    x"26985496",
    x"26981920",
    x"2697DDC2",
    x"2697A27B",
    x"2697674B",
    x"26972C32",
    x"2696F130",
    x"2696B646",
    x"26967B72",
    x"269640B5",
    x"2696060F",
    x"2695CB80",
    x"26959108",
    x"269556A7",
    x"26951C5D",
    x"2694E229",
    x"2694A80C",
    x"26946E06",
    x"26943416",
    x"2693FA3D",
    x"2693C07B",
    x"269386CF",
    x"26934D39",
    x"269313BA",
    x"2692DA52",
    x"2692A100",
    x"269267C4",
    x"26922E9F",
    x"2691F590",
    x"2691BC97",
    x"269183B4",
    x"26914AE8",
    x"26911232",
    x"2690D992",
    x"2690A108",
    x"26906894",
    x"26903036",
    x"268FF7EE",
    x"268FBFBC",
    x"268F87A0",
    x"268F4F9A",
    x"268F17AA",
    x"268EDFD0",
    x"268EA80B",
    x"268E705D",
    x"268E38C3",
    x"268E0140",
    x"268DC9D2",
    x"268D927A",
    x"268D5B38",
    x"268D240B",
    x"268CECF4",
    x"268CB5F2",
    x"268C7F06",
    x"268C482F",
    x"268C116D",
    x"268BDAC1",
    x"268BA42A",
    x"268B6DA9",
    x"268B373D",
    x"268B00E6",
    x"268ACAA4",
    x"268A9477",
    x"268A5E60",
    x"268A285E",
    x"2689F270",
    x"2689BC98",
    x"268986D5",
    x"26895127",
    x"26891B8E",
    x"2688E609",
    x"2688B09A",
    x"26887B3F",
    x"268845FA",
    x"268810C9",
    x"2687DBAD",
    x"2687A6A5",
    x"268771B2",
    x"26873CD4",
    x"2687080B",
    x"2686D356",
    x"26869EB6",
    x"26866A2A",
    x"268635B3",
    x"26860150",
    x"2685CD02",
    x"268598C8",
    x"268564A2",
    x"26853091",
    x"2684FC94",
    x"2684C8AC",
    x"268494D8",
    x"26846118",
    x"26842D6C",
    x"2683F9D4",
    x"2683C651",
    x"268392E1",
    x"26835F86",
    x"26832C3F",
    x"2682F90B",
    x"2682C5EC",
    x"268292E1",
    x"26825FE9",
    x"26822D06",
    x"2681FA36",
    x"2681C77A",
    x"268194D2",
    x"2681623E",
    x"26812FBD",
    x"2680FD51",
    x"2680CAF7",
    x"268098B2",
    x"26806680",
    x"26803462",
    x"26800257",
    x"267FA0C0",
    x"267F3CF9",
    x"267ED958",
    x"267E75DF",
    x"267E128C",
    x"267DAF61",
    x"267D4C5B",
    x"267CE97D",
    x"267C86C5",
    x"267C2434",
    x"267BC1C9",
    x"267B5F84",
    x"267AFD66",
    x"267A9B6E",
    x"267A399D",
    x"2679D7F1",
    x"2679766C",
    x"2679150D",
    x"2678B3D3",
    x"267852C0",
    x"2677F1D3",
    x"2677910B",
    x"26773069",
    x"2676CFED",
    x"26766F97",
    x"26760F66",
    x"2675AF5B",
    x"26754F75",
    x"2674EFB5",
    x"2674901A",
    x"267430A4",
    x"2673D154",
    x"26737229",
    x"26731323",
    x"2672B442",
    x"26725586",
    x"2671F6EF",
    x"2671987D",
    x"26713A30",
    x"2670DC07",
    x"26707E04",
    x"26702025",
    x"266FC26B",
    x"266F64D5",
    x"266F0764",
    x"266EAA17",
    x"266E4CEF",
    x"266DEFEB",
    x"266D930B",
    x"266D3650",
    x"266CD9B9",
    x"266C7D46",
    x"266C20F7",
    x"266BC4CC",
    x"266B68C5",
    x"266B0CE2",
    x"266AB123",
    x"266A5588",
    x"2669FA10",
    x"26699EBD",
    x"2669438C",
    x"2668E880",
    x"26688D97",
    x"266832D1",
    x"2667D82F",
    x"26677DB0",
    x"26672355",
    x"2666C91D",
    x"26666F08",
    x"26661516",
    x"2665BB47",
    x"2665619C",
    x"26650813",
    x"2664AEAD",
    x"2664556A",
    x"2663FC4A",
    x"2663A34D",
    x"26634A73",
    x"2662F1BB",
    x"26629926",
    x"266240B3",
    x"2661E863",
    x"26619036",
    x"2661382B",
    x"2660E042",
    x"2660887C",
    x"266030D7",
    x"265FD955",
    x"265F81F6",
    x"265F2AB8",
    x"265ED39C",
    x"265E7CA2",
    x"265E25CB",
    x"265DCF15",
    x"265D7881",
    x"265D220F",
    x"265CCBBE",
    x"265C7590",
    x"265C1F82",
    x"265BC997",
    x"265B73CD",
    x"265B1E24",
    x"265AC89D",
    x"265A7338",
    x"265A1DF3",
    x"2659C8D0",
    x"265973CE",
    x"26591EEE",
    x"2658CA2E",
    x"26587590",
    x"26582112",
    x"2657CCB6",
    x"2657787A",
    x"26572460",
    x"2656D066",
    x"26567C8D",
    x"265628D5",
    x"2655D53D",
    x"265581C6",
    x"26552E70",
    x"2654DB3A",
    x"26548824",
    x"2654352F",
    x"2653E25B",
    x"26538FA7",
    x"26533D13",
    x"2652EA9F",
    x"2652984B",
    x"26524618",
    x"2651F404",
    x"2651A211",
    x"2651503E",
    x"2650FE8A",
    x"2650ACF7",
    x"26505B83",
    x"26500A2F",
    x"264FB8FB",
    x"264F67E7",
    x"264F16F2",
    x"264EC61D",
    x"264E7567",
    x"264E24D1",
    x"264DD45B",
    x"264D8403",
    x"264D33CB",
    x"264CE3B3",
    x"264C93BA",
    x"264C43DF",
    x"264BF424",
    x"264BA489",
    x"264B550C",
    x"264B05AE",
    x"264AB66F",
    x"264A6750",
    x"264A184F",
    x"2649C96D",
    x"26497AA9",
    x"26492C05",
    x"2648DD7F",
    x"26488F18",
    x"264840CF",
    x"2647F2A5",
    x"2647A49A",
    x"264756AD",
    x"264708DE",
    x"2646BB2E",
    x"26466D9C",
    x"26462028",
    x"2645D2D2",
    x"2645859B",
    x"26453882",
    x"2644EB87",
    x"26449EAA",
    x"264451EB",
    x"2644054A",
    x"2643B8C7",
    x"26436C62",
    x"2643201A",
    x"2642D3F1",
    x"264287E5",
    x"26423BF6",
    x"2641F026",
    x"2641A473",
    x"264158DD",
    x"26410D65",
    x"2640C20B",
    x"264076CE",
    x"26402BAE",
    x"263FE0AC",
    x"263F95C6",
    x"263F4AFF",
    x"263F0054",
    x"263EB5C6",
    x"263E6B56",
    x"263E2102",
    x"263DD6CC",
    x"263D8CB3",
    x"263D42B6",
    x"263CF8D6",
    x"263CAF14",
    x"263C656E",
    x"263C1BE4",
    x"263BD278",
    x"263B8928",
    x"263B3FF5",
    x"263AF6DE",
    x"263AADE4",
    x"263A6506",
    x"263A1C45",
    x"2639D3A0",
    x"26398B18",
    x"263942AB",
    x"2638FA5B",
    x"2638B228",
    x"26386A10",
    x"26382215",
    x"2637DA36",
    x"26379272",
    x"26374ACB",
    x"26370340",
    x"2636BBD1",
    x"2636747D",
    x"26362D46",
    x"2635E62A",
    x"26359F2A",
    x"26355845",
    x"2635117D",
    x"2634CAD0",
    x"2634843E",
    x"26343DC8",
    x"2633F76E",
    x"2633B12F",
    x"26336B0C",
    x"26332503",
    x"2632DF17",
    x"26329945",
    x"2632538F",
    x"26320DF4",
    x"2631C874",
    x"2631830F",
    x"26313DC6",
    x"2630F897",
    x"2630B383",
    x"26306E8B",
    x"263029AD",
    x"262FE4EA",
    x"262FA042",
    x"262F5BB5",
    x"262F1742",
    x"262ED2EB",
    x"262E8EAE",
    x"262E4A8B",
    x"262E0683",
    x"262DC296",
    x"262D7EC3",
    x"262D3B0B",
    x"262CF76D",
    x"262CB3EA",
    x"262C7081",
    x"262C2D32",
    x"262BE9FD",
    x"262BA6E3",
    x"262B63E3",
    x"262B20FD",
    x"262ADE31",
    x"262A9B7F",
    x"262A58E8",
    x"262A166A",
    x"2629D406",
    x"262991BC",
    x"26294F8C",
    x"26290D76",
    x"2628CB7A",
    x"26288997",
    x"262847CE",
    x"2628061F",
    x"2627C489",
    x"2627830D",
    x"262741AB",
    x"26270062",
    x"2626BF33",
    x"26267E1D",
    x"26263D20",
    x"2625FC3D",
    x"2625BB73",
    x"26257AC3",
    x"26253A2B",
    x"2624F9AD",
    x"2624B948",
    x"262478FC",
    x"262438CA",
    x"2623F8B0",
    x"2623B8AF",
    x"262378C8",
    x"262338F9",
    x"2622F943",
    x"2622B9A6",
    x"26227A22",
    x"26223AB7",
    x"2621FB64",
    x"2621BC2A",
    x"26217D09",
    x"26213E01",
    x"2620FF11",
    x"2620C039",
    x"2620817B",
    x"262042D4",
    x"26200446",
    x"261FC5D1",
    x"261F8774",
    x"261F492F",
    x"261F0B03",
    x"261ECCEE",
    x"261E8EF2",
    x"261E510F",
    x"261E1343",
    x"261DD590",
    x"261D97F4",
    x"261D5A71",
    x"261D1D06",
    x"261CDFB2",
    x"261CA277",
    x"261C6553",
    x"261C2848",
    x"261BEB54",
    x"261BAE78",
    x"261B71B4",
    x"261B3507",
    x"261AF872",
    x"261ABBF5",
    x"261A7F8F",
    x"261A4341",
    x"261A070B",
    x"2619CAEC",
    x"26198EE4",
    x"261952F4",
    x"2619171B",
    x"2618DB5A",
    x"26189FB0",
    x"2618641D",
    x"261828A2",
    x"2617ED3D",
    x"2617B1F0",
    x"261776BA",
    x"26173B9C",
    x"26170094",
    x"2616C5A3",
    x"26168AC9",
    x"26165007",
    x"2616155B",
    x"2615DAC6",
    x"2615A048",
    x"261565E1",
    x"26152B90",
    x"2614F157",
    x"2614B734",
    x"26147D28",
    x"26144332",
    x"26140953",
    x"2613CF8B",
    x"261395D9",
    x"26135C3E",
    x"261322B9",
    x"2612E94A",
    x"2612AFF3",
    x"261276B1",
    x"26123D86",
    x"26120471",
    x"2611CB72",
    x"2611928A",
    x"261159B8",
    x"261120FC",
    x"2610E856",
    x"2610AFC6",
    x"2610774D",
    x"26103EE9",
    x"2610069C",
    x"260FCE64",
    x"260F9642",
    x"260F5E37",
    x"260F2641",
    x"260EEE61",
    x"260EB696",
    x"260E7EE2",
    x"260E4743",
    x"260E0FBA",
    x"260DD847",
    x"260DA0E9",
    x"260D69A1",
    x"260D326F",
    x"260CFB52",
    x"260CC44A",
    x"260C8D59",
    x"260C567C",
    x"260C1FB5",
    x"260BE903",
    x"260BB267",
    x"260B7BE0",
    x"260B456E",
    x"260B0F12",
    x"260AD8CA",
    x"260AA298",
    x"260A6C7B",
    x"260A3673",
    x"260A0081",
    x"2609CAA3",
    x"260994DA",
    x"26095F27",
    x"26092988",
    x"2608F3FE",
    x"2608BE89",
    x"26088929",
    x"260853DE",
    x"26081EA8",
    x"2607E986",
    x"2607B479",
    x"26077F81",
    x"26074A9E",
    x"260715CF",
    x"2606E115",
    x"2606AC6F",
    x"260677DE",
    x"26064361",
    x"26060EF9",
    x"2605DAA6",
    x"2605A667",
    x"2605723C",
    x"26053E25",
    x"26050A23",
    x"2604D635",
    x"2604A25C",
    x"26046E97",
    x"26043AE5",
    x"26040748",
    x"2603D3C0",
    x"2603A04B",
    x"26036CEA",
    x"2603399E",
    x"26030665",
    x"2602D341",
    x"2602A030",
    x"26026D34",
    x"26023A4B",
    x"26020776",
    x"2601D4B5",
    x"2601A208",
    x"26016F6F",
    x"26013CE9",
    x"26010A77",
    x"2600D819",
    x"2600A5CE",
    x"26007397",
    x"26004174",
    x"26000F64",
    x"25FFBAD0",
    x"25FF56FE",
    x"25FEF354",
    x"25FE8FD0",
    x"25FE2C73",
    x"25FDC93D",
    x"25FD662E",
    x"25FD0346",
    x"25FCA084",
    x"25FC3DE8",
    x"25FBDB73",
    x"25FB7925",
    x"25FB16FD",
    x"25FAB4FB",
    x"25FA531F",
    x"25F9F16A",
    x"25F98FDA",
    x"25F92E71",
    x"25F8CD2E",
    x"25F86C11",
    x"25F80B1A",
    x"25F7AA48",
    x"25F7499D",
    x"25F6E917",
    x"25F688B7",
    x"25F6287C",
    x"25F5C867",
    x"25F56877",
    x"25F508AD",
    x"25F4A909",
    x"25F44989",
    x"25F3EA2F",
    x"25F38AFA",
    x"25F32BEB",
    x"25F2CD00",
    x"25F26E3A",
    x"25F20F9A",
    x"25F1B11E",
    x"25F152C7",
    x"25F0F495",
    x"25F09688",
    x"25F038A0",
    x"25EFDADC",
    x"25EF7D3D",
    x"25EF1FC2",
    x"25EEC26C",
    x"25EE653A",
    x"25EE082D",
    x"25EDAB44",
    x"25ED4E7F",
    x"25ECF1DE",
    x"25EC9562",
    x"25EC390A",
    x"25EBDCD6",
    x"25EB80C5",
    x"25EB24D9",
    x"25EAC910",
    x"25EA6D6C",
    x"25EA11EB",
    x"25E9B68E",
    x"25E95B54",
    x"25E9003E",
    x"25E8A54C",
    x"25E84A7D",
    x"25E7EFD2",
    x"25E7954A",
    x"25E73AE5",
    x"25E6E0A4",
    x"25E68686",
    x"25E62C8B",
    x"25E5D2B3",
    x"25E578FE",
    x"25E51F6C",
    x"25E4C5FE",
    x"25E46CB2",
    x"25E41389",
    x"25E3BA82",
    x"25E3619F",
    x"25E308DE",
    x"25E2B040",
    x"25E257C4",
    x"25E1FF6B",
    x"25E1A735",
    x"25E14F21",
    x"25E0F72F",
    x"25E09F60",
    x"25E047B2",
    x"25DFF028",
    x"25DF98BF",
    x"25DF4178",
    x"25DEEA54",
    x"25DE9351",
    x"25DE3C71",
    x"25DDE5B2",
    x"25DD8F15",
    x"25DD389A",
    x"25DCE241",
    x"25DC8C09",
    x"25DC35F3",
    x"25DBDFFF",
    x"25DB8A2C",
    x"25DB347B",
    x"25DADEEB",
    x"25DA897D",
    x"25DA3430",
    x"25D9DF04",
    x"25D989FA",
    x"25D93510",
    x"25D8E048",
    x"25D88BA1",
    x"25D8371B",
    x"25D7E2B6",
    x"25D78E72",
    x"25D73A4F",
    x"25D6E64C",
    x"25D6926B",
    x"25D63EAA",
    x"25D5EB0A",
    x"25D5978A",
    x"25D5442B",
    x"25D4F0ED",
    x"25D49DCF",
    x"25D44AD2",
    x"25D3F7F5",
    x"25D3A538",
    x"25D3529C",
    x"25D3001F",
    x"25D2ADC4",
    x"25D25B88",
    x"25D2096C",
    x"25D1B770",
    x"25D16595",
    x"25D113D9",
    x"25D0C23D",
    x"25D070C1",
    x"25D01F65",
    x"25CFCE29",
    x"25CF7D0C",
    x"25CF2C0F",
    x"25CEDB32",
    x"25CE8A74",
    x"25CE39D5",
    x"25CDE956",
    x"25CD98F7",
    x"25CD48B7",
    x"25CCF896",
    x"25CCA895",
    x"25CC58B3",
    x"25CC08EF",
    x"25CBB94C",
    x"25CB69C7",
    x"25CB1A61",
    x"25CACB1A",
    x"25CA7BF2",
    x"25CA2CE9",
    x"25C9DDFF",
    x"25C98F34",
    x"25C94087",
    x"25C8F1F9",
    x"25C8A38A",
    x"25C8553A",
    x"25C80708",
    x"25C7B8F4",
    x"25C76AFF",
    x"25C71D28",
    x"25C6CF70",
    x"25C681D6",
    x"25C6345B",
    x"25C5E6FD",
    x"25C599BE",
    x"25C54C9D",
    x"25C4FF9A",
    x"25C4B2B6",
    x"25C465EF",
    x"25C41946",
    x"25C3CCBB",
    x"25C3804E",
    x"25C333FF",
    x"25C2E7CD",
    x"25C29BBA",
    x"25C24FC4",
    x"25C203EB",
    x"25C1B831",
    x"25C16C93",
    x"25C12114",
    x"25C0D5B2",
    x"25C08A6D",
    x"25C03F45",
    x"25BFF43B",
    x"25BFA94F",
    x"25BF5E7F",
    x"25BF13CD",
    x"25BEC938",
    x"25BE7EC0",
    x"25BE3465",
    x"25BDEA27",
    x"25BDA006",
    x"25BD5602",
    x"25BD0C1A",
    x"25BCC250",
    x"25BC78A3",
    x"25BC2F12",
    x"25BBE59E",
    x"25BB9C46",
    x"25BB530C",
    x"25BB09EE",
    x"25BAC0EC",
    x"25BA7807",
    x"25BA2F3E",
    x"25B9E692",
    x"25B99E02",
    x"25B9558E",
    x"25B90D37",
    x"25B8C4FC",
    x"25B87CDD",
    x"25B834DA",
    x"25B7ECF4",
    x"25B7A529",
    x"25B75D7B",
    x"25B715E8",
    x"25B6CE72",
    x"25B68717",
    x"25B63FD8",
    x"25B5F8B5",
    x"25B5B1AE",
    x"25B56AC2",
    x"25B523F2",
    x"25B4DD3E",
    x"25B496A6",
    x"25B45028",
    x"25B409C7",
    x"25B3C381",
    x"25B37D56",
    x"25B33747",
    x"25B2F153",
    x"25B2AB7A",
    x"25B265BD",
    x"25B2201B",
    x"25B1DA94",
    x"25B19528",
    x"25B14FD7",
    x"25B10AA2",
    x"25B0C587",
    x"25B08087",
    x"25B03BA3",
    x"25AFF6D9",
    x"25AFB22A",
    x"25AF6D96",
    x"25AF291C",
    x"25AEE4BD",
    x"25AEA079",
    x"25AE5C50",
    x"25AE1841",
    x"25ADD44D",
    x"25AD9073",
    x"25AD4CB4",
    x"25AD090F",
    x"25ACC585",
    x"25AC8215",
    x"25AC3EBF",
    x"25ABFB84",
    x"25ABB863",
    x"25AB755C",
    x"25AB326F",
    x"25AAEF9D",
    x"25AAACE4",
    x"25AA6A46",
    x"25AA27C1",
    x"25A9E556",
    x"25A9A306",
    x"25A960CF",
    x"25A91EB2",
    x"25A8DCAF",
    x"25A89AC6",
    x"25A858F6",
    x"25A81740",
    x"25A7D5A4",
    x"25A79421",
    x"25A752B8",
    x"25A71169",
    x"25A6D033",
    x"25A68F16",
    x"25A64E13",
    x"25A60D29",
    x"25A5CC59",
    x"25A58BA1",
    x"25A54B03",
    x"25A50A7F",
    x"25A4CA13",
    x"25A489C1",
    x"25A44988",
    x"25A40967",
    x"25A3C960",
    x"25A38972",
    x"25A3499D",
    x"25A309E1",
    x"25A2CA3D",
    x"25A28AB3",
    x"25A24B41",
    x"25A20BE8",
    x"25A1CCA7",
    x"25A18D80",
    x"25A14E71",
    x"25A10F7B",
    x"25A0D09D",
    x"25A091D8",
    x"25A0532B",
    x"25A01497",
    x"259FD61B",
    x"259F97B7",
    x"259F596C",
    x"259F1B39",
    x"259EDD1F",
    x"259E9F1D",
    x"259E6133",
    x"259E2361",
    x"259DE5A7",
    x"259DA805",
    x"259D6A7C",
    x"259D2D0A",
    x"259CEFB0",
    x"259CB26F",
    x"259C7545",
    x"259C3833",
    x"259BFB39",
    x"259BBE57",
    x"259B818C",
    x"259B44DA",
    x"259B083F",
    x"259ACBBB",
    x"259A8F4F",
    x"259A52FB",
    x"259A16BF",
    x"2599DA99",
    x"25999E8C",
    x"25996296",
    x"259926B7",
    x"2598EAEF",
    x"2598AF3F",
    x"259873A6",
    x"25983825",
    x"2597FCBB",
    x"2597C167",
    x"2597862B",
    x"25974B07",
    x"25970FF9",
    x"2596D502",
    x"25969A22",
    x"25965F5A",
    x"259624A8",
    x"2595EA0D",
    x"2595AF89",
    x"2595751C",
    x"25953AC5",
    x"25950086",
    x"2594C65D",
    x"25948C4B",
    x"2594524F",
    x"2594186B",
    x"2593DE9C",
    x"2593A4E5",
    x"25936B44",
    x"259331B9",
    x"2592F845",
    x"2592BEE7",
    x"259285A0",
    x"25924C6F",
    x"25921354",
    x"2591DA4F",
    x"2591A161",
    x"25916889",
    x"25912FC8",
    x"2590F71C",
    x"2590BE86",
    x"25908607",
    x"25904D9E",
    x"2590154A",
    x"258FDD0D",
    x"258FA4E6",
    x"258F6CD4",
    x"258F34D9",
    x"258EFCF3",
    x"258EC523",
    x"258E8D69",
    x"258E55C5",
    x"258E1E36",
    x"258DE6BD",
    x"258DAF5A",
    x"258D780C",
    x"258D40D4",
    x"258D09B1",
    x"258CD2A4",
    x"258C9BAD",
    x"258C64CB",
    x"258C2DFE",
    x"258BF747",
    x"258BC0A5",
    x"258B8A18",
    x"258B53A1",
    x"258B1D3F",
    x"258AE6F2",
    x"258AB0BA",
    x"258A7A98",
    x"258A448B",
    x"258A0E92",
    x"2589D8AF",
    x"2589A2E1",
    x"25896D28",
    x"25893784",
    x"258901F5",
    x"2588CC7A",
    x"25889715",
    x"258861C4",
    x"25882C88",
    x"2587F761",
    x"2587C24F",
    x"25878D52",
    x"25875869",
    x"25872395",
    x"2586EED5",
    x"2586BA2A",
    x"25868594",
    x"25865112",
    x"25861CA4",
    x"2585E84B",
    x"2585B407",
    x"25857FD7",
    x"25854BBB",
    x"258517B3",
    x"2584E3C0",
    x"2584AFE1",
    x"25847C17",
    x"25844860",
    x"258414BE",
    x"2583E130",
    x"2583ADB6",
    x"25837A51",
    x"258346FF",
    x"258313C1",
    x"2582E097",
    x"2582AD82",
    x"25827A80",
    x"25824792",
    x"258214B8",
    x"2581E1F2",
    x"2581AF3F",
    x"25817CA1",
    x"25814A16",
    x"2581179F",
    x"2580E53B",
    x"2580B2EC",
    x"258080B0",
    x"25804E87",
    x"25801C72",
    x"257FD4E2",
    x"257F7106",
    x"257F0D52",
    x"257EA9C4",
    x"257E465D",
    x"257DE31D",
    x"257D8004",
    x"257D1D11",
    x"257CBA45",
    x"257C579F",
    x"257BF520",
    x"257B92C8",
    x"257B3096",
    x"257ACE8A",
    x"257A6CA4",
    x"257A0AE5",
    x"2579A94C",
    x"257947D9",
    x"2578E68C",
    x"25788565",
    x"25782463",
    x"2577C388",
    x"257762D3",
    x"25770243",
    x"2576A1D9",
    x"25764194",
    x"2575E176",
    x"2575817C",
    x"257521A8",
    x"2574C1FA",
    x"25746271",
    x"2574030D",
    x"2573A3CE",
    x"257344B5",
    x"2572E5C1",
    x"257286F1",
    x"25722847",
    x"2571C9C2",
    x"25716B62",
    x"25710D26",
    x"2570AF0F",
    x"2570511D",
    x"256FF350",
    x"256F95A7",
    x"256F3823",
    x"256EDAC3",
    x"256E7D88",
    x"256E2071",
    x"256DC37F",
    x"256D66B0",
    x"256D0A06",
    x"256CAD81",
    x"256C511F",
    x"256BF4E1",
    x"256B98C8",
    x"256B3CD2",
    x"256AE100",
    x"256A8552",
    x"256A29C8",
    x"2569CE61",
    x"2569731F",
    x"256917FF",
    x"2568BD04",
    x"2568622C",
    x"25680777",
    x"2567ACE6",
    x"25675278",
    x"2566F82D",
    x"25669E06",
    x"25664402",
    x"2565EA21",
    x"25659063",
    x"256536C8",
    x"2564DD50",
    x"256483FB",
    x"25642AC9",
    x"2563D1BA",
    x"256378CD",
    x"25632003",
    x"2562C75C",
    x"25626ED8",
    x"25621676",
    x"2561BE36",
    x"25616619",
    x"25610E1E",
    x"2560B646",
    x"25605E90",
    x"256006FC",
    x"255FAF8A",
    x"255F583B",
    x"255F010D",
    x"255EAA02",
    x"255E5319",
    x"255DFC51",
    x"255DA5AB",
    x"255D4F28",
    x"255CF8C6",
    x"255CA285",
    x"255C4C67",
    x"255BF66A",
    x"255BA08E",
    x"255B4AD4",
    x"255AF53C",
    x"255A9FC5",
    x"255A4A6F",
    x"2559F53A",
    x"2559A027",
    x"25594B35",
    x"2558F664",
    x"2558A1B5",
    x"25584D26",
    x"2557F8B8",
    x"2557A46C",
    x"25575040",
    x"2556FC35",
    x"2556A84B",
    x"25565482",
    x"255600D9",
    x"2555AD51",
    x"255559E9",
    x"255506A3",
    x"2554B37C",
    x"25546076",
    x"25540D91",
    x"2553BACC",
    x"25536827",
    x"255315A2",
    x"2552C33E",
    x"255270FA",
    x"25521ED6",
    x"2551CCD2",
    x"25517AEE",
    x"2551292A",
    x"2550D786",
    x"25508601",
    x"2550349D",
    x"254FE358",
    x"254F9233",
    x"254F412E",
    x"254EF048",
    x"254E9F82",
    x"254E4EDC",
    x"254DFE55",
    x"254DADED",
    x"254D5DA5",
    x"254D0D7C",
    x"254CBD72",
    x"254C6D88",
    x"254C1DBD",
    x"254BCE10",
    x"254B7E84",
    x"254B2F16",
    x"254ADFC7",
    x"254A9097",
    x"254A4186",
    x"2549F294",
    x"2549A3C0",
    x"2549550C",
    x"25490676",
    x"2548B7FF",
    x"254869A6",
    x"25481B6C",
    x"2547CD51",
    x"25477F54",
    x"25473175",
    x"2546E3B5",
    x"25469613",
    x"25464890",
    x"2545FB2A",
    x"2545ADE3",
    x"254560BB",
    x"254513B0",
    x"2544C6C3",
    x"254479F5",
    x"25442D44",
    x"2543E0B1",
    x"2543943C",
    x"254347E5",
    x"2542FBAC",
    x"2542AF91",
    x"25426393",
    x"254217B3",
    x"2541CBF0",
    x"2541804C",
    x"254134C4",
    x"2540E95A",
    x"25409E0E",
    x"254052DF",
    x"254007CD",
    x"253FBCD9",
    x"253F7202",
    x"253F2748",
    x"253EDCAB",
    x"253E922B",
    x"253E47C9",
    x"253DFD83",
    x"253DB35B",
    x"253D694F",
    x"253D1F60",
    x"253CD58E",
    x"253C8BD9",
    x"253C4241",
    x"253BF8C6",
    x"253BAF67",
    x"253B6625",
    x"253B1CFF",
    x"253AD3F6",
    x"253A8B09",
    x"253A4239",
    x"2539F986",
    x"2539B0EE",
    x"25396873",
    x"25392015",
    x"2538D7D2",
    x"25388FAC",
    x"253847A2",
    x"2537FFB4",
    x"2537B7E2",
    x"2537702C",
    x"25372893",
    x"2536E115",
    x"253699B3",
    x"2536526D",
    x"25360B42",
    x"2535C434",
    x"25357D41",
    x"2535366A",
    x"2534EFAF",
    x"2534A90F",
    x"2534628A",
    x"25341C22",
    x"2533D5D4",
    x"25338FA3",
    x"2533498C",
    x"25330391",
    x"2532BDB1",
    x"253277ED",
    x"25323244",
    x"2531ECB6",
    x"2531A743",
    x"253161EB",
    x"25311CAE",
    x"2530D78D",
    x"25309286",
    x"25304D9A",
    x"253008C9",
    x"252FC413",
    x"252F7F78",
    x"252F3AF8",
    x"252EF692",
    x"252EB247",
    x"252E6E17",
    x"252E2A01",
    x"252DE606",
    x"252DA225",
    x"252D5E5F",
    x"252D1AB3",
    x"252CD722",
    x"252C93AB",
    x"252C504F",
    x"252C0D0D",
    x"252BC9E5",
    x"252B86D7",
    x"252B43E3",
    x"252B010A",
    x"252ABE4A",
    x"252A7BA5",
    x"252A391A",
    x"2529F6A9",
    x"2529B451",
    x"25297214",
    x"25292FF0",
    x"2528EDE6",
    x"2528ABF6",
    x"25286A20",
    x"25282863",
    x"2527E6C0",
    x"2527A537",
    x"252763C7",
    x"25272271",
    x"2526E134",
    x"2526A011",
    x"25265F07",
    x"25261E17",
    x"2525DD40",
    x"25259C82",
    x"25255BDD",
    x"25251B52",
    x"2524DAE0",
    x"25249A87",
    x"25245A47",
    x"25241A21",
    x"2523DA13",
    x"25239A1E",
    x"25235A42",
    x"25231A80",
    x"2522DAD6",
    x"25229B45",
    x"25225BCC",
    x"25221C6D",
    x"2521DD26",
    x"25219DF8",
    x"25215EE3",
    x"25211FE6",
    x"2520E102",
    x"2520A236",
    x"25206383",
    x"252024E8",
    x"251FE666",
    x"251FA7FC",
    x"251F69AB",
    x"251F2B72",
    x"251EED51",
    x"251EAF48",
    x"251E7158",
    x"251E3380",
    x"251DF5C0",
    x"251DB818",
    x"251D7A88",
    x"251D3D10",
    x"251CFFB0",
    x"251CC268",
    x"251C8538",
    x"251C4820",
    x"251C0B20",
    x"251BCE38",
    x"251B9167",
    x"251B54AE",
    x"251B180D",
    x"251ADB83",
    x"251A9F11",
    x"251A62B7",
    x"251A2674",
    x"2519EA49",
    x"2519AE35",
    x"25197239",
    x"25193654",
    x"2518FA86",
    x"2518BED0",
    x"25188331",
    x"251847AA",
    x"25180C39",
    x"2517D0E0",
    x"2517959E",
    x"25175A73",
    x"25171F5F",
    x"2516E463",
    x"2516A97D",
    x"25166EAE",
    x"251633F6",
    x"2515F956",
    x"2515BECC",
    x"25158459",
    x"251549FC",
    x"25150FB7",
    x"2514D588",
    x"25149B70",
    x"2514616E",
    x"25142784",
    x"2513EDB0",
    x"2513B3F2",
    x"25137A4B",
    x"251340BA",
    x"25130740",
    x"2512CDDD",
    x"25129490",
    x"25125B59",
    x"25122238",
    x"2511E92E",
    x"2511B03A",
    x"2511775C",
    x"25113E95",
    x"251105E3",
    x"2510CD48",
    x"251094C3",
    x"25105C54",
    x"251023FB",
    x"250FEBB8",
    x"250FB38B",
    x"250F7B74",
    x"250F4372",
    x"250F0B87",
    x"250ED3B1",
    x"250E9BF1",
    x"250E6447",
    x"250E2CB3",
    x"250DF534",
    x"250DBDCB",
    x"250D8678",
    x"250D4F3A",
    x"250D1812",
    x"250CE100",
    x"250CAA02",
    x"250C731B",
    x"250C3C49",
    x"250C058C",
    x"250BCEE4",
    x"250B9852",
    x"250B61D5",
    x"250B2B6E",
    x"250AF51B",
    x"250ABEDE",
    x"250A88B6",
    x"250A52A3",
    x"250A1CA6",
    x"2509E6BD",
    x"2509B0E9",
    x"25097B2B",
    x"25094581",
    x"25090FEC",
    x"2508DA6D",
    x"2508A502",
    x"25086FAC",
    x"25083A6A",
    x"2508053E",
    x"2507D026",
    x"25079B23",
    x"25076635",
    x"2507315C",
    x"2506FC97",
    x"2506C7E6",
    x"2506934A",
    x"25065EC3",
    x"25062A50",
    x"2505F5F2",
    x"2505C1A8",
    x"25058D73",
    x"25055952",
    x"25052545",
    x"2504F14D",
    x"2504BD68",
    x"25048999",
    x"250455DD",
    x"25042235",
    x"2503EEA2",
    x"2503BB23",
    x"250387B8",
    x"25035461",
    x"2503211E",
    x"2502EDEF",
    x"2502BAD4",
    x"250287CD",
    x"250254DA",
    x"250221FB",
    x"2501EF2F",
    x"2501BC78",
    x"250189D4",
    x"25015744",
    x"250124C8",
    x"2500F25F",
    x"2500C00B",
    x"25008DC9",
    x"25005B9C",
    x"25002982",
    x"24FFEEF7",
    x"24FF8B11",
    x"24FF2752",
    x"24FEC3BA",
    x"24FE6049",
    x"24FDFCFF",
    x"24FD99DC",
    x"24FD36DF",
    x"24FCD409",
    x"24FC7159",
    x"24FC0ED0",
    x"24FBAC6E",
    x"24FB4A31",
    x"24FAE81C",
    x"24FA862C",
    x"24FA2463",
    x"24F9C2C0",
    x"24F96143",
    x"24F8FFEC",
    x"24F89EBB",
    x"24F83DB0",
    x"24F7DCCA",
    x"24F77C0B",
    x"24F71B71",
    x"24F6BAFE",
    x"24F65AAF",
    x"24F5FA87",
    x"24F59A84",
    x"24F53AA6",
    x"24F4DAEE",
    x"24F47B5B",
    x"24F41BED",
    x"24F3BCA5",
    x"24F35D82",
    x"24F2FE84",
    x"24F29FAB",
    x"24F240F7",
    x"24F1E268",
    x"24F183FE",
    x"24F125B9",
    x"24F0C799",
    x"24F0699D",
    x"24F00BC6",
    x"24EFAE14",
    x"24EF5086",
    x"24EEF31D",
    x"24EE95D8",
    x"24EE38B8",
    x"24EDDBBC",
    x"24ED7EE4",
    x"24ED2231",
    x"24ECC5A2",
    x"24EC6936",
    x"24EC0CEF",
    x"24EBB0CC",
    x"24EB54CD",
    x"24EAF8F2",
    x"24EA9D3B",
    x"24EA41A7",
    x"24E9E637",
    x"24E98AEB",
    x"24E92FC3",
    x"24E8D4BE",
    x"24E879DD",
    x"24E81F1F",
    x"24E7C484",
    x"24E76A0D",
    x"24E70FB9",
    x"24E6B589",
    x"24E65B7C",
    x"24E60191",
    x"24E5A7CA",
    x"24E54E26",
    x"24E4F4A5",
    x"24E49B47",
    x"24E4420C",
    x"24E3E8F4",
    x"24E38FFE",
    x"24E3372B",
    x"24E2DE7B",
    x"24E285ED",
    x"24E22D82",
    x"24E1D53A",
    x"24E17D14",
    x"24E12510",
    x"24E0CD2F",
    x"24E07570",
    x"24E01DD3",
    x"24DFC658",
    x"24DF6F00",
    x"24DF17CA",
    x"24DEC0B5",
    x"24DE69C3",
    x"24DE12F3",
    x"24DDBC44",
    x"24DD65B8",
    x"24DD0F4D",
    x"24DCB904",
    x"24DC62DC",
    x"24DC0CD6",
    x"24DBB6F2",
    x"24DB612F",
    x"24DB0B8E",
    x"24DAB60E",
    x"24DA60B0",
    x"24DA0B73",
    x"24D9B657",
    x"24D9615C",
    x"24D90C83",
    x"24D8B7CB",
    x"24D86333",
    x"24D80EBD",
    x"24D7BA68",
    x"24D76633",
    x"24D71220",
    x"24D6BE2D",
    x"24D66A5B",
    x"24D616AA",
    x"24D5C31A",
    x"24D56FAA",
    x"24D51C5A",
    x"24D4C92B",
    x"24D4761D",
    x"24D4232F",
    x"24D3D062",
    x"24D37DB4",
    x"24D32B27",
    x"24D2D8BB",
    x"24D2866E",
    x"24D23442",
    x"24D1E235",
    x"24D19049",
    x"24D13E7C",
    x"24D0ECD0",
    x"24D09B43",
    x"24D049D7",
    x"24CFF88A",
    x"24CFA75D",
    x"24CF564F",
    x"24CF0561",
    x"24CEB493",
    x"24CE63E4",
    x"24CE1355",
    x"24CDC2E5",
    x"24CD7294",
    x"24CD2263",
    x"24CCD252",
    x"24CC825F",
    x"24CC328C",
    x"24CBE2D8",
    x"24CB9342",
    x"24CB43CC",
    x"24CAF475",
    x"24CAA53D",
    x"24CA5624",
    x"24CA072A",
    x"24C9B84F",
    x"24C96992",
    x"24C91AF4",
    x"24C8CC75",
    x"24C87E15",
    x"24C82FD3",
    x"24C7E1AF",
    x"24C793AA",
    x"24C745C4",
    x"24C6F7FC",
    x"24C6AA52",
    x"24C65CC7",
    x"24C60F5A",
    x"24C5C20B",
    x"24C574DA",
    x"24C527C7",
    x"24C4DAD3",
    x"24C48DFC",
    x"24C44144",
    x"24C3F4A9",
    x"24C3A82D",
    x"24C35BCE",
    x"24C30F8D",
    x"24C2C36A",
    x"24C27764",
    x"24C22B7C",
    x"24C1DFB2",
    x"24C19406",
    x"24C14877",
    x"24C0FD05",
    x"24C0B1B1",
    x"24C0667A",
    x"24C01B61",
    x"24BFD065",
    x"24BF8586",
    x"24BF3AC5",
    x"24BEF020",
    x"24BEA599",
    x"24BE5B2F",
    x"24BE10E2",
    x"24BDC6B2",
    x"24BD7C9E",
    x"24BD32A8",
    x"24BCE8CF",
    x"24BC9F12",
    x"24BC5573",
    x"24BC0BF0",
    x"24BBC289",
    x"24BB7940",
    x"24BB3012",
    x"24BAE702",
    x"24BA9E0E",
    x"24BA5536",
    x"24BA0C7B",
    x"24B9C3DD",
    x"24B97B5A",
    x"24B932F4",
    x"24B8EAAB",
    x"24B8A27D",
    x"24B85A6C",
    x"24B81276",
    x"24B7CA9D",
    x"24B782E0",
    x"24B73B3F",
    x"24B6F3BA",
    x"24B6AC50",
    x"24B66503",
    x"24B61DD1",
    x"24B5D6BC",
    x"24B58FC2",
    x"24B548E3",
    x"24B50221",
    x"24B4BB7A",
    x"24B474EE",
    x"24B42E7E",
    x"24B3E82A",
    x"24B3A1F1",
    x"24B35BD3",
    x"24B315D1",
    x"24B2CFEA",
    x"24B28A1F",
    x"24B2446E",
    x"24B1FED9",
    x"24B1B95F",
    x"24B17400",
    x"24B12EBD",
    x"24B0E994",
    x"24B0A486",
    x"24B05F93",
    x"24B01ABC",
    x"24AFD5FE",
    x"24AF915C",
    x"24AF4CD5",
    x"24AF0868",
    x"24AEC416",
    x"24AE7FDF",
    x"24AE3BC2",
    x"24ADF7C0",
    x"24ADB3D9",
    x"24AD700C",
    x"24AD2C59",
    x"24ACE8C1",
    x"24ACA543",
    x"24AC61E0",
    x"24AC1E97",
    x"24ABDB68",
    x"24AB9854",
    x"24AB5559",
    x"24AB1279",
    x"24AACFB3",
    x"24AA8D07",
    x"24AA4A74",
    x"24AA07FC",
    x"24A9C59E",
    x"24A9835A",
    x"24A94130",
    x"24A8FF1F",
    x"24A8BD28",
    x"24A87B4B",
    x"24A83988",
    x"24A7F7DE",
    x"24A7B64E",
    x"24A774D8",
    x"24A7337B",
    x"24A6F238",
    x"24A6B10E",
    x"24A66FFD",
    x"24A62F06",
    x"24A5EE29",
    x"24A5AD64",
    x"24A56CB9",
    x"24A52C27",
    x"24A4EBAF",
    x"24A4AB4F",
    x"24A46B09",
    x"24A42ADB",
    x"24A3EAC7",
    x"24A3AACC",
    x"24A36AEA",
    x"24A32B20",
    x"24A2EB70",
    x"24A2ABD9",
    x"24A26C5A",
    x"24A22CF4",
    x"24A1EDA7",
    x"24A1AE72",
    x"24A16F56",
    x"24A13053",
    x"24A0F169",
    x"24A0B297",
    x"24A073DD",
    x"24A0353C",
    x"249FF6B3",
    x"249FB843",
    x"249F79EB",
    x"249F3BAC",
    x"249EFD85",
    x"249EBF76",
    x"249E817F",
    x"249E43A1",
    x"249E05DA",
    x"249DC82C",
    x"249D8A96",
    x"249D4D18",
    x"249D0FB2",
    x"249CD264",
    x"249C952D",
    x"249C580F",
    x"249C1B09",
    x"249BDE1A",
    x"249BA143",
    x"249B6484",
    x"249B27DD",
    x"249AEB4D",
    x"249AAED5",
    x"249A7274",
    x"249A362B",
    x"2499F9FA",
    x"2499BDE0",
    x"249981DE",
    x"249945F2",
    x"24990A1F",
    x"2498CE63",
    x"249892BE",
    x"24985730",
    x"24981BB9",
    x"2497E05A",
    x"2497A512",
    x"249769E1",
    x"24972EC7",
    x"2496F3C5",
    x"2496B8D9",
    x"24967E04",
    x"24964347",
    x"249608A0",
    x"2495CE10",
    x"24959397",
    x"24955934",
    x"24951EE9",
    x"2494E4B4",
    x"2494AA96",
    x"2494708F",
    x"2494369E",
    x"2493FCC4",
    x"2493C301",
    x"24938954",
    x"24934FBE",
    x"2493163E",
    x"2492DCD4",
    x"2492A381",
    x"24926A44",
    x"2492311E",
    x"2491F80E",
    x"2491BF14",
    x"24918631",
    x"24914D63",
    x"249114AC",
    x"2490DC0B",
    x"2490A380",
    x"24906B0C",
    x"249032AD",
    x"248FFA64",
    x"248FC231",
    x"248F8A14",
    x"248F520D",
    x"248F1A1C",
    x"248EE241",
    x"248EAA7B",
    x"248E72CC",
    x"248E3B32",
    x"248E03AD",
    x"248DCC3F",
    x"248D94E6",
    x"248D5DA2",
    x"248D2675",
    x"248CEF5C",
    x"248CB85A",
    x"248C816C",
    x"248C4A95",
    x"248C13D2",
    x"248BDD25",
    x"248BA68D",
    x"248B700B",
    x"248B399E",
    x"248B0346",
    x"248ACD03",
    x"248A96D6",
    x"248A60BD",
    x"248A2ABA",
    x"2489F4CC",
    x"2489BEF3",
    x"2489892F",
    x"24895380",
    x"24891DE6",
    x"2488E860",
    x"2488B2F0",
    x"24887D94",
    x"2488484E",
    x"2488131C",
    x"2487DDFF",
    x"2487A8F7",
    x"24877403",
    x"24873F24",
    x"24870A5A",
    x"2486D5A4",
    x"2486A103",
    x"24866C76",
    x"248637FE",
    x"2486039A",
    x"2485CF4B",
    x"24859B10",
    x"248566EA",
    x"248532D8",
    x"2484FEDA",
    x"2484CAF1",
    x"2484971C",
    x"2484635B",
    x"24842FAE",
    x"2483FC15",
    x"2483C891",
    x"24839521",
    x"248361C5",
    x"24832E7C",
    x"2482FB48",
    x"2482C828",
    x"2482951C",
    x"24826224",
    x"24822F3F",
    x"2481FC6F",
    x"2481C9B2",
    x"24819709",
    x"24816474",
    x"248131F3",
    x"2480FF85",
    x"2480CD2B",
    x"24809AE5",
    x"248068B2",
    x"24803693",
    x"24800487",
    x"247FA51E",
    x"247F4155",
    x"247EDDB3",
    x"247E7A38",
    x"247E16E4",
    x"247DB3B6",
    x"247D50AF",
    x"247CEDCF",
    x"247C8B16",
    x"247C2883",
    x"247BC616",
    x"247B63D0",
    x"247B01B0",
    x"247A9FB6",
    x"247A3DE3",
    x"2479DC36",
    x"24797AAF",
    x"2479194E",
    x"2478B813",
    x"247856FE",
    x"2477F60F",
    x"24779546",
    x"247734A3",
    x"2476D425",
    x"247673CD",
    x"2476139A",
    x"2475B38E",
    x"247553A6",
    x"2474F3E4",
    x"24749448",
    x"247434D0",
    x"2473D57E",
    x"24737652",
    x"2473174A",
    x"2472B867",
    x"247259AA",
    x"2471FB11",
    x"24719C9E",
    x"24713E4F",
    x"2470E025",
    x"24708220",
    x"2470243F",
    x"246FC683",
    x"246F68EC",
    x"246F0B79",
    x"246EAE2B",
    x"246E5101",
    x"246DF3FC",
    x"246D971B",
    x"246D3A5E",
    x"246CDDC5",
    x"246C8151",
    x"246C2500",
    x"246BC8D4",
    x"246B6CCB",
    x"246B10E7",
    x"246AB526",
    x"246A5989",
    x"2469FE10",
    x"2469A2BB",
    x"24694789",
    x"2468EC7B",
    x"24689190",
    x"246836C9",
    x"2467DC25",
    x"246781A5",
    x"24672748",
    x"2466CD0E",
    x"246672F8",
    x"24661904",
    x"2465BF34",
    x"24656587",
    x"24650BFD",
    x"2464B296",
    x"24645951",
    x"24640030",
    x"2463A731",
    x"24634E55",
    x"2462F59C",
    x"24629D05",
    x"24624491",
    x"2461EC40",
    x"24619411",
    x"24613C04",
    x"2460E41A",
    x"24608C52",
    x"246034AC",
    x"245FDD29",
    x"245F85C7",
    x"245F2E88",
    x"245ED76B",
    x"245E8070",
    x"245E2997",
    x"245DD2DF",
    x"245D7C4A",
    x"245D25D6",
    x"245CCF84",
    x"245C7954",
    x"245C2345",
    x"245BCD58",
    x"245B778D",
    x"245B21E3",
    x"245ACC5A",
    x"245A76F3",
    x"245A21AE",
    x"2459CC89",
    x"24597786",
    x"245922A4",
    x"2458CDE3",
    x"24587943",
    x"245824C4",
    x"2457D066",
    x"24577C29",
    x"2457280D",
    x"2456D412",
    x"24568037",
    x"24562C7E",
    x"2455D8E5",
    x"2455856C",
    x"24553214",
    x"2454DEDD",
    x"24548BC6",
    x"245438D0",
    x"2453E5FA",
    x"24539344",
    x"245340AF",
    x"2452EE3A",
    x"24529BE5",
    x"245249B0",
    x"2451F79B",
    x"2451A5A6",
    x"245153D2",
    x"2451021D",
    x"2450B088",
    x"24505F13",
    x"24500DBE",
    x"244FBC88",
    x"244F6B72",
    x"244F1A7C",
    x"244EC9A6",
    x"244E78EF",
    x"244E2857",
    x"244DD7DF",
    x"244D8786",
    x"244D374D",
    x"244CE733",
    x"244C9738",
    x"244C475D",
    x"244BF7A1",
    x"244BA804",
    x"244B5885",
    x"244B0926",
    x"244AB9E6",
    x"244A6AC5",
    x"244A1BC3",
    x"2449CCDF",
    x"24497E1B",
    x"24492F75",
    x"2448E0EE",
    x"24489285",
    x"2448443B",
    x"2447F610",
    x"2447A803",
    x"24475A15",
    x"24470C45",
    x"2446BE93",
    x"24467100",
    x"2446238B",
    x"2445D634",
    x"244588FB",
    x"24453BE1",
    x"2444EEE4",
    x"2444A206",
    x"24445546",
    x"244408A4",
    x"2443BC1F",
    x"24436FB9",
    x"24432370",
    x"2442D745",
    x"24428B38",
    x"24423F48",
    x"2441F376",
    x"2441A7C2",
    x"24415C2B",
    x"244110B2",
    x"2440C556",
    x"24407A18",
    x"24402EF7",
    x"243FE3F3",
    x"243F990D",
    x"243F4E43",
    x"243F0397",
    x"243EB909",
    x"243E6E97",
    x"243E2442",
    x"243DDA0A",
    x"243D8FF0",
    x"243D45F2",
    x"243CFC11",
    x"243CB24D",
    x"243C68A6",
    x"243C1F1B",
    x"243BD5AD",
    x"243B8C5C",
    x"243B4328",
    x"243AFA10",
    x"243AB114",
    x"243A6836",
    x"243A1F73",
    x"2439D6CD",
    x"24398E43",
    x"243945D6",
    x"2438FD85",
    x"2438B550",
    x"24386D37",
    x"2438253A",
    x"2437DD5A",
    x"24379595",
    x"24374DED",
    x"24370661",
    x"2436BEF0",
    x"2436779B",
    x"24363063",
    x"2435E946",
    x"2435A244",
    x"24355B5F",
    x"24351495",
    x"2434CDE7",
    x"24348754",
    x"243440DD",
    x"2433FA81",
    x"2433B441",
    x"24336E1C",
    x"24332813",
    x"2432E225",
    x"24329C52",
    x"2432569B",
    x"243210FF",
    x"2431CB7E",
    x"24318618",
    x"243140CD",
    x"2430FB9D",
    x"2430B688",
    x"2430718F",
    x"24302CB0",
    x"242FE7EC",
    x"242FA342",
    x"242F5EB4",
    x"242F1A40",
    x"242ED5E8",
    x"242E91A9",
    x"242E4D86",
    x"242E097D",
    x"242DC58E",
    x"242D81BA",
    x"242D3E01",
    x"242CFA62",
    x"242CB6DD",
    x"242C7373",
    x"242C3023",
    x"242BECED",
    x"242BA9D2",
    x"242B66D1",
    x"242B23EA",
    x"242AE11D",
    x"242A9E6A",
    x"242A5BD1",
    x"242A1952",
    x"2429D6ED",
    x"242994A2",
    x"24295271",
    x"2429105A",
    x"2428CE5C",
    x"24288C78",
    x"24284AAE",
    x"242808FE",
    x"2427C767",
    x"242785EA",
    x"24274487",
    x"2427033D",
    x"2426C20C",
    x"242680F5",
    x"24263FF7",
    x"2425FF13",
    x"2425BE48",
    x"24257D96",
    x"24253CFE",
    x"2424FC7F",
    x"2424BC19",
    x"24247BCC",
    x"24243B98",
    x"2423FB7D",
    x"2423BB7C",
    x"24237B93",
    x"24233BC3",
    x"2422FC0C",
    x"2422BC6E",
    x"24227CE9",
    x"24223D7C",
    x"2421FE29",
    x"2421BEEE",
    x"24217FCC",
    x"242140C2",
    x"242101D1",
    x"2420C2F9",
    x"24208439",
    x"24204591",
    x"24200702",
    x"241FC88C",
    x"241F8A2E",
    x"241F4BE8",
    x"241F0DBA",
    x"241ECFA5",
    x"241E91A8",
    x"241E53C3",
    x"241E15F7",
    x"241DD842",
    x"241D9AA6",
    x"241D5D21",
    x"241D1FB5",
    x"241CE261",
    x"241CA524",
    x"241C67FF",
    x"241C2AF3",
    x"241BEDFE",
    x"241BB121",
    x"241B745C",
    x"241B37AE",
    x"241AFB18",
    x"241ABE9A",
    x"241A8233",
    x"241A45E4",
    x"241A09AC",
    x"2419CD8C",
    x"24199184",
    x"24195593",
    x"241919B9",
    x"2418DDF7",
    x"2418A24C",
    x"241866B8",
    x"24182B3B",
    x"2417EFD6",
    x"2417B488",
    x"24177951",
    x"24173E31",
    x"24170328",
    x"2416C837",
    x"24168D5C",
    x"24165298",
    x"241617EB",
    x"2415DD56",
    x"2415A2D6",
    x"2415686E",
    x"24152E1D",
    x"2414F3E2",
    x"2414B9BE",
    x"24147FB1",
    x"241445BB",
    x"24140BDB",
    x"2413D211",
    x"2413985F",
    x"24135EC2",
    x"2413253C",
    x"2412EBCD",
    x"2412B274",
    x"24127932",
    x"24124006",
    x"241206F0",
    x"2411CDF0",
    x"24119507",
    x"24115C34",
    x"24112377",
    x"2410EAD0",
    x"2410B23F",
    x"241079C5",
    x"24104160",
    x"24100912",
    x"240FD0D9",
    x"240F98B6",
    x"240F60AA",
    x"240F28B3",
    x"240EF0D2",
    x"240EB907",
    x"240E8151",
    x"240E49B2",
    x"240E1228",
    x"240DDAB4",
    x"240DA355",
    x"240D6C0C",
    x"240D34D8",
    x"240CFDBB",
    x"240CC6B2",
    x"240C8FBF",
    x"240C58E2",
    x"240C221A",
    x"240BEB67",
    x"240BB4CA",
    x"240B7E42",
    x"240B47CF",
    x"240B1172",
    x"240ADB2A",
    x"240AA4F7",
    x"240A6ED9",
    x"240A38D0",
    x"240A02DC",
    x"2409CCFE",
    x"24099734",
    x"24096180",
    x"24092BE0",
    x"2408F655",
    x"2408C0E0",
    x"24088B7F",
    x"24085633",
    x"240820FB",
    x"2407EBD9",
    x"2407B6CB",
    x"240781D2",
    x"24074CEE",
    x"2407181E",
    x"2406E363",
    x"2406AEBC",
    x"24067A2A",
    x"240645AD",
    x"24061144",
    x"2405DCEF",
    x"2405A8AF",
    x"24057484",
    x"2405406C",
    x"24050C69",
    x"2404D87A",
    x"2404A4A0",
    x"240470DA",
    x"24043D28",
    x"2404098A",
    x"2403D600",
    x"2403A28B",
    x"24036F29",
    x"24033BDC",
    x"240308A3",
    x"2402D57D",
    x"2402A26C",
    x"24026F6E",
    x"24023C85",
    x"240209AF",
    x"2401D6ED",
    x"2401A43F",
    x"240171A5",
    x"24013F1E",
    x"24010CAC",
    x"2400DA4C",
    x"2400A801",
    x"240075C9",
    x"240043A5",
    x"24001194",
    x"23FFBF2E",
    x"23FF5B5B",
    x"23FEF7AF",
    x"23FE942A",
    x"23FE30CB",
    x"23FDCD94",
    x"23FD6A83",
    x"23FD0798",
    x"23FCA4D5",
    x"23FC4238",
    x"23FBDFC1",
    x"23FB7D71",
    x"23FB1B47",
    x"23FAB943",
    x"23FA5766",
    x"23F9F5AF",
    x"23F9941E",
    x"23F932B3",
    x"23F8D16F",
    x"23F87050",
    x"23F80F57",
    x"23F7AE84",
    x"23F74DD6",
    x"23F6ED4F",
    x"23F68CED",
    x"23F62CB1",
    x"23F5CC9A",
    x"23F56CA9",
    x"23F50CDD",
    x"23F4AD37",
    x"23F44DB6",
    x"23F3EE5A",
    x"23F38F24",
    x"23F33012",
    x"23F2D126",
    x"23F2725F",
    x"23F213BD",
    x"23F1B53F",
    x"23F156E7",
    x"23F0F8B4",
    x"23F09AA5",
    x"23F03CBB",
    x"23EFDEF5",
    x"23EF8154",
    x"23EF23D8",
    x"23EEC680",
    x"23EE694D",
    x"23EE0C3E",
    x"23EDAF54",
    x"23ED528D",
    x"23ECF5EB",
    x"23EC996D",
    x"23EC3D13",
    x"23EBE0DD",
    x"23EB84CB",
    x"23EB28DE",
    x"23EACD14",
    x"23EA716D",
    x"23EA15EB",
    x"23E9BA8C",
    x"23E95F51",
    x"23E9043A",
    x"23E8A946",
    x"23E84E75",
    x"23E7F3C8",
    x"23E7993F",
    x"23E73ED9",
    x"23E6E496",
    x"23E68A76",
    x"23E6307A",
    x"23E5D6A0",
    x"23E57CEA",
    x"23E52357",
    x"23E4C9E6",
    x"23E47099",
    x"23E4176E",
    x"23E3BE67",
    x"23E36582",
    x"23E30CBF",
    x"23E2B420",
    x"23E25BA3",
    x"23E20348",
    x"23E1AB10",
    x"23E152FA",
    x"23E0FB07",
    x"23E0A336",
    x"23E04B88",
    x"23DFF3FB",
    x"23DF9C91",
    x"23DF4549",
    x"23DEEE23",
    x"23DE971F",
    x"23DE403D",
    x"23DDE97D",
    x"23DD92DE",
    x"23DD3C62",
    x"23DCE607",
    x"23DC8FCE",
    x"23DC39B7",
    x"23DBE3C1",
    x"23DB8DED",
    x"23DB383A",
    x"23DAE2A9",
    x"23DA8D39",
    x"23DA37EA",
    x"23D9E2BD",
    x"23D98DB1",
    x"23D938C7",
    x"23D8E3FD",
    x"23D88F54",
    x"23D83ACD",
    x"23D7E666",
    x"23D79221",
    x"23D73DFC",
    x"23D6E9F9",
    x"23D69616",
    x"23D64253",
    x"23D5EEB2",
    x"23D59B31",
    x"23D547D0",
    x"23D4F491",
    x"23D4A171",
    x"23D44E72",
    x"23D3FB94",
    x"23D3A8D6",
    x"23D35638",
    x"23D303BB",
    x"23D2B15D",
    x"23D25F20",
    x"23D20D03",
    x"23D1BB06",
    x"23D16929",
    x"23D1176C",
    x"23D0C5CE",
    x"23D07451",
    x"23D022F4",
    x"23CFD1B6",
    x"23CF8098",
    x"23CF2F99",
    x"23CEDEBA",
    x"23CE8DFB",
    x"23CE3D5C",
    x"23CDECDB",
    x"23CD9C7A",
    x"23CD4C39",
    x"23CCFC17",
    x"23CCAC14",
    x"23CC5C30",
    x"23CC0C6C",
    x"23CBBCC7",
    x"23CB6D41",
    x"23CB1DD9",
    x"23CACE91",
    x"23CA7F68",
    x"23CA305E",
    x"23C9E172",
    x"23C992A5",
    x"23C943F8",
    x"23C8F568",
    x"23C8A6F8",
    x"23C858A6",
    x"23C80A73",
    x"23C7BC5E",
    x"23C76E67",
    x"23C7208F",
    x"23C6D2D6",
    x"23C6853B",
    x"23C637BE",
    x"23C5EA5F",
    x"23C59D1F",
    x"23C54FFC",
    x"23C502F8",
    x"23C4B612",
    x"23C4694A",
    x"23C41CA0",
    x"23C3D014",
    x"23C383A5",
    x"23C33755",
    x"23C2EB22",
    x"23C29F0D",
    x"23C25316",
    x"23C2073C",
    x"23C1BB80",
    x"23C16FE2",
    x"23C12461",
    x"23C0D8FD",
    x"23C08DB7",
    x"23C0428E",
    x"23BFF783",
    x"23BFAC95",
    x"23BF61C4",
    x"23BF1711",
    x"23BECC7A",
    x"23BE8201",
    x"23BE37A5",
    x"23BDED65",
    x"23BDA343",
    x"23BD593E",
    x"23BD0F55",
    x"23BCC58A",
    x"23BC7BDB",
    x"23BC3249",
    x"23BBE8D4",
    x"23BB9F7B",
    x"23BB563F",
    x"23BB0D20",
    x"23BAC41D",
    x"23BA7B37",
    x"23BA326D",
    x"23B9E9BF",
    x"23B9A12E",
    x"23B958B9",
    x"23B91061",
    x"23B8C824",
    x"23B88004",
    x"23B83800",
    x"23B7F019",
    x"23B7A84D",
    x"23B7609D",
    x"23B71909",
    x"23B6D191",
    x"23B68A36",
    x"23B642F5",
    x"23B5FBD1",
    x"23B5B4C9",
    x"23B56DDC",
    x"23B5270B",
    x"23B4E055",
    x"23B499BC",
    x"23B4533D",
    x"23B40CDB",
    x"23B3C693",
    x"23B38067",
    x"23B33A57",
    x"23B2F462",
    x"23B2AE88",
    x"23B268C9",
    x"23B22326",
    x"23B1DD9E",
    x"23B19831",
    x"23B152DF",
    x"23B10DA8",
    x"23B0C88C",
    x"23B0838B",
    x"23B03EA6",
    x"23AFF9DB",
    x"23AFB52A",
    x"23AF7095",
    x"23AF2C1A",
    x"23AEE7BB",
    x"23AEA375",
    x"23AE5F4B",
    x"23AE1B3B",
    x"23ADD746",
    x"23AD936B",
    x"23AD4FAA",
    x"23AD0C04",
    x"23ACC879",
    x"23AC8508",
    x"23AC41B1",
    x"23ABFE74",
    x"23ABBB52",
    x"23AB784A",
    x"23AB355C",
    x"23AAF288",
    x"23AAAFCF",
    x"23AA6D2F",
    x"23AA2AA9",
    x"23A9E83E",
    x"23A9A5EC",
    x"23A963B4",
    x"23A92196",
    x"23A8DF92",
    x"23A89DA7",
    x"23A85BD7",
    x"23A81A20",
    x"23A7D882",
    x"23A796FE",
    x"23A75594",
    x"23A71444",
    x"23A6D30C",
    x"23A691EF",
    x"23A650EA",
    x"23A60FFF",
    x"23A5CF2E",
    x"23A58E76",
    x"23A54DD7",
    x"23A50D51",
    x"23A4CCE4",
    x"23A48C91",
    x"23A44C56",
    x"23A40C35",
    x"23A3CC2D",
    x"23A38C3D",
    x"23A34C67",
    x"23A30CAA",
    x"23A2CD05",
    x"23A28D7A",
    x"23A24E07",
    x"23A20EAD",
    x"23A1CF6B",
    x"23A19043",
    x"23A15133",
    x"23A1123B",
    x"23A0D35C",
    x"23A09496",
    x"23A055E8",
    x"23A01753",
    x"239FD8D6",
    x"239F9A71",
    x"239F5C25",
    x"239F1DF1",
    x"239EDFD6",
    x"239EA1D3",
    x"239E63E7",
    x"239E2614",
    x"239DE85A",
    x"239DAAB7",
    x"239D6D2C",
    x"239D2FBA",
    x"239CF25F",
    x"239CB51C",
    x"239C77F1",
    x"239C3ADF",
    x"239BFDE3",
    x"239BC100",
    x"239B8435",
    x"239B4781",
    x"239B0AE5",
    x"239ACE60",
    x"239A91F4",
    x"239A559E",
    x"239A1961",
    x"2399DD3B",
    x"2399A12C",
    x"23996535",
    x"23992955",
    x"2398ED8C",
    x"2398B1DB",
    x"23987641",
    x"23983ABF",
    x"2397FF53",
    x"2397C3FF",
    x"239788C2",
    x"23974D9C",
    x"2397128E",
    x"2396D796",
    x"23969CB5",
    x"239661EB",
    x"23962739",
    x"2395EC9D",
    x"2395B218",
    x"239577AA",
    x"23953D52",
    x"23950312",
    x"2394C8E8",
    x"23948ED5",
    x"239454D8",
    x"23941AF2",
    x"2393E123",
    x"2393A76B",
    x"23936DC8",
    x"2393343D",
    x"2392FAC8",
    x"2392C169",
    x"23928821",
    x"23924EEF",
    x"239215D3",
    x"2391DCCD",
    x"2391A3DE",
    x"23916B05",
    x"23913243",
    x"2390F996",
    x"2390C100",
    x"2390887F",
    x"23905015",
    x"239017C1",
    x"238FDF82",
    x"238FA75A",
    x"238F6F48",
    x"238F374B",
    x"238EFF65",
    x"238EC794",
    x"238E8FD9",
    x"238E5833",
    x"238E20A4",
    x"238DE92A",
    x"238DB1C5",
    x"238D7A77",
    x"238D433E",
    x"238D0C1A",
    x"238CD50C",
    x"238C9E14",
    x"238C6731",
    x"238C3063",
    x"238BF9AB",
    x"238BC308",
    x"238B8C7B",
    x"238B5602",
    x"238B1F9F",
    x"238AE952",
    x"238AB319",
    x"238A7CF6",
    x"238A46E8",
    x"238A10EE",
    x"2389DB0A",
    x"2389A53B",
    x"23896F81",
    x"238939DC",
    x"2389044C",
    x"2388CED1",
    x"2388996A",
    x"23886419",
    x"23882EDC",
    x"2387F9B4",
    x"2387C4A1",
    x"23878FA3",
    x"23875AB9",
    x"238725E4",
    x"2386F123",
    x"2386BC77",
    x"238687E0",
    x"2386535D",
    x"23861EEF",
    x"2385EA95",
    x"2385B650",
    x"2385821F",
    x"23854E02",
    x"238519FA",
    x"2384E606",
    x"2384B226",
    x"23847E5A",
    x"23844AA3",
    x"23841700",
    x"2383E371",
    x"2383AFF6",
    x"23837C90",
    x"2383493D",
    x"238315FE",
    x"2382E2D4",
    x"2382AFBD",
    x"23827CBB",
    x"238249CC",
    x"238216F1",
    x"2381E42A",
    x"2381B177",
    x"23817ED7",
    x"23814C4C",
    x"238119D4",
    x"2380E76F",
    x"2380B51F",
    x"238082E2",
    x"238050B9",
    x"23801EA3",
    x"237FD941",
    x"237F7564",
    x"237F11AD",
    x"237EAE1E",
    x"237E4AB5",
    x"237DE774",
    x"237D8459",
    x"237D2164",
    x"237CBE96",
    x"237C5BEF",
    x"237BF96F",
    x"237B9714",
    x"237B34E1",
    x"237AD2D3",
    x"237A70EC",
    x"237A0F2B",
    x"2379AD90",
    x"23794C1B",
    x"2378EACC",
    x"237889A4",
    x"237828A1",
    x"2377C7C4",
    x"2377670D",
    x"2377067B",
    x"2376A610",
    x"237645CA",
    x"2375E5A9",
    x"237585AE",
    x"237525D9",
    x"2374C629",
    x"2374669E",
    x"23740738",
    x"2373A7F8",
    x"237348DD",
    x"2372E9E7",
    x"23728B16",
    x"23722C6B",
    x"2371CDE4",
    x"23716F82",
    x"23711145",
    x"2370B32C",
    x"23705539",
    x"236FF76A",
    x"236F99BF",
    x"236F3C3A",
    x"236EDED8",
    x"236E819B",
    x"236E2483",
    x"236DC78F",
    x"236D6ABF",
    x"236D0E13",
    x"236CB18C",
    x"236C5529",
    x"236BF8E9",
    x"236B9CCE",
    x"236B40D7",
    x"236AE504",
    x"236A8954",
    x"236A2DC8",
    x"2369D260",
    x"2369771C",
    x"23691BFB",
    x"2368C0FE",
    x"23686624",
    x"23680B6E",
    x"2367B0DB",
    x"2367566C",
    x"2366FC20",
    x"2366A1F7",
    x"236647F1",
    x"2365EE0F",
    x"2365944F",
    x"23653AB3",
    x"2364E139",
    x"236487E3",
    x"23642EAF",
    x"2363D59E",
    x"23637CB0",
    x"236323E5",
    x"2362CB3C",
    x"236272B6",
    x"23621A53",
    x"2361C212",
    x"236169F3",
    x"236111F7",
    x"2360BA1D",
    x"23606265",
    x"23600AD0",
    x"235FB35D",
    x"235F5C0C",
    x"235F04DD",
    x"235EADD0",
    x"235E56E5",
    x"235E001C",
    x"235DA975",
    x"235D52F0",
    x"235CFC8C",
    x"235CA64A",
    x"235C502A",
    x"235BFA2C",
    x"235BA44F",
    x"235B4E93",
    x"235AF8F9",
    x"235AA381",
    x"235A4E2A",
    x"2359F8F4",
    x"2359A3DF",
    x"23594EEC",
    x"2358FA1A",
    x"2358A568",
    x"235850D8",
    x"2357FC69",
    x"2357A81B",
    x"235753EE",
    x"2356FFE2",
    x"2356ABF6",
    x"2356582B",
    x"23560481",
    x"2355B0F8",
    x"23555D8F",
    x"23550A47",
    x"2354B71F",
    x"23546417",
    x"23541131",
    x"2353BE6A",
    x"23536BC4",
    x"2353193E",
    x"2352C6D8",
    x"23527492",
    x"2352226D",
    x"2351D068",
    x"23517E82",
    x"23512CBD",
    x"2350DB17",
    x"23508991",
    x"2350382C",
    x"234FE6E6",
    x"234F95BF",
    x"234F44B9",
    x"234EF3D2",
    x"234EA30A",
    x"234E5262",
    x"234E01DA",
    x"234DB171",
    x"234D6127",
    x"234D10FD",
    x"234CC0F2",
    x"234C7106",
    x"234C2139",
    x"234BD18C",
    x"234B81FE",
    x"234B328E",
    x"234AE33E",
    x"234A940D",
    x"234A44FB",
    x"2349F607",
    x"2349A732",
    x"2349587C",
    x"234909E5",
    x"2348BB6D",
    x"23486D13",
    x"23481ED7",
    x"2347D0BB",
    x"234782BC",
    x"234734DC",
    x"2346E71B",
    x"23469978",
    x"23464BF3",
    x"2345FE8D",
    x"2345B144",
    x"2345641A",
    x"2345170E",
    x"2344CA20",
    x"23447D50",
    x"2344309E",
    x"2343E40A",
    x"23439794",
    x"23434B3C",
    x"2342FF01",
    x"2342B2E4",
    x"234266E5",
    x"23421B04",
    x"2341CF40",
    x"2341839A",
    x"23413811",
    x"2340ECA6",
    x"2340A159",
    x"23405628",
    x"23400B15",
    x"233FC01F",
    x"233F7547",
    x"233F2A8C",
    x"233EDFEE",
    x"233E956D",
    x"233E4B09",
    x"233E00C2",
    x"233DB698",
    x"233D6C8C",
    x"233D229C",
    x"233CD8C9",
    x"233C8F12",
    x"233C4579",
    x"233BFBFC",
    x"233BB29C",
    x"233B6958",
    x"233B2032",
    x"233AD727",
    x"233A8E39",
    x"233A4568",
    x"2339FCB3",
    x"2339B41B",
    x"23396B9E",
    x"2339233F",
    x"2338DAFB",
    x"233892D4",
    x"23384AC8",
    x"233802D9",
    x"2337BB06",
    x"2337734F",
    x"23372BB4",
    x"2336E435",
    x"23369CD2",
    x"2336558A",
    x"23360E5F",
    x"2335C74F",
    x"2335805B",
    x"23353983",
    x"2334F2C6",
    x"2334AC25",
    x"233465A0",
    x"23341F36",
    x"2333D8E7",
    x"233392B4",
    x"23334C9D",
    x"233306A0",
    x"2332C0BF",
    x"23327AFA",
    x"2332354F",
    x"2331EFC0",
    x"2331AA4C",
    x"233164F3",
    x"23311FB5",
    x"2330DA92",
    x"2330958A",
    x"2330509D",
    x"23300BCB",
    x"232FC714",
    x"232F8278",
    x"232F3DF6",
    x"232EF98F",
    x"232EB543",
    x"232E7112",
    x"232E2CFB",
    x"232DE8FF",
    x"232DA51D",
    x"232D6156",
    x"232D1DA9",
    x"232CDA16",
    x"232C969E",
    x"232C5341",
    x"232C0FFD",
    x"232BCCD4",
    x"232B89C5",
    x"232B46D1",
    x"232B03F6",
    x"232AC135",
    x"232A7E8F",
    x"232A3C03",
    x"2329F990",
    x"2329B738",
    x"232974F9",
    x"232932D4",
    x"2328F0C9",
    x"2328AED8",
    x"23286D01",
    x"23282B43",
    x"2327E99F",
    x"2327A814",
    x"232766A3",
    x"2327254C",
    x"2326E40E",
    x"2326A2EA",
    x"232661DF",
    x"232620ED",
    x"2325E015",
    x"23259F56",
    x"23255EB1",
    x"23251E24",
    x"2324DDB1",
    x"23249D57",
    x"23245D16",
    x"23241CEE",
    x"2323DCE0",
    x"23239CEA",
    x"23235D0D",
    x"23231D49",
    x"2322DD9E",
    x"23229E0C",
    x"23225E93",
    x"23221F32",
    x"2321DFEA",
    x"2321A0BB",
    x"232161A5",
    x"232122A7",
    x"2320E3C2",
    x"2320A4F5",
    x"23206641",
    x"232027A5",
    x"231FE922",
    x"231FAAB7",
    x"231F6C64",
    x"231F2E2A",
    x"231EF008",
    x"231EB1FF",
    x"231E740D",
    x"231E3634",
    x"231DF873",
    x"231DBACA",
    x"231D7D39",
    x"231D3FC0",
    x"231D025F",
    x"231CC516",
    x"231C87E5",
    x"231C4ACC",
    x"231C0DCB",
    x"231BD0E1",
    x"231B940F",
    x"231B5756",
    x"231B1AB3",
    x"231ADE29",
    x"231AA1B6",
    x"231A655A",
    x"231A2916",
    x"2319ECEA",
    x"2319B0D5",
    x"231974D8",
    x"231938F2",
    x"2318FD24",
    x"2318C16C",
    x"231885CC",
    x"23184A44",
    x"23180ED2",
    x"2317D378",
    x"23179835",
    x"23175D09",
    x"231721F4",
    x"2316E6F7",
    x"2316AC10",
    x"23167140",
    x"23163688",
    x"2315FBE6",
    x"2315C15B",
    x"231586E7",
    x"23154C89",
    x"23151243",
    x"2314D813",
    x"23149DFA",
    x"231463F8",
    x"23142A0C",
    x"2313F037",
    x"2313B678",
    x"23137CD0",
    x"2313433F",
    x"231309C4",
    x"2312D05F",
    x"23129711",
    x"23125DD9",
    x"231224B7",
    x"2311EBAC",
    x"2311B2B7",
    x"231179D9",
    x"23114110",
    x"2311085E",
    x"2310CFC2",
    x"2310973B",
    x"23105ECB",
    x"23102671",
    x"230FEE2D",
    x"230FB5FF",
    x"230F7DE7",
    x"230F45E5",
    x"230F0DF9",
    x"230ED622",
    x"230E9E61",
    x"230E66B6",
    x"230E2F21",
    x"230DF7A1",
    x"230DC038",
    x"230D88E3",
    x"230D51A5",
    x"230D1A7B",
    x"230CE368",
    x"230CAC6A",
    x"230C7581",
    x"230C3EAE",
    x"230C07F0",
    x"230BD148",
    x"230B9AB5",
    x"230B6437",
    x"230B2DCE",
    x"230AF77B",
    x"230AC13D",
    x"230A8B14",
    x"230A5500",
    x"230A1F02",
    x"2309E918",
    x"2309B344",
    x"23097D84",
    x"230947DA",
    x"23091244",
    x"2308DCC3",
    x"2308A757",
    x"23087201",
    x"23083CBE",
    x"23080791",
    x"2307D278",
    x"23079D75",
    x"23076885",
    x"230733AB",
    x"2306FEE5",
    x"2306CA34",
    x"23069597",
    x"2306610F",
    x"23062C9B",
    x"2305F83C",
    x"2305C3F1",
    x"23058FBB",
    x"23055B99",
    x"2305278B",
    x"2304F392",
    x"2304BFAD",
    x"23048BDC",
    x"23045820",
    x"23042477",
    x"2303F0E3",
    x"2303BD63",
    x"230389F7",
    x"2303569F",
    x"2303235C",
    x"2302F02C",
    x"2302BD10",
    x"23028A08",
    x"23025714",
    x"23022434",
    x"2301F168",
    x"2301BEAF",
    x"23018C0B",
    x"2301597A",
    x"230126FD",
    x"2300F494",
    x"2300C23E",
    x"23008FFC",
    x"23005DCD",
    x"23002BB3",
    x"22FFF356",
    x"22FF8F6F",
    x"22FF2BAE",
    x"22FEC815",
    x"22FE64A2",
    x"22FE0156",
    x"22FD9E31",
    x"22FD3B33",
    x"22FCD85B",
    x"22FC75AA",
    x"22FC131F",
    x"22FBB0BB",
    x"22FB4E7D",
    x"22FAEC65",
    x"22FA8A74",
    x"22FA28A9",
    x"22F9C704",
    x"22F96586",
    x"22F9042D",
    x"22F8A2FA",
    x"22F841EE",
    x"22F7E107",
    x"22F78046",
    x"22F71FAA",
    x"22F6BF35",
    x"22F65EE5",
    x"22F5FEBB",
    x"22F59EB6",
    x"22F53ED7",
    x"22F4DF1D",
    x"22F47F88",
    x"22F42019",
    x"22F3C0CF",
    x"22F361AB",
    x"22F302AB",
    x"22F2A3D1",
    x"22F2451B",
    x"22F1E68B",
    x"22F1881F",
    x"22F129D8",
    x"22F0CBB6",
    x"22F06DB9",
    x"22F00FE0",
    x"22EFB22D",
    x"22EF549D",
    x"22EEF732",
    x"22EE99EC",
    x"22EE3CCA",
    x"22EDDFCD",
    x"22ED82F3",
    x"22ED263E",
    x"22ECC9AD",
    x"22EC6D41",
    x"22EC10F8",
    x"22EBB4D3",
    x"22EB58D3",
    x"22EAFCF6",
    x"22EAA13D",
    x"22EA45A8",
    x"22E9EA37",
    x"22E98EE9",
    x"22E933BF",
    x"22E8D8B9",
    x"22E87DD6",
    x"22E82316",
    x"22E7C87A",
    x"22E76E02",
    x"22E713AC",
    x"22E6B97A",
    x"22E65F6B",
    x"22E60580",
    x"22E5ABB7",
    x"22E55212",
    x"22E4F88F",
    x"22E49F2F",
    x"22E445F3",
    x"22E3ECD9",
    x"22E393E2",
    x"22E33B0D",
    x"22E2E25B",
    x"22E289CC",
    x"22E23160",
    x"22E1D916",
    x"22E180EE",
    x"22E128E9",
    x"22E0D106",
    x"22E07946",
    x"22E021A7",
    x"22DFCA2B",
    x"22DF72D1",
    x"22DF1B9A",
    x"22DEC484",
    x"22DE6D90",
    x"22DE16BE",
    x"22DDC00E",
    x"22DD6980",
    x"22DD1314",
    x"22DCBCC9",
    x"22DC66A0",
    x"22DC1099",
    x"22DBBAB3",
    x"22DB64EF",
    x"22DB0F4C",
    x"22DAB9CB",
    x"22DA646B",
    x"22DA0F2D",
    x"22D9BA0F",
    x"22D96513",
    x"22D91038",
    x"22D8BB7F",
    x"22D866E6",
    x"22D8126E",
    x"22D7BE17",
    x"22D769E2",
    x"22D715CD",
    x"22D6C1D9",
    x"22D66E05",
    x"22D61A53",
    x"22D5C6C1",
    x"22D5734F",
    x"22D51FFF",
    x"22D4CCCE",
    x"22D479BF",
    x"22D426CF",
    x"22D3D400",
    x"22D38152",
    x"22D32EC3",
    x"22D2DC55",
    x"22D28A07",
    x"22D237D9",
    x"22D1E5CB",
    x"22D193DE",
    x"22D14210",
    x"22D0F062",
    x"22D09ED4",
    x"22D04D66",
    x"22CFFC18",
    x"22CFAAE9",
    x"22CF59DA",
    x"22CF08EB",
    x"22CEB81B",
    x"22CE676B",
    x"22CE16DA",
    x"22CDC669",
    x"22CD7617",
    x"22CD25E5",
    x"22CCD5D2",
    x"22CC85DE",
    x"22CC3609",
    x"22CBE653",
    x"22CB96BD",
    x"22CB4746",
    x"22CAF7ED",
    x"22CAA8B4",
    x"22CA599A",
    x"22CA0A9E",
    x"22C9BBC1",
    x"22C96D03",
    x"22C91E64",
    x"22C8CFE3",
    x"22C88182",
    x"22C8333E",
    x"22C7E51A",
    x"22C79713",
    x"22C7492C",
    x"22C6FB62",
    x"22C6ADB7",
    x"22C6602A",
    x"22C612BC",
    x"22C5C56C",
    x"22C5783A",
    x"22C52B26",
    x"22C4DE30",
    x"22C49158",
    x"22C4449E",
    x"22C3F803",
    x"22C3AB85",
    x"22C35F25",
    x"22C312E2",
    x"22C2C6BE",
    x"22C27AB7",
    x"22C22ECE",
    x"22C1E302",
    x"22C19755",
    x"22C14BC4",
    x"22C10051",
    x"22C0B4FC",
    x"22C069C4",
    x"22C01EA9",
    x"22BFD3AC",
    x"22BF88CC",
    x"22BF3E09",
    x"22BEF363",
    x"22BEA8DB",
    x"22BE5E6F",
    x"22BE1421",
    x"22BDC9F0",
    x"22BD7FDB",
    x"22BD35E4",
    x"22BCEC09",
    x"22BCA24B",
    x"22BC58AA",
    x"22BC0F26",
    x"22BBC5BF",
    x"22BB7C74",
    x"22BB3345",
    x"22BAEA34",
    x"22BAA13E",
    x"22BA5866",
    x"22BA0FA9",
    x"22B9C709",
    x"22B97E86",
    x"22B9361E",
    x"22B8EDD3",
    x"22B8A5A5",
    x"22B85D92",
    x"22B8159C",
    x"22B7CDC1",
    x"22B78603",
    x"22B73E60",
    x"22B6F6DA",
    x"22B6AF70",
    x"22B66821",
    x"22B620EE",
    x"22B5D9D7",
    x"22B592DC",
    x"22B54BFC",
    x"22B50539",
    x"22B4BE90",
    x"22B47804",
    x"22B43193",
    x"22B3EB3D",
    x"22B3A503",
    x"22B35EE4",
    x"22B318E1",
    x"22B2D2F9",
    x"22B28D2C",
    x"22B2477A",
    x"22B201E4",
    x"22B1BC69",
    x"22B17709",
    x"22B131C4",
    x"22B0EC9A",
    x"22B0A78B",
    x"22B06297",
    x"22B01DBE",
    x"22AFD900",
    x"22AF945C",
    x"22AF4FD4",
    x"22AF0B66",
    x"22AEC713",
    x"22AE82DA",
    x"22AE3EBD",
    x"22ADFAB9",
    x"22ADB6D1",
    x"22AD7303",
    x"22AD2F4F",
    x"22ACEBB6",
    x"22ACA837",
    x"22AC64D2",
    x"22AC2188",
    x"22ABDE58",
    x"22AB9B42",
    x"22AB5847",
    x"22AB1565",
    x"22AAD29E",
    x"22AA8FF1",
    x"22AA4D5D",
    x"22AA0AE4",
    x"22A9C885",
    x"22A98640",
    x"22A94414",
    x"22A90202",
    x"22A8C00A",
    x"22A87E2C",
    x"22A83C68",
    x"22A7FABD",
    x"22A7B92C",
    x"22A777B4",
    x"22A73656",
    x"22A6F512",
    x"22A6B3E7",
    x"22A672D5",
    x"22A631DD",
    x"22A5F0FE",
    x"22A5B039",
    x"22A56F8D",
    x"22A52EFA",
    x"22A4EE80",
    x"22A4AE1F",
    x"22A46DD8",
    x"22A42DAA",
    x"22A3ED94",
    x"22A3AD98",
    x"22A36DB5",
    x"22A32DEA",
    x"22A2EE39",
    x"22A2AEA0",
    x"22A26F20",
    x"22A22FB9",
    x"22A1F06B",
    x"22A1B135",
    x"22A17219",
    x"22A13314",
    x"22A0F429",
    x"22A0B556",
    x"22A0769B",
    x"22A037F9",
    x"229FF96F",
    x"229FBAFE",
    x"229F7CA5",
    x"229F3E65",
    x"229F003C",
    x"229EC22C",
    x"229E8435",
    x"229E4655",
    x"229E088E",
    x"229DCADE",
    x"229D8D47",
    x"229D4FC8",
    x"229D1261",
    x"229CD512",
    x"229C97DA",
    x"229C5ABB",
    x"229C1DB4",
    x"229BE0C4",
    x"229BA3EC",
    x"229B672C",
    x"229B2A83",
    x"229AEDF3",
    x"229AB179",
    x"229A7518",
    x"229A38CE",
    x"2299FC9B",
    x"2299C081",
    x"2299847D",
    x"22994891",
    x"22990CBC",
    x"2298D0FF",
    x"22989559",
    x"229859CA",
    x"22981E53",
    x"2297E2F3",
    x"2297A7AA",
    x"22976C78",
    x"2297315D",
    x"2296F659",
    x"2296BB6C",
    x"22968097",
    x"229645D8",
    x"22960B30",
    x"2295D09F",
    x"22959625",
    x"22955BC2",
    x"22952175",
    x"2294E740",
    x"2294AD21",
    x"22947318",
    x"22943927",
    x"2293FF4C",
    x"2293C587",
    x"22938BD9",
    x"22935242",
    x"229318C1",
    x"2292DF57",
    x"2292A603",
    x"22926CC5",
    x"2292339E",
    x"2291FA8D",
    x"2291C192",
    x"229188AD",
    x"22914FDF",
    x"22911727",
    x"2290DE85",
    x"2290A5F9",
    x"22906D83",
    x"22903524",
    x"228FFCDA",
    x"228FC4A6",
    x"228F8C88",
    x"228F5480",
    x"228F1C8E",
    x"228EE4B2",
    x"228EACEB",
    x"228E753B",
    x"228E3DA0",
    x"228E061B",
    x"228DCEAB",
    x"228D9751",
    x"228D600D",
    x"228D28DE",
    x"228CF1C5",
    x"228CBAC1",
    x"228C83D3",
    x"228C4CFA",
    x"228C1637",
    x"228BDF89",
    x"228BA8F0",
    x"228B726D",
    x"228B3BFF",
    x"228B05A6",
    x"228ACF62",
    x"228A9934",
    x"228A631B",
    x"228A2D17",
    x"2289F727",
    x"2289C14D",
    x"22898B88",
    x"228955D8",
    x"2289203D",
    x"2288EAB7",
    x"2288B546",
    x"22887FEA",
    x"22884AA2",
    x"2288156F",
    x"2287E051",
    x"2287AB48",
    x"22877653",
    x"22874174",
    x"22870CA8",
    x"2286D7F2",
    x"2286A350",
    x"22866EC2",
    x"22863A49",
    x"228605E5",
    x"2285D194",
    x"22859D59",
    x"22856931",
    x"2285351F",
    x"22850120",
    x"2284CD36",
    x"22849960",
    x"2284659E",
    x"228431F0",
    x"2283FE57",
    x"2283CAD2",
    x"22839760",
    x"22836403",
    x"228330BA",
    x"2282FD85",
    x"2282CA64",
    x"22829757",
    x"2282645E",
    x"22823179",
    x"2281FEA7",
    x"2281CBEA",
    x"22819940",
    x"228166AA",
    x"22813428",
    x"228101B9",
    x"2280CF5E",
    x"22809D17",
    x"22806AE4",
    x"228038C4",
    x"228006B7",
    x"227FA97D",
    x"227F45B2",
    x"227EE20E",
    x"227E7E91",
    x"227E1B3B",
    x"227DB80C",
    x"227D5504",
    x"227CF222",
    x"227C8F66",
    x"227C2CD2",
    x"227BCA63",
    x"227B681C",
    x"227B05FA",
    x"227AA3FF",
    x"227A422A",
    x"2279E07B",
    x"22797EF2",
    x"22791D90",
    x"2278BC53",
    x"22785B3D",
    x"2277FA4C",
    x"22779981",
    x"227738DC",
    x"2276D85D",
    x"22767803",
    x"227617CF",
    x"2275B7C0",
    x"227557D7",
    x"2274F814",
    x"22749876",
    x"227438FD",
    x"2273D9A9",
    x"22737A7B",
    x"22731B71",
    x"2272BC8D",
    x"22725DCE",
    x"2271FF34",
    x"2271A0BF",
    x"2271426E",
    x"2270E443",
    x"2270863C",
    x"2270285A",
    x"226FCA9C",
    x"226F6D04",
    x"226F0F8F",
    x"226EB23F",
    x"226E5514",
    x"226DF80D",
    x"226D9B2A",
    x"226D3E6C",
    x"226CE1D1",
    x"226C855B",
    x"226C2909",
    x"226BCCDB",
    x"226B70D1",
    x"226B14EB",
    x"226AB929",
    x"226A5D8A",
    x"226A0210",
    x"2269A6B9",
    x"22694B85",
    x"2268F076",
    x"22689589",
    x"22683AC1",
    x"2267E01C",
    x"2267859A",
    x"22672B3B",
    x"2266D100",
    x"226676E8",
    x"22661CF3",
    x"2265C321",
    x"22656973",
    x"22650FE7",
    x"2264B67E",
    x"22645D38",
    x"22640415",
    x"2263AB15",
    x"22635238",
    x"2262F97D",
    x"2262A0E5",
    x"2262486F",
    x"2261F01C",
    x"226197EB",
    x"22613FDD",
    x"2260E7F2",
    x"22609028",
    x"22603881",
    x"225FE0FC",
    x"225F8999",
    x"225F3258",
    x"225EDB3A",
    x"225E843D",
    x"225E2D62",
    x"225DD6AA",
    x"225D8013",
    x"225D299E",
    x"225CD34A",
    x"225C7D18",
    x"225C2708",
    x"225BD11A",
    x"225B7B4D",
    x"225B25A2",
    x"225AD018",
    x"225A7AAF",
    x"225A2568",
    x"2259D042",
    x"22597B3D",
    x"22592659",
    x"2258D197",
    x"22587CF6",
    x"22582875",
    x"2257D416",
    x"22577FD8",
    x"22572BBA",
    x"2256D7BE",
    x"225683E2",
    x"22563026",
    x"2255DC8C",
    x"22558912",
    x"225535B9",
    x"2254E280",
    x"22548F68",
    x"22543C70",
    x"2253E999",
    x"225396E2",
    x"2253444B",
    x"2252F1D4",
    x"22529F7E",
    x"22524D48",
    x"2251FB31",
    x"2251A93B",
    x"22515765",
    x"225105AF",
    x"2250B419",
    x"225062A2",
    x"2250114C",
    x"224FC015",
    x"224F6EFE",
    x"224F1E06",
    x"224ECD2E",
    x"224E7C76",
    x"224E2BDD",
    x"224DDB64",
    x"224D8B0A",
    x"224D3ACF",
    x"224CEAB4",
    x"224C9AB7",
    x"224C4ADB",
    x"224BFB1D",
    x"224BAB7E",
    x"224B5BFF",
    x"224B0C9F",
    x"224ABD5D",
    x"224A6E3B",
    x"224A1F37",
    x"2249D052",
    x"2249818C",
    x"224932E5",
    x"2248E45C",
    x"224895F3",
    x"224847A7",
    x"2247F97B",
    x"2247AB6C",
    x"22475D7D",
    x"22470FAB",
    x"2246C1F8",
    x"22467464",
    x"224626ED",
    x"2245D995",
    x"22458C5B",
    x"22453F40",
    x"2244F242",
    x"2244A562",
    x"224458A1",
    x"22440BFD",
    x"2243BF77",
    x"22437310",
    x"224326C5",
    x"2242DA99",
    x"22428E8B",
    x"2242429A",
    x"2241F6C7",
    x"2241AB11",
    x"22415F79",
    x"224113FE",
    x"2240C8A1",
    x"22407D62",
    x"2240323F",
    x"223FE73A",
    x"223F9C53",
    x"223F5188",
    x"223F06DB",
    x"223EBC4B",
    x"223E71D8",
    x"223E2782",
    x"223DDD49",
    x"223D932D",
    x"223D492E",
    x"223CFF4C",
    x"223CB587",
    x"223C6BDE",
    x"223C2252",
    x"223BD8E3",
    x"223B8F91",
    x"223B465B",
    x"223AFD42",
    x"223AB445",
    x"223A6B65",
    x"223A22A1",
    x"2239D9FA",
    x"2239916F",
    x"22394900",
    x"223900AE",
    x"2238B878",
    x"2238705E",
    x"22382860",
    x"2237E07E",
    x"223798B9",
    x"2237510F",
    x"22370981",
    x"2236C20F",
    x"22367ABA",
    x"22363380",
    x"2235EC61",
    x"2235A55F",
    x"22355E78",
    x"223517AD",
    x"2234D0FE",
    x"22348A6A",
    x"223443F1",
    x"2233FD95",
    x"2233B753",
    x"2233712D",
    x"22332B23",
    x"2232E534",
    x"22329F60",
    x"223259A7",
    x"2232140A",
    x"2231CE88",
    x"22318920",
    x"223143D4",
    x"2230FEA3",
    x"2230B98D",
    x"22307492",
    x"22302FB2",
    x"222FEAED",
    x"222FA643",
    x"222F61B3",
    x"222F1D3E",
    x"222ED8E4",
    x"222E94A5",
    x"222E5080",
    x"222E0C76",
    x"222DC886",
    x"222D84B1",
    x"222D40F7",
    x"222CFD57",
    x"222CB9D1",
    x"222C7665",
    x"222C3314",
    x"222BEFDE",
    x"222BACC1",
    x"222B69BF",
    x"222B26D6",
    x"222AE408",
    x"222AA154",
    x"222A5EBA",
    x"222A1C3A",
    x"2229D9D4",
    x"22299788",
    x"22295556",
    x"2229133D",
    x"2228D13F",
    x"22288F5A",
    x"22284D8F",
    x"22280BDD",
    x"2227CA45",
    x"222788C7",
    x"22274762",
    x"22270617",
    x"2226C4E6",
    x"222683CE",
    x"222642CF",
    x"222601E9",
    x"2225C11D",
    x"2225806A",
    x"22253FD1",
    x"2224FF51",
    x"2224BEE9",
    x"22247E9B",
    x"22243E66",
    x"2223FE4B",
    x"2223BE48",
    x"22237E5E",
    x"22233E8D",
    x"2222FED5",
    x"2222BF36",
    x"22227FB0",
    x"22224042",
    x"222200ED",
    x"2221C1B1",
    x"2221828E",
    x"22214383",
    x"22210491",
    x"2220C5B8",
    x"222086F7",
    x"2220484E",
    x"222009BE",
    x"221FCB47",
    x"221F8CE8",
    x"221F4EA1",
    x"221F1072",
    x"221ED25C",
    x"221E945E",
    x"221E5678",
    x"221E18AA",
    x"221DDAF5",
    x"221D9D57",
    x"221D5FD2",
    x"221D2264",
    x"221CE50F",
    x"221CA7D1",
    x"221C6AAC",
    x"221C2D9E",
    x"221BF0A8",
    x"221BB3CA",
    x"221B7704",
    x"221B3A55",
    x"221AFDBE",
    x"221AC13F",
    x"221A84D7",
    x"221A4887",
    x"221A0C4E",
    x"2219D02D",
    x"22199424",
    x"22195832",
    x"22191C57",
    x"2218E093",
    x"2218A4E7",
    x"22186953",
    x"22182DD5",
    x"2217F26F",
    x"2217B720",
    x"22177BE8",
    x"221740C7",
    x"221705BD",
    x"2216CACA",
    x"22168FEF",
    x"2216552A",
    x"22161A7C",
    x"2215DFE5",
    x"2215A565",
    x"22156AFC",
    x"221530AA",
    x"2214F66E",
    x"2214BC49",
    x"2214823B",
    x"22144843",
    x"22140E62",
    x"2213D498",
    x"22139AE4",
    x"22136147",
    x"221327C0",
    x"2212EE50",
    x"2212B4F6",
    x"22127BB2",
    x"22124285",
    x"2212096F",
    x"2211D06E",
    x"22119784",
    x"22115EB0",
    x"221125F2",
    x"2210ED4A",
    x"2210B4B8",
    x"22107C3D",
    x"221043D7",
    x"22100B88",
    x"220FD34E",
    x"220F9B2B",
    x"220F631D",
    x"220F2B25",
    x"220EF343",
    x"220EBB77",
    x"220E83C1",
    x"220E4C20",
    x"220E1495",
    x"220DDD20",
    x"220DA5C1",
    x"220D6E77",
    x"220D3742",
    x"220D0023",
    x"220CC91A",
    x"220C9226",
    x"220C5B48",
    x"220C247F",
    x"220BEDCB",
    x"220BB72D",
    x"220B80A4",
    x"220B4A31",
    x"220B13D2",
    x"220ADD89",
    x"220AA755",
    x"220A7136",
    x"220A3B2D",
    x"220A0538",
    x"2209CF59",
    x"2209998E",
    x"220963D9",
    x"22092E38",
    x"2208F8AD",
    x"2208C336",
    x"22088DD4",
    x"22085887",
    x"2208234F",
    x"2207EE2B",
    x"2207B91D",
    x"22078423",
    x"22074F3E",
    x"22071A6D",
    x"2206E5B1",
    x"2206B109",
    x"22067C77",
    x"220647F8",
    x"2206138E",
    x"2205DF39",
    x"2205AAF8",
    x"220576CB",
    x"220542B3",
    x"22050EAF",
    x"2204DAC0",
    x"2204A6E4",
    x"2204731D",
    x"22043F6A",
    x"22040BCC",
    x"2203D841",
    x"2203A4CB",
    x"22037168",
    x"22033E1A",
    x"22030AE0",
    x"2202D7BA",
    x"2202A4A7",
    x"220271A9",
    x"22023EBF",
    x"22020BE8",
    x"2201D925",
    x"2201A676",
    x"220173DB",
    x"22014154",
    x"22010EE0",
    x"2200DC80",
    x"2200AA34",
    x"220077FB",
    x"220045D6",
    x"220013C5",
    x"21FFC38D",
    x"21FF5FB8",
    x"21FEFC0A",
    x"21FE9883",
    x"21FE3523",
    x"21FDD1EA",
    x"21FD6ED7",
    x"21FD0BEB",
    x"21FCA926",
    x"21FC4687",
    x"21FBE40F",
    x"21FB81BD",
    x"21FB1F91",
    x"21FABD8C",
    x"21FA5BAD",
    x"21F9F9F5",
    x"21F99862",
    x"21F936F6",
    x"21F8D5AF",
    x"21F8748F",
    x"21F81394",
    x"21F7B2BF",
    x"21F75210",
    x"21F6F187",
    x"21F69124",
    x"21F630E6",
    x"21F5D0CD",
    x"21F570DB",
    x"21F5110D",
    x"21F4B165",
    x"21F451E3",
    x"21F3F285",
    x"21F3934D",
    x"21F3343A",
    x"21F2D54C",
    x"21F27683",
    x"21F217E0",
    x"21F1B961",
    x"21F15B07",
    x"21F0FCD2",
    x"21F09EC1",
    x"21F040D6",
    x"21EFE30F",
    x"21EF856C",
    x"21EF27EE",
    x"21EECA95",
    x"21EE6D60",
    x"21EE1050",
    x"21EDB363",
    x"21ED569B",
    x"21ECF9F8",
    x"21EC9D78",
    x"21EC411D",
    x"21EBE4E5",
    x"21EB88D2",
    x"21EB2CE2",
    x"21EAD117",
    x"21EA756F",
    x"21EA19EB",
    x"21E9BE8B",
    x"21E9634E",
    x"21E90835",
    x"21E8AD40",
    x"21E8526E",
    x"21E7F7BF",
    x"21E79D34",
    x"21E742CC",
    x"21E6E888",
    x"21E68E67",
    x"21E63469",
    x"21E5DA8E",
    x"21E580D6",
    x"21E52741",
    x"21E4CDCF",
    x"21E47480",
    x"21E41B54",
    x"21E3C24B",
    x"21E36964",
    x"21E310A1",
    x"21E2B7FF",
    x"21E25F81",
    x"21E20725",
    x"21E1AEEB",
    x"21E156D4",
    x"21E0FEDF",
    x"21E0A70D",
    x"21E04F5D",
    x"21DFF7CF",
    x"21DFA063",
    x"21DF491A",
    x"21DEF1F2",
    x"21DE9AED",
    x"21DE4409",
    x"21DDED47",
    x"21DD96A8",
    x"21DD402A",
    x"21DCE9CD",
    x"21DC9393",
    x"21DC3D7A",
    x"21DBE783",
    x"21DB91AD",
    x"21DB3BF9",
    x"21DAE666",
    x"21DA90F5",
    x"21DA3BA5",
    x"21D9E676",
    x"21D99169",
    x"21D93C7D",
    x"21D8E7B2",
    x"21D89308",
    x"21D83E7F",
    x"21D7EA17",
    x"21D795D0",
    x"21D741AA",
    x"21D6EDA5",
    x"21D699C0",
    x"21D645FD",
    x"21D5F25A",
    x"21D59ED7",
    x"21D54B75",
    x"21D4F834",
    x"21D4A514",
    x"21D45213",
    x"21D3FF33",
    x"21D3AC74",
    x"21D359D5",
    x"21D30756",
    x"21D2B4F7",
    x"21D262B8",
    x"21D2109A",
    x"21D1BE9B",
    x"21D16CBD",
    x"21D11AFE",
    x"21D0C960",
    x"21D077E1",
    x"21D02682",
    x"21CFD543",
    x"21CF8423",
    x"21CF3324",
    x"21CEE243",
    x"21CE9183",
    x"21CE40E2",
    x"21CDF060",
    x"21CD9FFE",
    x"21CD4FBB",
    x"21CCFF98",
    x"21CCAF93",
    x"21CC5FAE",
    x"21CC0FE9",
    x"21CBC042",
    x"21CB70BA",
    x"21CB2152",
    x"21CAD208",
    x"21CA82DE",
    x"21CA33D2",
    x"21C9E4E5",
    x"21C99617",
    x"21C94768",
    x"21C8F8D7",
    x"21C8AA66",
    x"21C85C12",
    x"21C80DDE",
    x"21C7BFC8",
    x"21C771D0",
    x"21C723F7",
    x"21C6D63C",
    x"21C6889F",
    x"21C63B21",
    x"21C5EDC1",
    x"21C5A07F",
    x"21C5535C",
    x"21C50656",
    x"21C4B96F",
    x"21C46CA5",
    x"21C41FFA",
    x"21C3D36C",
    x"21C386FD",
    x"21C33AAB",
    x"21C2EE77",
    x"21C2A260",
    x"21C25668",
    x"21C20A8D",
    x"21C1BED0",
    x"21C17330",
    x"21C127AE",
    x"21C0DC49",
    x"21C09101",
    x"21C045D7",
    x"21BFFACB",
    x"21BFAFDC",
    x"21BF6509",
    x"21BF1A55",
    x"21BECFBD",
    x"21BE8542",
    x"21BE3AE5",
    x"21BDF0A4",
    x"21BDA681",
    x"21BD5C7A",
    x"21BD1290",
    x"21BCC8C4",
    x"21BC7F14",
    x"21BC3580",
    x"21BBEC0A",
    x"21BBA2B0",
    x"21BB5973",
    x"21BB1052",
    x"21BAC74E",
    x"21BA7E66",
    x"21BA359B",
    x"21B9ECEC",
    x"21B9A45A",
    x"21B95BE4",
    x"21B9138A",
    x"21B8CB4D",
    x"21B8832B",
    x"21B83B26",
    x"21B7F33D",
    x"21B7AB70",
    x"21B763BF",
    x"21B71C2A",
    x"21B6D4B1",
    x"21B68D54",
    x"21B64613",
    x"21B5FEED",
    x"21B5B7E4",
    x"21B570F6",
    x"21B52A23",
    x"21B4E36D",
    x"21B49CD2",
    x"21B45652",
    x"21B40FEE",
    x"21B3C9A6",
    x"21B38379",
    x"21B33D67",
    x"21B2F771",
    x"21B2B196",
    x"21B26BD6",
    x"21B22631",
    x"21B1E0A8",
    x"21B19B3A",
    x"21B155E7",
    x"21B110AF",
    x"21B0CB92",
    x"21B08690",
    x"21B041A9",
    x"21AFFCDC",
    x"21AFB82B",
    x"21AF7394",
    x"21AF2F19",
    x"21AEEAB8",
    x"21AEA671",
    x"21AE6246",
    x"21AE1E35",
    x"21ADDA3E",
    x"21AD9662",
    x"21AD52A1",
    x"21AD0EF9",
    x"21ACCB6D",
    x"21AC87FB",
    x"21AC44A3",
    x"21AC0165",
    x"21ABBE41",
    x"21AB7B38",
    x"21AB3849",
    x"21AAF574",
    x"21AAB2B9",
    x"21AA7019",
    x"21AA2D92",
    x"21A9EB25",
    x"21A9A8D2",
    x"21A96699",
    x"21A9247A",
    x"21A8E275",
    x"21A8A089",
    x"21A85EB7",
    x"21A81CFF",
    x"21A7DB60",
    x"21A799DC",
    x"21A75870",
    x"21A7171E",
    x"21A6D5E6",
    x"21A694C7",
    x"21A653C2",
    x"21A612D6",
    x"21A5D203",
    x"21A5914A",
    x"21A550AA",
    x"21A51023",
    x"21A4CFB5",
    x"21A48F61",
    x"21A44F25",
    x"21A40F03",
    x"21A3CEF9",
    x"21A38F09",
    x"21A34F32",
    x"21A30F73",
    x"21A2CFCD",
    x"21A29041",
    x"21A250CD",
    x"21A21172",
    x"21A1D22F",
    x"21A19305",
    x"21A153F4",
    x"21A114FC",
    x"21A0D61C",
    x"21A09754",
    x"21A058A6",
    x"21A01A0F",
    x"219FDB91",
    x"219F9D2C",
    x"219F5EDE",
    x"219F20AA",
    x"219EE28D",
    x"219EA489",
    x"219E669C",
    x"219E28C8",
    x"219DEB0C",
    x"219DAD69",
    x"219D6FDD",
    x"219D3269",
    x"219CF50E",
    x"219CB7CA",
    x"219C7A9E",
    x"219C3D8A",
    x"219C008E",
    x"219BC3AA",
    x"219B86DD",
    x"219B4A28",
    x"219B0D8B",
    x"219AD106",
    x"219A9498",
    x"219A5842",
    x"219A1C03",
    x"2199DFDC",
    x"2199A3CC",
    x"219967D4",
    x"21992BF3",
    x"2198F029",
    x"2198B477",
    x"219878DC",
    x"21983D59",
    x"219801EC",
    x"2197C697",
    x"21978B59",
    x"21975032",
    x"21971523",
    x"2196DA2A",
    x"21969F48",
    x"2196647D",
    x"219629CA",
    x"2195EF2D",
    x"2195B4A7",
    x"21957A38",
    x"21953FDF",
    x"2195059E",
    x"2194CB73",
    x"2194915F",
    x"21945761",
    x"21941D7A",
    x"2193E3AA",
    x"2193A9F1",
    x"2193704D",
    x"219336C1",
    x"2192FD4B",
    x"2192C3EB",
    x"21928AA2",
    x"2192516F",
    x"21921852",
    x"2191DF4C",
    x"2191A65B",
    x"21916D82",
    x"219134BE",
    x"2190FC10",
    x"2190C379",
    x"21908AF8",
    x"2190528C",
    x"21901A37",
    x"218FE1F8",
    x"218FA9CF",
    x"218F71BB",
    x"218F39BE",
    x"218F01D6",
    x"218ECA04",
    x"218E9248",
    x"218E5AA2",
    x"218E2311",
    x"218DEB97",
    x"218DB431",
    x"218D7CE2",
    x"218D45A8",
    x"218D0E83",
    x"218CD774",
    x"218CA07B",
    x"218C6997",
    x"218C32C9",
    x"218BFC0F",
    x"218BC56C",
    x"218B8EDD",
    x"218B5864",
    x"218B2200",
    x"218AEBB1",
    x"218AB578",
    x"218A7F54",
    x"218A4944",
    x"218A134A",
    x"2189DD65",
    x"2189A795",
    x"218971DA",
    x"21893C34",
    x"218906A3",
    x"2188D127",
    x"21889BC0",
    x"2188666E",
    x"21883130",
    x"2187FC07",
    x"2187C6F3",
    x"218791F4",
    x"21875D09",
    x"21872833",
    x"2186F372",
    x"2186BEC5",
    x"21868A2D",
    x"218655A9",
    x"2186213A",
    x"2185ECDF",
    x"2185B899",
    x"21858467",
    x"21855049",
    x"21851C40",
    x"2184E84B",
    x"2184B46A",
    x"2184809E",
    x"21844CE6",
    x"21841942",
    x"2183E5B2",
    x"2183B236",
    x"21837ECF",
    x"21834B7B",
    x"2183183C",
    x"2182E510",
    x"2182B1F9",
    x"21827EF5",
    x"21824C06",
    x"2182192A",
    x"2181E662",
    x"2181B3AE",
    x"2181810E",
    x"21814E81",
    x"21811C08",
    x"2180E9A3",
    x"2180B752",
    x"21808514",
    x"218052EA",
    x"218020D3",
    x"217FDDA0",
    x"217F79C1",
    x"217F1609",
    x"217EB278",
    x"217E4F0E",
    x"217DEBCA",
    x"217D88AE",
    x"217D25B8",
    x"217CC2E8",
    x"217C603F",
    x"217BFDBD",
    x"217B9B61",
    x"217B392B",
    x"217AD71C",
    x"217A7533",
    x"217A1371",
    x"2179B1D4",
    x"2179505E",
    x"2178EF0D",
    x"21788DE3",
    x"21782CDF",
    x"2177CC00",
    x"21776B47",
    x"21770AB4",
    x"2176AA47",
    x"217649FF",
    x"2175E9DD",
    x"217589E0",
    x"21752A09",
    x"2174CA57",
    x"21746ACB",
    x"21740B64",
    x"2173AC22",
    x"21734D05",
    x"2172EE0E",
    x"21728F3B",
    x"2172308E",
    x"2171D206",
    x"217173A2",
    x"21711563",
    x"2170B749",
    x"21705954",
    x"216FFB83",
    x"216F9DD7",
    x"216F4050",
    x"216EE2ED",
    x"216E85AF",
    x"216E2895",
    x"216DCB9F",
    x"216D6ECE",
    x"216D1220",
    x"216CB597",
    x"216C5933",
    x"216BFCF2",
    x"216BA0D5",
    x"216B44DC",
    x"216AE907",
    x"216A8D56",
    x"216A31C9",
    x"2169D65F",
    x"21697B19",
    x"21691FF7",
    x"2168C4F8",
    x"21686A1D",
    x"21680F65",
    x"2167B4D1",
    x"21675A60",
    x"21670012",
    x"2166A5E8",
    x"21664BE1",
    x"2165F1FD",
    x"2165983C",
    x"21653E9E",
    x"2164E523",
    x"21648BCB",
    x"21643295",
    x"2163D983",
    x"21638094",
    x"216327C7",
    x"2162CF1C",
    x"21627695",
    x"21621E30",
    x"2161C5ED",
    x"21616DCD",
    x"216115CF",
    x"2160BDF4",
    x"2160663B",
    x"21600EA4",
    x"215FB730",
    x"215F5FDD",
    x"215F08AD",
    x"215EB19E",
    x"215E5AB2",
    x"215E03E7",
    x"215DAD3F",
    x"215D56B8",
    x"215D0053",
    x"215CAA10",
    x"215C53EE",
    x"215BFDEE",
    x"215BA810",
    x"215B5253",
    x"215AFCB7",
    x"215AA73D",
    x"215A51E5",
    x"2159FCAD",
    x"2159A797",
    x"215952A2",
    x"2158FDCF",
    x"2158A91C",
    x"2158548B",
    x"2158001A",
    x"2157ABCB",
    x"2157579C",
    x"2157038E",
    x"2156AFA1",
    x"21565BD5",
    x"21560829",
    x"2155B49E",
    x"21556134",
    x"21550DEA",
    x"2154BAC1",
    x"215467B9",
    x"215414D0",
    x"2153C208",
    x"21536F61",
    x"21531CD9",
    x"2152CA72",
    x"2152782B",
    x"21522604",
    x"2151D3FD",
    x"21518217",
    x"21513050",
    x"2150DEA9",
    x"21508D22",
    x"21503BBB",
    x"214FEA73",
    x"214F994B",
    x"214F4843",
    x"214EF75B",
    x"214EA692",
    x"214E55E9",
    x"214E055F",
    x"214DB4F5",
    x"214D64AA",
    x"214D147E",
    x"214CC471",
    x"214C7484",
    x"214C24B6",
    x"214BD508",
    x"214B8578",
    x"214B3607",
    x"214AE6B6",
    x"214A9783",
    x"214A486F",
    x"2149F97B",
    x"2149AAA4",
    x"21495BED",
    x"21490D55",
    x"2148BEDB",
    x"21487080",
    x"21482243",
    x"2147D425",
    x"21478625",
    x"21473844",
    x"2146EA81",
    x"21469CDD",
    x"21464F57",
    x"214601EF",
    x"2145B4A5",
    x"2145677A",
    x"21451A6C",
    x"2144CD7D",
    x"214480AC",
    x"214433F8",
    x"2143E763",
    x"21439AEC",
    x"21434E92",
    x"21430256",
    x"2142B638",
    x"21426A38",
    x"21421E55",
    x"2141D290",
    x"214186E9",
    x"21413B5F",
    x"2140EFF2",
    x"2140A4A3",
    x"21405972",
    x"21400E5D",
    x"213FC366",
    x"213F788D",
    x"213F2DD0",
    x"213EE331",
    x"213E98AF",
    x"213E4E4A",
    x"213E0401",
    x"213DB9D6",
    x"213D6FC8",
    x"213D25D7",
    x"213CDC03",
    x"213C924B",
    x"213C48B0",
    x"213BFF32",
    x"213BB5D1",
    x"213B6C8C",
    x"213B2364",
    x"213ADA59",
    x"213A916A",
    x"213A4897",
    x"2139FFE1",
    x"2139B747",
    x"21396ECA",
    x"21392669",
    x"2138DE24",
    x"213895FB",
    x"21384DEE",
    x"213805FE",
    x"2137BE2A",
    x"21377671",
    x"21372ED5",
    x"2136E755",
    x"21369FF0",
    x"213658A8",
    x"2136117B",
    x"2135CA6A",
    x"21358375",
    x"21353C9C",
    x"2134F5DE",
    x"2134AF3B",
    x"213468B5",
    x"2134224A",
    x"2133DBFA",
    x"213395C6",
    x"21334FAD",
    x"213309AF",
    x"2132C3CD",
    x"21327E06",
    x"2132385B",
    x"2131F2CA",
    x"2131AD55",
    x"213167FB",
    x"213122BC",
    x"2130DD98",
    x"2130988F",
    x"213053A1",
    x"21300ECD",
    x"212FCA15",
    x"212F8578",
    x"212F40F5",
    x"212EFC8D",
    x"212EB83F",
    x"212E740D",
    x"212E2FF5",
    x"212DEBF7",
    x"212DA814",
    x"212D644C",
    x"212D209E",
    x"212CDD0B",
    x"212C9991",
    x"212C5633",
    x"212C12EE",
    x"212BCFC4",
    x"212B8CB4",
    x"212B49BE",
    x"212B06E2",
    x"212AC420",
    x"212A8179",
    x"212A3EEB",
    x"2129FC78",
    x"2129BA1E",
    x"212977DE",
    x"212935B8",
    x"2128F3AC",
    x"2128B1BA",
    x"21286FE1",
    x"21282E23",
    x"2127EC7D",
    x"2127AAF2",
    x"21276980",
    x"21272827",
    x"2126E6E8",
    x"2126A5C3",
    x"212664B7",
    x"212623C4",
    x"2125E2EB",
    x"2125A22B",
    x"21256184",
    x"212520F7",
    x"2124E082",
    x"2124A027",
    x"21245FE5",
    x"21241FBC",
    x"2123DFAD",
    x"21239FB6",
    x"21235FD8",
    x"21232013",
    x"2122E067",
    x"2122A0D3",
    x"21226159",
    x"212221F7",
    x"2121E2AE",
    x"2121A37E",
    x"21216467",
    x"21212568",
    x"2120E681",
    x"2120A7B4",
    x"212068FE",
    x"21202A62",
    x"211FEBDD",
    x"211FAD71",
    x"211F6F1E",
    x"211F30E3",
    x"211EF2C0",
    x"211EB4B5",
    x"211E76C2",
    x"211E38E8",
    x"211DFB26",
    x"211DBD7C",
    x"211D7FEA",
    x"211D4270",
    x"211D050E",
    x"211CC7C4",
    x"211C8A92",
    x"211C4D78",
    x"211C1075",
    x"211BD38B",
    x"211B96B8",
    x"211B59FD",
    x"211B1D5A",
    x"211AE0CE",
    x"211AA45A",
    x"211A67FE",
    x"211A2BB9",
    x"2119EF8C",
    x"2119B376",
    x"21197777",
    x"21193B90",
    x"2118FFC1",
    x"2118C409",
    x"21188868",
    x"21184CDE",
    x"2118116C",
    x"2117D610",
    x"21179ACC",
    x"21175F9F",
    x"2117248A",
    x"2116E98B",
    x"2116AEA3",
    x"211673D2",
    x"21163919",
    x"2115FE76",
    x"2115C3EA",
    x"21158975",
    x"21154F16",
    x"211514CF",
    x"2114DA9E",
    x"2114A084",
    x"21146681",
    x"21142C94",
    x"2113F2BE",
    x"2113B8FE",
    x"21137F55",
    x"211345C3",
    x"21130C47",
    x"2112D2E1",
    x"21129992",
    x"21126059",
    x"21122737",
    x"2111EE2B",
    x"2111B535",
    x"21117C55",
    x"2111438C",
    x"21110AD8",
    x"2110D23B",
    x"211099B4",
    x"21106143",
    x"211028E8",
    x"210FF0A3",
    x"210FB874",
    x"210F805B",
    x"210F4858",
    x"210F106A",
    x"210ED893",
    x"210EA0D1",
    x"210E6925",
    x"210E318F",
    x"210DFA0F",
    x"210DC2A4",
    x"210D8B4E",
    x"210D540F",
    x"210D1CE5",
    x"210CE5D0",
    x"210CAED1",
    x"210C77E8",
    x"210C4114",
    x"210C0A55",
    x"210BD3AB",
    x"210B9D17",
    x"210B6699",
    x"210B302F",
    x"210AF9DB",
    x"210AC39C",
    x"210A8D72",
    x"210A575E",
    x"210A215E",
    x"2109EB73",
    x"2109B59E",
    x"21097FDE",
    x"21094A32",
    x"2109149C",
    x"2108DF1A",
    x"2108A9AD",
    x"21087455",
    x"21083F12",
    x"210809E4",
    x"2107D4CB",
    x"21079FC6",
    x"21076AD6",
    x"210735FA",
    x"21070134",
    x"2106CC81",
    x"210697E4",
    x"2106635B",
    x"21062EE6",
    x"2105FA86",
    x"2105C63A",
    x"21059203",
    x"21055DE0",
    x"210529D2",
    x"2104F5D8",
    x"2104C1F2",
    x"21048E20",
    x"21045A63",
    x"210426BA",
    x"2103F325",
    x"2103BFA4",
    x"21038C37",
    x"210358DE",
    x"21032599",
    x"2102F269",
    x"2102BF4C",
    x"21028C43",
    x"2102594E",
    x"2102266D",
    x"2101F3A0",
    x"2101C0E7",
    x"21018E42",
    x"21015BB0",
    x"21012932",
    x"2100F6C8",
    x"2100C471",
    x"2100922E",
    x"21005FFF",
    x"21002DE3",
    x"20FFF7B6",
    x"20FF93CD",
    x"20FF300B",
    x"20FECC6F",
    x"20FE68FB",
    x"20FE05AD",
    x"20FDA287",
    x"20FD3F86",
    x"20FCDCAD",
    x"20FC79FA",
    x"20FC176E",
    x"20FBB508",
    x"20FB52C8",
    x"20FAF0AF",
    x"20FA8EBC",
    x"20FA2CEF",
    x"20F9CB49",
    x"20F969C9",
    x"20F9086E",
    x"20F8A73A",
    x"20F8462C",
    x"20F7E543",
    x"20F78480",
    x"20F723E4",
    x"20F6C36C",
    x"20F6631B",
    x"20F602EF",
    x"20F5A2E9",
    x"20F54308",
    x"20F4E34C",
    x"20F483B6",
    x"20F42445",
    x"20F3C4FA",
    x"20F365D3",
    x"20F306D2",
    x"20F2A7F6",
    x"20F2493F",
    x"20F1EAAD",
    x"20F18C40",
    x"20F12DF7",
    x"20F0CFD4",
    x"20F071D5",
    x"20F013FB",
    x"20EFB645",
    x"20EF58B4",
    x"20EEFB48",
    x"20EE9E00",
    x"20EE40DC",
    x"20EDE3DD",
    x"20ED8702",
    x"20ED2A4C",
    x"20ECCDB9",
    x"20EC714B",
    x"20EC1501",
    x"20EBB8DB",
    x"20EB5CD8",
    x"20EB00FA",
    x"20EAA540",
    x"20EA49A9",
    x"20E9EE36",
    x"20E992E7",
    x"20E937BB",
    x"20E8DCB3",
    x"20E881CF",
    x"20E8270E",
    x"20E7CC70",
    x"20E771F6",
    x"20E7179F",
    x"20E6BD6C",
    x"20E6635B",
    x"20E6096E",
    x"20E5AFA4",
    x"20E555FD",
    x"20E4FC79",
    x"20E4A317",
    x"20E449D9",
    x"20E3F0BE",
    x"20E397C5",
    x"20E33EEF",
    x"20E2E63C",
    x"20E28DAB",
    x"20E2353D",
    x"20E1DCF2",
    x"20E184C9",
    x"20E12CC2",
    x"20E0D4DE",
    x"20E07D1C",
    x"20E0257C",
    x"20DFCDFE",
    x"20DF76A3",
    x"20DF1F6A",
    x"20DEC852",
    x"20DE715D",
    x"20DE1A8A",
    x"20DDC3D8",
    x"20DD6D49",
    x"20DD16DB",
    x"20DCC08F",
    x"20DC6A64",
    x"20DC145C",
    x"20DBBE75",
    x"20DB68AF",
    x"20DB130B",
    x"20DABD88",
    x"20DA6827",
    x"20DA12E7",
    x"20D9BDC8",
    x"20D968CA",
    x"20D913EE",
    x"20D8BF33",
    x"20D86A99",
    x"20D8161F",
    x"20D7C1C7",
    x"20D76D90",
    x"20D7197A",
    x"20D6C584",
    x"20D671AF",
    x"20D61DFB",
    x"20D5CA68",
    x"20D576F5",
    x"20D523A3",
    x"20D4D071",
    x"20D47D60",
    x"20D42A6F",
    x"20D3D79F",
    x"20D384EF",
    x"20D3325F",
    x"20D2DFEF",
    x"20D28DA0",
    x"20D23B71",
    x"20D1E962",
    x"20D19772",
    x"20D145A3",
    x"20D0F3F4",
    x"20D0A265",
    x"20D050F5",
    x"20CFFFA5",
    x"20CFAE75",
    x"20CF5D65",
    x"20CF0C74",
    x"20CEBBA3",
    x"20CE6AF2",
    x"20CE1A60",
    x"20CDC9ED",
    x"20CD799A",
    x"20CD2966",
    x"20CCD952",
    x"20CC895C",
    x"20CC3986",
    x"20CBE9CF",
    x"20CB9A38",
    x"20CB4ABF",
    x"20CAFB65",
    x"20CAAC2B",
    x"20CA5D0F",
    x"20CA0E12",
    x"20C9BF34",
    x"20C97074",
    x"20C921D4",
    x"20C8D352",
    x"20C884EF",
    x"20C836AA",
    x"20C7E884",
    x"20C79A7C",
    x"20C74C93",
    x"20C6FEC9",
    x"20C6B11C",
    x"20C6638E",
    x"20C6161E",
    x"20C5C8CD",
    x"20C57B9A",
    x"20C52E84",
    x"20C4E18D",
    x"20C494B4",
    x"20C447F9",
    x"20C3FB5C",
    x"20C3AEDD",
    x"20C3627B",
    x"20C31638",
    x"20C2CA12",
    x"20C27E0A",
    x"20C2321F",
    x"20C1E653",
    x"20C19AA3",
    x"20C14F12",
    x"20C1039E",
    x"20C0B847",
    x"20C06D0E",
    x"20C021F2",
    x"20BFD6F3",
    x"20BF8C12",
    x"20BF414E",
    x"20BEF6A7",
    x"20BEAC1D",
    x"20BE61B0",
    x"20BE1761",
    x"20BDCD2E",
    x"20BD8318",
    x"20BD3920",
    x"20BCEF44",
    x"20BCA585",
    x"20BC5BE2",
    x"20BC125D",
    x"20BBC8F4",
    x"20BB7FA8",
    x"20BB3678",
    x"20BAED65",
    x"20BAA46F",
    x"20BA5B95",
    x"20BA12D7",
    x"20B9CA36",
    x"20B981B1",
    x"20B93949",
    x"20B8F0FC",
    x"20B8A8CC",
    x"20B860B9",
    x"20B818C1",
    x"20B7D0E5",
    x"20B78926",
    x"20B74182",
    x"20B6F9FA",
    x"20B6B28F",
    x"20B66B3F",
    x"20B6240B",
    x"20B5DCF3",
    x"20B595F6",
    x"20B54F16",
    x"20B50851",
    x"20B4C1A7",
    x"20B47B19",
    x"20B434A7",
    x"20B3EE50",
    x"20B3A815",
    x"20B361F5",
    x"20B31BF0",
    x"20B2D607",
    x"20B29039",
    x"20B24A86",
    x"20B204EF",
    x"20B1BF72",
    x"20B17A11",
    x"20B134CB",
    x"20B0EFA0",
    x"20B0AA90",
    x"20B0659B",
    x"20B020C0",
    x"20AFDC01",
    x"20AF975C",
    x"20AF52D3",
    x"20AF0E64",
    x"20AECA0F",
    x"20AE85D6",
    x"20AE41B7",
    x"20ADFDB3",
    x"20ADB9C9",
    x"20AD75F9",
    x"20AD3244",
    x"20ACEEAA",
    x"20ACAB2A",
    x"20AC67C4",
    x"20AC2479",
    x"20ABE148",
    x"20AB9E31",
    x"20AB5B34",
    x"20AB1852",
    x"20AAD589",
    x"20AA92DB",
    x"20AA5046",
    x"20AA0DCC",
    x"20A9CB6C",
    x"20A98925",
    x"20A946F9",
    x"20A904E6",
    x"20A8C2ED",
    x"20A8810D",
    x"20A83F48",
    x"20A7FD9C",
    x"20A7BC0A",
    x"20A77A91",
    x"20A73932",
    x"20A6F7EC",
    x"20A6B6C0",
    x"20A675AE",
    x"20A634B4",
    x"20A5F3D4",
    x"20A5B30E",
    x"20A57260",
    x"20A531CC",
    x"20A4F152",
    x"20A4B0F0",
    x"20A470A7",
    x"20A43078",
    x"20A3F061",
    x"20A3B064",
    x"20A37080",
    x"20A330B4",
    x"20A2F102",
    x"20A2B168",
    x"20A271E7",
    x"20A2327F",
    x"20A1F32F",
    x"20A1B3F9",
    x"20A174DB",
    x"20A135D6",
    x"20A0F6E9",
    x"20A0B815",
    x"20A07959",
    x"20A03AB6",
    x"209FFC2B",
    x"209FBDB9",
    x"209F7F5F",
    x"209F411D",
    x"209F02F4",
    x"209EC4E3",
    x"209E86EA",
    x"209E490A",
    x"209E0B41",
    x"209DCD91",
    x"209D8FF8",
    x"209D5278",
    x"209D1510",
    x"209CD7C0",
    x"209C9A87",
    x"209C5D67",
    x"209C205E",
    x"209BE36E",
    x"209BA695",
    x"209B69D4",
    x"209B2D2A",
    x"209AF098",
    x"209AB41E",
    x"209A77BC",
    x"209A3B71",
    x"2099FF3D",
    x"2099C321",
    x"2099871D",
    x"20994B30",
    x"20990F5A",
    x"2098D39C",
    x"209897F5",
    x"20985C65",
    x"209820EC",
    x"2097E58B",
    x"2097AA41",
    x"20976F0E",
    x"209733F2",
    x"2096F8ED",
    x"2096BE00",
    x"20968329",
    x"20964869",
    x"20960DC0",
    x"2095D32F",
    x"209598B3",
    x"20955E4F",
    x"20952402",
    x"2094E9CB",
    x"2094AFAB",
    x"209475A2",
    x"20943BAF",
    x"209401D3",
    x"2093C80E",
    x"20938E5F",
    x"209354C7",
    x"20931B45",
    x"2092E1D9",
    x"2092A884",
    x"20926F46",
    x"2092361D",
    x"2091FD0B",
    x"2091C410",
    x"20918B2A",
    x"2091525B",
    x"209119A2",
    x"2090E0FF",
    x"2090A872",
    x"20906FFB",
    x"2090379A",
    x"208FFF50",
    x"208FC71B",
    x"208F8EFC",
    x"208F56F3",
    x"208F1F00",
    x"208EE723",
    x"208EAF5C",
    x"208E77AA",
    x"208E400E",
    x"208E0888",
    x"208DD117",
    x"208D99BD",
    x"208D6277",
    x"208D2B48",
    x"208CF42E",
    x"208CBD29",
    x"208C863A",
    x"208C4F60",
    x"208C189C",
    x"208BE1ED",
    x"208BAB53",
    x"208B74CF",
    x"208B3E60",
    x"208B0806",
    x"208AD1C2",
    x"208A9B92",
    x"208A6578",
    x"208A2F73",
    x"2089F983",
    x"2089C3A8",
    x"20898DE2",
    x"20895831",
    x"20892295",
    x"2088ED0E",
    x"2088B79C",
    x"2088823F",
    x"20884CF6",
    x"208817C3",
    x"2087E2A4",
    x"2087AD9A",
    x"208778A4",
    x"208743C3",
    x"20870EF7",
    x"2086DA40",
    x"2086A59D",
    x"2086710E",
    x"20863C94",
    x"2086082F",
    x"2085D3DE",
    x"20859FA1",
    x"20856B79",
    x"20853765",
    x"20850366",
    x"2084CF7B",
    x"20849BA4",
    x"208467E1",
    x"20843433",
    x"20840098",
    x"2083CD12",
    x"208399A0",
    x"20836642",
    x"208332F8",
    x"2082FFC2",
    x"2082CCA0",
    x"20829992",
    x"20826698",
    x"208233B2",
    x"208200E0",
    x"2081CE21",
    x"20819B77",
    x"208168E0",
    x"2081365D",
    x"208103EE",
    x"2080D192",
    x"20809F4A",
    x"20806D15",
    x"20803AF5",
    x"208008E7",
    x"207FADDB",
    x"207F4A0F",
    x"207EE669",
    x"207E82EB",
    x"207E1F93",
    x"207DBC62",
    x"207D5958",
    x"207CF674",
    x"207C93B7",
    x"207C3121",
    x"207BCEB1",
    x"207B6C67",
    x"207B0A44",
    x"207AA847",
    x"207A4671",
    x"2079E4C0",
    x"20798336",
    x"207921D2",
    x"2078C094",
    x"20785F7B",
    x"2077FE89",
    x"20779DBC",
    x"20773D16",
    x"2076DC95",
    x"20767C39",
    x"20761C04",
    x"2075BBF3",
    x"20755C09",
    x"2074FC43",
    x"20749CA4",
    x"20743D29",
    x"2073DDD4",
    x"20737EA4",
    x"20731F99",
    x"2072C0B3",
    x"207261F2",
    x"20720357",
    x"2071A4E0",
    x"2071468E",
    x"2070E861",
    x"20708A58",
    x"20702C74",
    x"206FCEB5",
    x"206F711B",
    x"206F13A5",
    x"206EB654",
    x"206E5927",
    x"206DFC1E",
    x"206D9F3A",
    x"206D4279",
    x"206CE5DE",
    x"206C8966",
    x"206C2D12",
    x"206BD0E3",
    x"206B74D7",
    x"206B18EF",
    x"206ABD2C",
    x"206A618C",
    x"206A060F",
    x"2069AAB7",
    x"20694F82",
    x"2068F471",
    x"20689983",
    x"20683EB9",
    x"2067E412",
    x"2067898E",
    x"20672F2E",
    x"2066D4F2",
    x"20667AD8",
    x"206620E2",
    x"2065C70E",
    x"20656D5E",
    x"206513D1",
    x"2064BA67",
    x"2064611F",
    x"206407FB",
    x"2063AEF9",
    x"2063561A",
    x"2062FD5E",
    x"2062A4C4",
    x"20624C4D",
    x"2061F3F8",
    x"20619BC6",
    x"206143B7",
    x"2060EBC9",
    x"206093FE",
    x"20603C56",
    x"205FE4CF",
    x"205F8D6B",
    x"205F3629",
    x"205EDF09",
    x"205E880B",
    x"205E312E",
    x"205DDA74",
    x"205D83DC",
    x"205D2D65",
    x"205CD710",
    x"205C80DD",
    x"205C2ACC",
    x"205BD4DC",
    x"205B7F0D",
    x"205B2960",
    x"205AD3D5",
    x"205A7E6B",
    x"205A2922",
    x"2059D3FB",
    x"20597EF4",
    x"20592A0F",
    x"2058D54C",
    x"205880A9",
    x"20582C27",
    x"2057D7C6",
    x"20578386",
    x"20572F68",
    x"2056DB69",
    x"2056878C",
    x"205633CF",
    x"2055E034",
    x"20558CB8",
    x"2055395E",
    x"2054E623",
    x"2054930A",
    x"20544011",
    x"2053ED38",
    x"20539A7F",
    x"205347E7",
    x"2052F56F",
    x"2052A317",
    x"205250E0",
    x"2051FEC8",
    x"2051ACD1",
    x"20515AF9",
    x"20510941",
    x"2050B7AA",
    x"20506632",
    x"205014DA",
    x"204FC3A2",
    x"204F7289",
    x"204F2190",
    x"204ED0B7",
    x"204E7FFD",
    x"204E2F63",
    x"204DDEE8",
    x"204D8E8D",
    x"204D3E51",
    x"204CEE34",
    x"204C9E37",
    x"204C4E58",
    x"204BFE99",
    x"204BAEF9",
    x"204B5F79",
    x"204B1017",
    x"204AC0D4",
    x"204A71B0",
    x"204A22AB",
    x"2049D3C5",
    x"204984FE",
    x"20493655",
    x"2048E7CB",
    x"20489960",
    x"20484B13",
    x"2047FCE5",
    x"2047AED6",
    x"204760E5",
    x"20471312",
    x"2046C55E",
    x"204677C8",
    x"20462A50",
    x"2045DCF7",
    x"20458FBC",
    x"2045429F",
    x"2044F5A0",
    x"2044A8BF",
    x"20445BFC",
    x"20440F57",
    x"2043C2D0",
    x"20437667",
    x"20432A1B",
    x"2042DDEE",
    x"204291DE",
    x"204245EC",
    x"2041FA17",
    x"2041AE60",
    x"204162C7",
    x"2041174B",
    x"2040CBED",
    x"204080AC",
    x"20403588",
    x"203FEA82",
    x"203F9F99",
    x"203F54CD",
    x"203F0A1F",
    x"203EBF8D",
    x"203E7519",
    x"203E2AC2",
    x"203DE088",
    x"203D966A",
    x"203D4C6A",
    x"203D0287",
    x"203CB8C0",
    x"203C6F16",
    x"203C2589",
    x"203BDC19",
    x"203B92C5",
    x"203B498E",
    x"203B0074",
    x"203AB776",
    x"203A6E94",
    x"203A25D0",
    x"2039DD27",
    x"2039949B",
    x"20394C2B",
    x"203903D7",
    x"2038BBA0",
    x"20387385",
    x"20382B86",
    x"2037E3A3",
    x"20379BDC",
    x"20375431",
    x"20370CA2",
    x"2036C52F",
    x"20367DD8",
    x"2036369D",
    x"2035EF7D",
    x"2035A879",
    x"20356192",
    x"20351AC5",
    x"2034D415",
    x"20348D80",
    x"20344706",
    x"203400A8",
    x"2033BA66",
    x"2033743E",
    x"20332E33",
    x"2032E842",
    x"2032A26D",
    x"20325CB3",
    x"20321715",
    x"2031D191",
    x"20318C29",
    x"203146DC",
    x"203101AA",
    x"2030BC93",
    x"20307796",
    x"203032B5",
    x"202FEDEF",
    x"202FA943",
    x"202F64B2",
    x"202F203C",
    x"202EDBE1",
    x"202E97A1",
    x"202E537B",
    x"202E0F6F",
    x"202DCB7F",
    x"202D87A8",
    x"202D43ED",
    x"202D004B",
    x"202CBCC4",
    x"202C7958",
    x"202C3606",
    x"202BF2CE",
    x"202BAFB0",
    x"202B6CAC",
    x"202B29C3",
    x"202AE6F4",
    x"202AA43F",
    x"202A61A3",
    x"202A1F22",
    x"2029DCBB",
    x"20299A6E",
    x"2029583A",
    x"20291621",
    x"2028D421",
    x"2028923B",
    x"2028506F",
    x"20280EBC",
    x"2027CD23",
    x"20278BA4",
    x"20274A3E",
    x"202708F2",
    x"2026C7BF",
    x"202686A6",
    x"202645A6",
    x"202604C0",
    x"2025C3F2",
    x"2025833E",
    x"202542A4",
    x"20250222",
    x"2024C1BA",
    x"2024816B",
    x"20244135",
    x"20240118",
    x"2023C114",
    x"20238129",
    x"20234157",
    x"2023019E",
    x"2022C1FE",
    x"20228277",
    x"20224308",
    x"202203B2",
    x"2021C475",
    x"20218551",
    x"20214645",
    x"20210752",
    x"2020C877",
    x"202089B5",
    x"20204B0C",
    x"20200C7B",
    x"201FCE02",
    x"201F8FA2",
    x"201F515A",
    x"201F132A",
    x"201ED513",
    x"201E9714",
    x"201E592D",
    x"201E1B5E",
    x"201DDDA7",
    x"201DA009",
    x"201D6282",
    x"201D2514",
    x"201CE7BD",
    x"201CAA7F",
    x"201C6D58",
    x"201C3049",
    x"201BF352",
    x"201BB673",
    x"201B79AC",
    x"201B3CFC",
    x"201B0064",
    x"201AC3E4",
    x"201A877B",
    x"201A4B2A",
    x"201A0EF0",
    x"2019D2CE",
    x"201996C4",
    x"20195AD0",
    x"20191EF5",
    x"2018E330",
    x"2018A783",
    x"20186BED",
    x"2018306F",
    x"2017F507",
    x"2017B9B7",
    x"20177E7E",
    x"2017435C",
    x"20170852",
    x"2016CD5E",
    x"20169281",
    x"201657BB",
    x"20161D0D",
    x"2015E275",
    x"2015A7F4",
    x"20156D8A",
    x"20153336",
    x"2014F8FA",
    x"2014BED4",
    x"201484C4",
    x"20144ACC",
    x"201410EA",
    x"2013D71F",
    x"20139D6A",
    x"201363CC",
    x"20132A44",
    x"2012F0D3",
    x"2012B778",
    x"20127E33",
    x"20124505",
    x"20120BED",
    x"2011D2EC",
    x"20119A01",
    x"2011612C",
    x"2011286D",
    x"2010EFC4",
    x"2010B731",
    x"20107EB5",
    x"2010464E",
    x"20100DFE",
    x"200FD5C3",
    x"200F9D9F",
    x"200F6590",
    x"200F2D97",
    x"200EF5B5",
    x"200EBDE8",
    x"200E8630",
    x"200E4E8F",
    x"200E1703",
    x"200DDF8D",
    x"200DA82C",
    x"200D70E1",
    x"200D39AC",
    x"200D028C",
    x"200CCB82",
    x"200C948D",
    x"200C5DAE",
    x"200C26E4",
    x"200BF030",
    x"200BB990",
    x"200B8307",
    x"200B4C92",
    x"200B1633",
    x"200ADFE9",
    x"200AA9B4",
    x"200A7394",
    x"200A3D89",
    x"200A0794",
    x"2009D1B4",
    x"20099BE8",
    x"20096632",
    x"20093090",
    x"2008FB04",
    x"2008C58C",
    x"20089029",
    x"20085ADC",
    x"200825A2",
    x"2007F07E",
    x"2007BB6F",
    x"20078674",
    x"2007518D",
    x"20071CBC",
    x"2006E7FF",
    x"2006B357",
    x"20067EC3",
    x"20064A44",
    x"200615D9",
    x"2005E183",
    x"2005AD41",
    x"20057913",
    x"200544FA",
    x"200510F5",
    x"2004DD05",
    x"2004A929",
    x"20047561",
    x"200441AD",
    x"20040E0D",
    x"2003DA82",
    x"2003A70B",
    x"200373A7",
    x"20034058",
    x"20030D1D",
    x"2002D9F6",
    x"2002A6E3",
    x"200273E4",
    x"200240F8",
    x"20020E21",
    x"2001DB5D",
    x"2001A8AD",
    x"20017611",
    x"20014389",
    x"20011115",
    x"2000DEB4",
    x"2000AC67",
    x"20007A2D",
    x"20004807",
    x"200015F5",
    x"1FFFC7EC",
    x"1FFF6416",
    x"1FFF0066",
    x"1FFE9CDD",
    x"1FFE397B",
    x"1FFDD640",
    x"1FFD732C",
    x"1FFD103E",
    x"1FFCAD77",
    x"1FFC4AD7",
    x"1FFBE85D",
    x"1FFB8609",
    x"1FFB23DC",
    x"1FFAC1D5",
    x"1FFA5FF5",
    x"1FF9FE3A",
    x"1FF99CA6",
    x"1FF93B38",
    x"1FF8D9F0",
    x"1FF878CD",
    x"1FF817D1",
    x"1FF7B6FB",
    x"1FF7564A",
    x"1FF6F5BF",
    x"1FF6955A",
    x"1FF6351B",
    x"1FF5D501",
    x"1FF5750C",
    x"1FF5153D",
    x"1FF4B594",
    x"1FF4560F",
    x"1FF3F6B0",
    x"1FF39777",
    x"1FF33862",
    x"1FF2D973",
    x"1FF27AA8",
    x"1FF21C03",
    x"1FF1BD82",
    x"1FF15F27",
    x"1FF100F0",
    x"1FF0A2DE",
    x"1FF044F1",
    x"1FEFE728",
    x"1FEF8984",
    x"1FEF2C05",
    x"1FEECEAA",
    x"1FEE7173",
    x"1FEE1461",
    x"1FEDB773",
    x"1FED5AAA",
    x"1FECFE04",
    x"1FECA183",
    x"1FEC4526",
    x"1FEBE8ED",
    x"1FEB8CD8",
    x"1FEB30E7",
    x"1FEAD51A",
    x"1FEA7971",
    x"1FEA1DEB",
    x"1FE9C289",
    x"1FE9674B",
    x"1FE90C30",
    x"1FE8B13A",
    x"1FE85666",
    x"1FE7FBB6",
    x"1FE7A129",
    x"1FE746C0",
    x"1FE6EC7A",
    x"1FE69257",
    x"1FE63858",
    x"1FE5DE7B",
    x"1FE584C2",
    x"1FE52B2C",
    x"1FE4D1B8",
    x"1FE47868",
    x"1FE41F3A",
    x"1FE3C62F",
    x"1FE36D47",
    x"1FE31482",
    x"1FE2BBDF",
    x"1FE2635F",
    x"1FE20B02",
    x"1FE1B2C6",
    x"1FE15AAE",
    x"1FE102B8",
    x"1FE0AAE4",
    x"1FE05332",
    x"1FDFFBA3",
    x"1FDFA435",
    x"1FDF4CEA",
    x"1FDEF5C1",
    x"1FDE9EBA",
    x"1FDE47D5",
    x"1FDDF112",
    x"1FDD9A71",
    x"1FDD43F2",
    x"1FDCED94",
    x"1FDC9758",
    x"1FDC413E",
    x"1FDBEB45",
    x"1FDB956E",
    x"1FDB3FB8",
    x"1FDAEA24",
    x"1FDA94B1",
    x"1FDA3F60",
    x"1FD9EA30",
    x"1FD99521",
    x"1FD94033",
    x"1FD8EB67",
    x"1FD896BB",
    x"1FD84231",
    x"1FD7EDC8",
    x"1FD7997F",
    x"1FD74558",
    x"1FD6F151",
    x"1FD69D6B",
    x"1FD649A6",
    x"1FD5F601",
    x"1FD5A27E",
    x"1FD54F1B",
    x"1FD4FBD8",
    x"1FD4A8B6",
    x"1FD455B4",
    x"1FD402D3",
    x"1FD3B012",
    x"1FD35D71",
    x"1FD30AF1",
    x"1FD2B891",
    x"1FD26651",
    x"1FD21431",
    x"1FD1C231",
    x"1FD17051",
    x"1FD11E91",
    x"1FD0CCF1",
    x"1FD07B71",
    x"1FD02A11",
    x"1FCFD8D0",
    x"1FCF87AF",
    x"1FCF36AE",
    x"1FCEE5CC",
    x"1FCE950B",
    x"1FCE4468",
    x"1FCDF3E5",
    x"1FCDA381",
    x"1FCD533D",
    x"1FCD0318",
    x"1FCCB313",
    x"1FCC632D",
    x"1FCC1365",
    x"1FCBC3BD",
    x"1FCB7434",
    x"1FCB24CB",
    x"1FCAD580",
    x"1FCA8654",
    x"1FCA3747",
    x"1FC9E859",
    x"1FC99989",
    x"1FC94AD9",
    x"1FC8FC47",
    x"1FC8ADD3",
    x"1FC85F7F",
    x"1FC81149",
    x"1FC7C331",
    x"1FC77538",
    x"1FC7275E",
    x"1FC6D9A2",
    x"1FC68C04",
    x"1FC63E84",
    x"1FC5F123",
    x"1FC5A3E0",
    x"1FC556BB",
    x"1FC509B4",
    x"1FC4BCCB",
    x"1FC47000",
    x"1FC42354",
    x"1FC3D6C5",
    x"1FC38A54",
    x"1FC33E01",
    x"1FC2F1CB",
    x"1FC2A5B4",
    x"1FC259BA",
    x"1FC20DDE",
    x"1FC1C21F",
    x"1FC1767E",
    x"1FC12AFB",
    x"1FC0DF94",
    x"1FC0944C",
    x"1FC04921",
    x"1FBFFE13",
    x"1FBFB322",
    x"1FBF684F",
    x"1FBF1D99",
    x"1FBED300",
    x"1FBE8884",
    x"1FBE3E25",
    x"1FBDF3E3",
    x"1FBDA9BE",
    x"1FBD5FB7",
    x"1FBD15CC",
    x"1FBCCBFD",
    x"1FBC824C",
    x"1FBC38B8",
    x"1FBBEF40",
    x"1FBBA5E5",
    x"1FBB5CA6",
    x"1FBB1384",
    x"1FBACA7F",
    x"1FBA8196",
    x"1FBA38CA",
    x"1FB9F01A",
    x"1FB9A786",
    x"1FB95F0F",
    x"1FB916B4",
    x"1FB8CE75",
    x"1FB88653",
    x"1FB83E4C",
    x"1FB7F662",
    x"1FB7AE94",
    x"1FB766E1",
    x"1FB71F4B",
    x"1FB6D7D1",
    x"1FB69073",
    x"1FB64930",
    x"1FB60209",
    x"1FB5BAFF",
    x"1FB5740F",
    x"1FB52D3C",
    x"1FB4E684",
    x"1FB49FE8",
    x"1FB45967",
    x"1FB41302",
    x"1FB3CCB8",
    x"1FB3868A",
    x"1FB34077",
    x"1FB2FA80",
    x"1FB2B4A3",
    x"1FB26EE2",
    x"1FB2293D",
    x"1FB1E3B2",
    x"1FB19E43",
    x"1FB158EF",
    x"1FB113B5",
    x"1FB0CE97",
    x"1FB08994",
    x"1FB044AC",
    x"1FAFFFDE",
    x"1FAFBB2C",
    x"1FAF7694",
    x"1FAF3217",
    x"1FAEEDB5",
    x"1FAEA96D",
    x"1FAE6540",
    x"1FAE212E",
    x"1FADDD37",
    x"1FAD9959",
    x"1FAD5597",
    x"1FAD11EF",
    x"1FACCE61",
    x"1FAC8AED",
    x"1FAC4794",
    x"1FAC0455",
    x"1FABC131",
    x"1FAB7E26",
    x"1FAB3B36",
    x"1FAAF860",
    x"1FAAB5A4",
    x"1FAA7302",
    x"1FAA307A",
    x"1FA9EE0C",
    x"1FA9ABB8",
    x"1FA9697E",
    x"1FA9275E",
    x"1FA8E557",
    x"1FA8A36B",
    x"1FA86198",
    x"1FA81FDE",
    x"1FA7DE3F",
    x"1FA79CB9",
    x"1FA75B4C",
    x"1FA719F9",
    x"1FA6D8C0",
    x"1FA697A0",
    x"1FA6569A",
    x"1FA615AC",
    x"1FA5D4D9",
    x"1FA5941E",
    x"1FA5537D",
    x"1FA512F5",
    x"1FA4D286",
    x"1FA49230",
    x"1FA451F4",
    x"1FA411D0",
    x"1FA3D1C6",
    x"1FA391D4",
    x"1FA351FC",
    x"1FA3123C",
    x"1FA2D296",
    x"1FA29308",
    x"1FA25393",
    x"1FA21437",
    x"1FA1D4F3",
    x"1FA195C8",
    x"1FA156B6",
    x"1FA117BC",
    x"1FA0D8DB",
    x"1FA09A13",
    x"1FA05B63",
    x"1FA01CCC",
    x"1F9FDE4D",
    x"1F9F9FE6",
    x"1F9F6198",
    x"1F9F2362",
    x"1F9EE544",
    x"1F9EA73F",
    x"1F9E6951",
    x"1F9E2B7C",
    x"1F9DEDBF",
    x"1F9DB01A",
    x"1F9D728E",
    x"1F9D3519",
    x"1F9CF7BC",
    x"1F9CBA77",
    x"1F9C7D4B",
    x"1F9C4036",
    x"1F9C0338",
    x"1F9BC653",
    x"1F9B8985",
    x"1F9B4CD0",
    x"1F9B1031",
    x"1F9AD3AB",
    x"1F9A973C",
    x"1F9A5AE5",
    x"1F9A1EA5",
    x"1F99E27D",
    x"1F99A66C",
    x"1F996A73",
    x"1F992E91",
    x"1F98F2C6",
    x"1F98B713",
    x"1F987B77",
    x"1F983FF3",
    x"1F980485",
    x"1F97C92F",
    x"1F978DF0",
    x"1F9752C8",
    x"1F9717B7",
    x"1F96DCBE",
    x"1F96A1DB",
    x"1F96670F",
    x"1F962C5A",
    x"1F95F1BD",
    x"1F95B736",
    x"1F957CC5",
    x"1F95426C",
    x"1F95082A",
    x"1F94CDFE",
    x"1F9493E9",
    x"1F9459EA",
    x"1F942002",
    x"1F93E631",
    x"1F93AC76",
    x"1F9372D2",
    x"1F933945",
    x"1F92FFCE",
    x"1F92C66D",
    x"1F928D23",
    x"1F9253EF",
    x"1F921AD1",
    x"1F91E1CA",
    x"1F91A8D9",
    x"1F916FFE",
    x"1F913739",
    x"1F90FE8B",
    x"1F90C5F2",
    x"1F908D70",
    x"1F905504",
    x"1F901CAE",
    x"1F8FE46D",
    x"1F8FAC43",
    x"1F8F742F",
    x"1F8F3C30",
    x"1F8F0448",
    x"1F8ECC75",
    x"1F8E94B8",
    x"1F8E5D11",
    x"1F8E257F",
    x"1F8DEE03",
    x"1F8DB69D",
    x"1F8D7F4D",
    x"1F8D4812",
    x"1F8D10EC",
    x"1F8CD9DD",
    x"1F8CA2E2",
    x"1F8C6BFD",
    x"1F8C352E",
    x"1F8BFE74",
    x"1F8BC7CF",
    x"1F8B9140",
    x"1F8B5AC6",
    x"1F8B2461",
    x"1F8AEE11",
    x"1F8AB7D7",
    x"1F8A81B1",
    x"1F8A4BA1",
    x"1F8A15A6",
    x"1F89DFC0",
    x"1F89A9F0",
    x"1F897434",
    x"1F893E8D",
    x"1F8908FB",
    x"1F88D37E",
    x"1F889E16",
    x"1F8868C2",
    x"1F883384",
    x"1F87FE5A",
    x"1F87C945",
    x"1F879445",
    x"1F875F59",
    x"1F872A82",
    x"1F86F5C0",
    x"1F86C112",
    x"1F868C79",
    x"1F8657F4",
    x"1F862384",
    x"1F85EF29",
    x"1F85BAE1",
    x"1F8586AF",
    x"1F855290",
    x"1F851E86",
    x"1F84EA90",
    x"1F84B6AF",
    x"1F8482E2",
    x"1F844F29",
    x"1F841B84",
    x"1F83E7F3",
    x"1F83B477",
    x"1F83810E",
    x"1F834DBA",
    x"1F831A79",
    x"1F82E74D",
    x"1F82B435",
    x"1F828130",
    x"1F824E40",
    x"1F821B63",
    x"1F81E89A",
    x"1F81B5E5",
    x"1F818344",
    x"1F8150B7",
    x"1F811E3D",
    x"1F80EBD7",
    x"1F80B985",
    x"1F808746",
    x"1F80551B",
    x"1F802304",
    x"1F7FE200",
    x"1F7F7E1F",
    x"1F7F1A65",
    x"1F7EB6D2",
    x"1F7E5366",
    x"1F7DF021",
    x"1F7D8D03",
    x"1F7D2A0B",
    x"1F7CC73A",
    x"1F7C648F",
    x"1F7C020B",
    x"1F7B9FAE",
    x"1F7B3D76",
    x"1F7ADB66",
    x"1F7A797B",
    x"1F7A17B7",
    x"1F79B619",
    x"1F7954A0",
    x"1F78F34E",
    x"1F789222",
    x"1F78311C",
    x"1F77D03C",
    x"1F776F81",
    x"1F770EED",
    x"1F76AE7E",
    x"1F764E34",
    x"1F75EE11",
    x"1F758E12",
    x"1F752E3A",
    x"1F74CE86",
    x"1F746EF8",
    x"1F740F90",
    x"1F73B04C",
    x"1F73512E",
    x"1F72F235",
    x"1F729361",
    x"1F7234B2",
    x"1F71D627",
    x"1F7177C2",
    x"1F711982",
    x"1F70BB66",
    x"1F705D6F",
    x"1F6FFF9D",
    x"1F6FA1F0",
    x"1F6F4467",
    x"1F6EE702",
    x"1F6E89C2",
    x"1F6E2CA7",
    x"1F6DCFAF",
    x"1F6D72DC",
    x"1F6D162E",
    x"1F6CB9A3",
    x"1F6C5D3D",
    x"1F6C00FA",
    x"1F6BA4DC",
    x"1F6B48E1",
    x"1F6AED0B",
    x"1F6A9158",
    x"1F6A35C9",
    x"1F69DA5E",
    x"1F697F17",
    x"1F6923F3",
    x"1F68C8F2",
    x"1F686E16",
    x"1F68135C",
    x"1F67B8C7",
    x"1F675E54",
    x"1F670405",
    x"1F66A9D9",
    x"1F664FD0",
    x"1F65F5EB",
    x"1F659C28",
    x"1F654289",
    x"1F64E90C",
    x"1F648FB2",
    x"1F64367C",
    x"1F63DD68",
    x"1F638477",
    x"1F632BA8",
    x"1F62D2FD",
    x"1F627A74",
    x"1F62220D",
    x"1F61C9C9",
    x"1F6171A7",
    x"1F6119A8",
    x"1F60C1CB",
    x"1F606A11",
    x"1F601278",
    x"1F5FBB02",
    x"1F5F63AE",
    x"1F5F0C7C",
    x"1F5EB56C",
    x"1F5E5E7F",
    x"1F5E07B3",
    x"1F5DB109",
    x"1F5D5A80",
    x"1F5D041A",
    x"1F5CADD5",
    x"1F5C57B2",
    x"1F5C01B1",
    x"1F5BABD1",
    x"1F5B5612",
    x"1F5B0075",
    x"1F5AAAFA",
    x"1F5A55A0",
    x"1F5A0067",
    x"1F59AB4F",
    x"1F595659",
    x"1F590184",
    x"1F58ACD0",
    x"1F58583D",
    x"1F5803CB",
    x"1F57AF7A",
    x"1F575B4A",
    x"1F57073B",
    x"1F56B34C",
    x"1F565F7F",
    x"1F560BD2",
    x"1F55B845",
    x"1F5564DA",
    x"1F55118F",
    x"1F54BE64",
    x"1F546B5A",
    x"1F541870",
    x"1F53C5A7",
    x"1F5372FE",
    x"1F532075",
    x"1F52CE0C",
    x"1F527BC4",
    x"1F52299C",
    x"1F51D793",
    x"1F5185AB",
    x"1F5133E3",
    x"1F50E23B",
    x"1F5090B2",
    x"1F503F49",
    x"1F4FEE01",
    x"1F4F9CD8",
    x"1F4F4BCE",
    x"1F4EFAE4",
    x"1F4EAA1A",
    x"1F4E596F",
    x"1F4E08E4",
    x"1F4DB878",
    x"1F4D682C",
    x"1F4D17FF",
    x"1F4CC7F1",
    x"1F4C7803",
    x"1F4C2833",
    x"1F4BD883",
    x"1F4B88F2",
    x"1F4B3980",
    x"1F4AEA2D",
    x"1F4A9AF9",
    x"1F4A4BE4",
    x"1F49FCEE",
    x"1F49AE17",
    x"1F495F5E",
    x"1F4910C4",
    x"1F48C249",
    x"1F4873EC",
    x"1F4825AE",
    x"1F47D78F",
    x"1F47898E",
    x"1F473BAB",
    x"1F46EDE7",
    x"1F46A042",
    x"1F4652BA",
    x"1F460551",
    x"1F45B806",
    x"1F456AD9",
    x"1F451DCA",
    x"1F44D0DA",
    x"1F448407",
    x"1F443753",
    x"1F43EABC",
    x"1F439E43",
    x"1F4351E8",
    x"1F4305AB",
    x"1F42B98C",
    x"1F426D8A",
    x"1F4221A6",
    x"1F41D5E0",
    x"1F418A37",
    x"1F413EAC",
    x"1F40F33E",
    x"1F40A7EE",
    x"1F405CBB",
    x"1F4011A5",
    x"1F3FC6AD",
    x"1F3F7BD2",
    x"1F3F3114",
    x"1F3EE674",
    x"1F3E9BF0",
    x"1F3E518A",
    x"1F3E0741",
    x"1F3DBD14",
    x"1F3D7305",
    x"1F3D2912",
    x"1F3CDF3D",
    x"1F3C9584",
    x"1F3C4BE8",
    x"1F3C0269",
    x"1F3BB906",
    x"1F3B6FC0",
    x"1F3B2697",
    x"1F3ADD8A",
    x"1F3A949A",
    x"1F3A4BC6",
    x"1F3A030F",
    x"1F39BA74",
    x"1F3971F5",
    x"1F392992",
    x"1F38E14C",
    x"1F389922",
    x"1F385115",
    x"1F380923",
    x"1F37C14E",
    x"1F377994",
    x"1F3731F7",
    x"1F36EA75",
    x"1F36A30F",
    x"1F365BC6",
    x"1F361498",
    x"1F35CD86",
    x"1F35868F",
    x"1F353FB4",
    x"1F34F8F5",
    x"1F34B252",
    x"1F346BCA",
    x"1F34255E",
    x"1F33DF0D",
    x"1F3398D7",
    x"1F3352BD",
    x"1F330CBF",
    x"1F32C6DB",
    x"1F328113",
    x"1F323B67",
    x"1F31F5D5",
    x"1F31B05E",
    x"1F316B03",
    x"1F3125C3",
    x"1F30E09E",
    x"1F309B93",
    x"1F3056A4",
    x"1F3011D0",
    x"1F2FCD16",
    x"1F2F8877",
    x"1F2F43F3",
    x"1F2EFF8A",
    x"1F2EBB3C",
    x"1F2E7708",
    x"1F2E32EF",
    x"1F2DEEF0",
    x"1F2DAB0C",
    x"1F2D6743",
    x"1F2D2393",
    x"1F2CDFFF",
    x"1F2C9C84",
    x"1F2C5924",
    x"1F2C15DF",
    x"1F2BD2B3",
    x"1F2B8FA2",
    x"1F2B4CAB",
    x"1F2B09CE",
    x"1F2AC70B",
    x"1F2A8463",
    x"1F2A41D4",
    x"1F29FF5F",
    x"1F29BD04",
    x"1F297AC4",
    x"1F29389D",
    x"1F28F68F",
    x"1F28B49C",
    x"1F2872C2",
    x"1F283102",
    x"1F27EF5C",
    x"1F27ADCF",
    x"1F276C5C",
    x"1F272B03",
    x"1F26E9C3",
    x"1F26A89C",
    x"1F26678F",
    x"1F26269B",
    x"1F25E5C1",
    x"1F25A500",
    x"1F256458",
    x"1F2523C9",
    x"1F24E354",
    x"1F24A2F8",
    x"1F2462B4",
    x"1F24228A",
    x"1F23E279",
    x"1F23A281",
    x"1F2362A2",
    x"1F2322DC",
    x"1F22E32F",
    x"1F22A39B",
    x"1F22641F",
    x"1F2224BD",
    x"1F21E573",
    x"1F21A641",
    x"1F216729",
    x"1F212829",
    x"1F20E941",
    x"1F20AA73",
    x"1F206BBC",
    x"1F202D1E",
    x"1F1FEE99",
    x"1F1FB02C",
    x"1F1F71D7",
    x"1F1F339B",
    x"1F1EF577",
    x"1F1EB76B",
    x"1F1E7978",
    x"1F1E3B9C",
    x"1F1DFDD9",
    x"1F1DC02E",
    x"1F1D829B",
    x"1F1D4520",
    x"1F1D07BD",
    x"1F1CCA72",
    x"1F1C8D3F",
    x"1F1C5023",
    x"1F1C1320",
    x"1F1BD635",
    x"1F1B9961",
    x"1F1B5CA5",
    x"1F1B2000",
    x"1F1AE374",
    x"1F1AA6FF",
    x"1F1A6AA1",
    x"1F1A2E5B",
    x"1F19F22D",
    x"1F19B616",
    x"1F197A17",
    x"1F193E2F",
    x"1F19025E",
    x"1F18C6A5",
    x"1F188B03",
    x"1F184F78",
    x"1F181405",
    x"1F17D8A9",
    x"1F179D64",
    x"1F176236",
    x"1F17271F",
    x"1F16EC1F",
    x"1F16B136",
    x"1F167665",
    x"1F163BAA",
    x"1F160106",
    x"1F15C679",
    x"1F158C03",
    x"1F1551A4",
    x"1F15175B",
    x"1F14DD29",
    x"1F14A30E",
    x"1F14690A",
    x"1F142F1C",
    x"1F13F545",
    x"1F13BB85",
    x"1F1381DB",
    x"1F134847",
    x"1F130ECA",
    x"1F12D564",
    x"1F129C13",
    x"1F1262DA",
    x"1F1229B6",
    x"1F11F0A9",
    x"1F11B7B2",
    x"1F117ED2",
    x"1F114607",
    x"1F110D53",
    x"1F10D4B5",
    x"1F109C2D",
    x"1F1063BB",
    x"1F102B5F",
    x"1F0FF319",
    x"1F0FBAE9",
    x"1F0F82CF",
    x"1F0F4ACB",
    x"1F0F12DC",
    x"1F0EDB04",
    x"1F0EA341",
    x"1F0E6B94",
    x"1F0E33FD",
    x"1F0DFC7C",
    x"1F0DC510",
    x"1F0D8DBA",
    x"1F0D5679",
    x"1F0D1F4E",
    x"1F0CE839",
    x"1F0CB139",
    x"1F0C7A4E",
    x"1F0C4379",
    x"1F0C0CB9",
    x"1F0BD60F",
    x"1F0B9F7A",
    x"1F0B68FB",
    x"1F0B3290",
    x"1F0AFC3B",
    x"1F0AC5FB",
    x"1F0A8FD0",
    x"1F0A59BB",
    x"1F0A23BA",
    x"1F09EDCF",
    x"1F09B7F8",
    x"1F098237",
    x"1F094C8B",
    x"1F0916F3",
    x"1F08E171",
    x"1F08AC03",
    x"1F0876AA",
    x"1F084166",
    x"1F080C37",
    x"1F07D71D",
    x"1F07A217",
    x"1F076D26",
    x"1F07384A",
    x"1F070382",
    x"1F06CECF",
    x"1F069A31",
    x"1F0665A7",
    x"1F063131",
    x"1F05FCD0",
    x"1F05C884",
    x"1F05944C",
    x"1F056028",
    x"1F052C18",
    x"1F04F81D",
    x"1F04C437",
    x"1F049064",
    x"1F045CA6",
    x"1F0428FC",
    x"1F03F566",
    x"1F03C1E4",
    x"1F038E76",
    x"1F035B1D",
    x"1F0327D7",
    x"1F02F4A6",
    x"1F02C188",
    x"1F028E7E",
    x"1F025B89",
    x"1F0228A7",
    x"1F01F5D9",
    x"1F01C31F",
    x"1F019078",
    x"1F015DE6",
    x"1F012B67",
    x"1F00F8FC",
    x"1F00C6A4",
    x"1F009461",
    x"1F006231",
    x"1F003014",
    x"1EFFFC16",
    x"1EFF982B",
    x"1EFF3467",
    x"1EFED0CA",
    x"1EFE6D54",
    x"1EFE0A05",
    x"1EFDA6DC",
    x"1EFD43DA",
    x"1EFCE0FF",
    x"1EFC7E4A",
    x"1EFC1BBC",
    x"1EFBB955",
    x"1EFB5714",
    x"1EFAF4F9",
    x"1EFA9304",
    x"1EFA3136",
    x"1EF9CF8E",
    x"1EF96E0C",
    x"1EF90CB0",
    x"1EF8AB7A",
    x"1EF84A6A",
    x"1EF7E980",
    x"1EF788BB",
    x"1EF7281D",
    x"1EF6C7A4",
    x"1EF66751",
    x"1EF60723",
    x"1EF5A71B",
    x"1EF54739",
    x"1EF4E77B",
    x"1EF487E4",
    x"1EF42871",
    x"1EF3C924",
    x"1EF369FC",
    x"1EF30AF9",
    x"1EF2AC1C",
    x"1EF24D63",
    x"1EF1EECF",
    x"1EF19060",
    x"1EF13216",
    x"1EF0D3F1",
    x"1EF075F1",
    x"1EF01815",
    x"1EEFBA5E",
    x"1EEF5CCB",
    x"1EEEFF5D",
    x"1EEEA214",
    x"1EEE44EF",
    x"1EEDE7EE",
    x"1EED8B11",
    x"1EED2E59",
    x"1EECD1C5",
    x"1EEC7555",
    x"1EEC190A",
    x"1EEBBCE2",
    x"1EEB60DE",
    x"1EEB04FE",
    x"1EEAA942",
    x"1EEA4DAA",
    x"1EE9F235",
    x"1EE996E5",
    x"1EE93BB7",
    x"1EE8E0AE",
    x"1EE885C8",
    x"1EE82B05",
    x"1EE7D066",
    x"1EE775EB",
    x"1EE71B92",
    x"1EE6C15D",
    x"1EE6674B",
    x"1EE60D5C",
    x"1EE5B391",
    x"1EE559E8",
    x"1EE50062",
    x"1EE4A700",
    x"1EE44DC0",
    x"1EE3F4A3",
    x"1EE39BA9",
    x"1EE342D1",
    x"1EE2EA1C",
    x"1EE2918A",
    x"1EE2391B",
    x"1EE1E0CE",
    x"1EE188A3",
    x"1EE1309B",
    x"1EE0D8B5",
    x"1EE080F2",
    x"1EE02950",
    x"1EDFD1D1",
    x"1EDF7A74",
    x"1EDF233A",
    x"1EDECC21",
    x"1EDE752A",
    x"1EDE1E55",
    x"1EDDC7A2",
    x"1EDD7111",
    x"1EDD1AA2",
    x"1EDCC455",
    x"1EDC6E29",
    x"1EDC181E",
    x"1EDBC236",
    x"1EDB6C6F",
    x"1EDB16C9",
    x"1EDAC145",
    x"1EDA6BE2",
    x"1EDA16A1",
    x"1ED9C180",
    x"1ED96C81",
    x"1ED917A4",
    x"1ED8C2E7",
    x"1ED86E4B",
    x"1ED819D1",
    x"1ED7C577",
    x"1ED7713E",
    x"1ED71D27",
    x"1ED6C930",
    x"1ED67559",
    x"1ED621A4",
    x"1ED5CE0F",
    x"1ED57A9B",
    x"1ED52747",
    x"1ED4D414",
    x"1ED48102",
    x"1ED42E0F",
    x"1ED3DB3E",
    x"1ED3888C",
    x"1ED335FB",
    x"1ED2E38A",
    x"1ED29139",
    x"1ED23F09",
    x"1ED1ECF8",
    x"1ED19B07",
    x"1ED14937",
    x"1ED0F786",
    x"1ED0A5F5",
    x"1ED05484",
    x"1ED00333",
    x"1ECFB202",
    x"1ECF60F0",
    x"1ECF0FFE",
    x"1ECEBF2C",
    x"1ECE6E79",
    x"1ECE1DE5",
    x"1ECDCD71",
    x"1ECD7D1D",
    x"1ECD2CE8",
    x"1ECCDCD2",
    x"1ECC8CDB",
    x"1ECC3D04",
    x"1ECBED4B",
    x"1ECB9DB2",
    x"1ECB4E38",
    x"1ECAFEDD",
    x"1ECAAFA1",
    x"1ECA6084",
    x"1ECA1186",
    x"1EC9C2A6",
    x"1EC973E6",
    x"1EC92544",
    x"1EC8D6C1",
    x"1EC8885C",
    x"1EC83A16",
    x"1EC7EBEF",
    x"1EC79DE6",
    x"1EC74FFB",
    x"1EC7022F",
    x"1EC6B481",
    x"1EC666F2",
    x"1EC61981",
    x"1EC5CC2E",
    x"1EC57EF9",
    x"1EC531E3",
    x"1EC4E4EA",
    x"1EC49810",
    x"1EC44B54",
    x"1EC3FEB5",
    x"1EC3B235",
    x"1EC365D2",
    x"1EC3198D",
    x"1EC2CD66",
    x"1EC2815D",
    x"1EC23571",
    x"1EC1E9A3",
    x"1EC19DF2",
    x"1EC1525F",
    x"1EC106EA",
    x"1EC0BB92",
    x"1EC07057",
    x"1EC0253A",
    x"1EBFDA3A",
    x"1EBF8F58",
    x"1EBF4492",
    x"1EBEF9EA",
    x"1EBEAF5F",
    x"1EBE64F1",
    x"1EBE1AA0",
    x"1EBDD06C",
    x"1EBD8655",
    x"1EBD3C5B",
    x"1EBCF27E",
    x"1EBCA8BE",
    x"1EBC5F1A",
    x"1EBC1594",
    x"1EBBCC29",
    x"1EBB82DC",
    x"1EBB39AB",
    x"1EBAF097",
    x"1EBAA79F",
    x"1EBA5EC4",
    x"1EBA1605",
    x"1EB9CD63",
    x"1EB984DD",
    x"1EB93C73",
    x"1EB8F426",
    x"1EB8ABF4",
    x"1EB863DF",
    x"1EB81BE6",
    x"1EB7D409",
    x"1EB78C49",
    x"1EB744A4",
    x"1EB6FD1B",
    x"1EB6B5AE",
    x"1EB66E5D",
    x"1EB62728",
    x"1EB5E00E",
    x"1EB59911",
    x"1EB5522F",
    x"1EB50B68",
    x"1EB4C4BE",
    x"1EB47E2F",
    x"1EB437BB",
    x"1EB3F163",
    x"1EB3AB27",
    x"1EB36505",
    x"1EB31F00",
    x"1EB2D915",
    x"1EB29346",
    x"1EB24D92",
    x"1EB207F9",
    x"1EB1C27C",
    x"1EB17D1A",
    x"1EB137D2",
    x"1EB0F2A6",
    x"1EB0AD95",
    x"1EB0689E",
    x"1EB023C3",
    x"1EAFDF02",
    x"1EAF9A5D",
    x"1EAF55D2",
    x"1EAF1162",
    x"1EAECD0C",
    x"1EAE88D1",
    x"1EAE44B1",
    x"1EAE00AC",
    x"1EADBCC1",
    x"1EAD78F0",
    x"1EAD353A",
    x"1EACF19F",
    x"1EACAE1D",
    x"1EAC6AB7",
    x"1EAC276A",
    x"1EABE438",
    x"1EABA120",
    x"1EAB5E22",
    x"1EAB1B3E",
    x"1EAAD875",
    x"1EAA95C5",
    x"1EAA5330",
    x"1EAA10B4",
    x"1EA9CE52",
    x"1EA98C0B",
    x"1EA949DD",
    x"1EA907C9",
    x"1EA8C5CF",
    x"1EA883EF",
    x"1EA84228",
    x"1EA8007B",
    x"1EA7BEE7",
    x"1EA77D6E",
    x"1EA73C0D",
    x"1EA6FAC7",
    x"1EA6B99A",
    x"1EA67886",
    x"1EA6378B",
    x"1EA5F6AA",
    x"1EA5B5E3",
    x"1EA57534",
    x"1EA5349F",
    x"1EA4F423",
    x"1EA4B3C0",
    x"1EA47377",
    x"1EA43346",
    x"1EA3F32F",
    x"1EA3B330",
    x"1EA3734B",
    x"1EA3337E",
    x"1EA2F3CA",
    x"1EA2B430",
    x"1EA274AE",
    x"1EA23544",
    x"1EA1F5F4",
    x"1EA1B6BC",
    x"1EA1779D",
    x"1EA13897",
    x"1EA0F9A9",
    x"1EA0BAD4",
    x"1EA07C17",
    x"1EA03D73",
    x"1E9FFEE7",
    x"1E9FC074",
    x"1E9F8219",
    x"1E9F43D6",
    x"1E9F05AC",
    x"1E9EC799",
    x"1E9E89A0",
    x"1E9E4BBE",
    x"1E9E0DF4",
    x"1E9DD043",
    x"1E9D92AA",
    x"1E9D5528",
    x"1E9D17BF",
    x"1E9CDA6E",
    x"1E9C9D35",
    x"1E9C6013",
    x"1E9C2309",
    x"1E9BE618",
    x"1E9BA93E",
    x"1E9B6C7B",
    x"1E9B2FD1",
    x"1E9AF33E",
    x"1E9AB6C3",
    x"1E9A7A5F",
    x"1E9A3E13",
    x"1E9A01DF",
    x"1E99C5C2",
    x"1E9989BC",
    x"1E994DCE",
    x"1E9911F7",
    x"1E98D638",
    x"1E989A90",
    x"1E985EFF",
    x"1E982386",
    x"1E97E824",
    x"1E97ACD9",
    x"1E9771A5",
    x"1E973688",
    x"1E96FB82",
    x"1E96C093",
    x"1E9685BB",
    x"1E964AFB",
    x"1E961051",
    x"1E95D5BE",
    x"1E959B42",
    x"1E9560DD",
    x"1E95268E",
    x"1E94EC57",
    x"1E94B236",
    x"1E94782B",
    x"1E943E38",
    x"1E94045B",
    x"1E93CA94",
    x"1E9390E4",
    x"1E93574B",
    x"1E931DC8",
    x"1E92E45C",
    x"1E92AB06",
    x"1E9271C6",
    x"1E92389D",
    x"1E91FF8A",
    x"1E91C68D",
    x"1E918DA7",
    x"1E9154D7",
    x"1E911C1C",
    x"1E90E379",
    x"1E90AAEB",
    x"1E907273",
    x"1E903A11",
    x"1E9001C6",
    x"1E8FC990",
    x"1E8F9170",
    x"1E8F5966",
    x"1E8F2172",
    x"1E8EE994",
    x"1E8EB1CC",
    x"1E8E7A19",
    x"1E8E427C",
    x"1E8E0AF5",
    x"1E8DD384",
    x"1E8D9C28",
    x"1E8D64E2",
    x"1E8D2DB1",
    x"1E8CF696",
    x"1E8CBF91",
    x"1E8C88A0",
    x"1E8C51C6",
    x"1E8C1B01",
    x"1E8BE451",
    x"1E8BADB6",
    x"1E8B7731",
    x"1E8B40C1",
    x"1E8B0A66",
    x"1E8AD421",
    x"1E8A9DF1",
    x"1E8A67D6",
    x"1E8A31D0",
    x"1E89FBDF",
    x"1E89C603",
    x"1E89903C",
    x"1E895A8A",
    x"1E8924ED",
    x"1E88EF65",
    x"1E88B9F2",
    x"1E888494",
    x"1E884F4B",
    x"1E881A16",
    x"1E87E4F6",
    x"1E87AFEB",
    x"1E877AF5",
    x"1E874613",
    x"1E871146",
    x"1E86DC8D",
    x"1E86A7EA",
    x"1E86735A",
    x"1E863EDF",
    x"1E860A79",
    x"1E85D627",
    x"1E85A1EA",
    x"1E856DC1",
    x"1E8539AC",
    x"1E8505AC",
    x"1E84D1C0",
    x"1E849DE8",
    x"1E846A24",
    x"1E843675",
    x"1E8402DA",
    x"1E83CF53",
    x"1E839BE0",
    x"1E836881",
    x"1E833536",
    x"1E8301FF",
    x"1E82CEDD",
    x"1E829BCE",
    x"1E8268D3",
    x"1E8235EC",
    x"1E820319",
    x"1E81D059",
    x"1E819DAE",
    x"1E816B16",
    x"1E813892",
    x"1E810622",
    x"1E80D3C5",
    x"1E80A17C",
    x"1E806F47",
    x"1E803D26",
    x"1E800B17",
    x"1E7FB23A",
    x"1E7F4E6C",
    x"1E7EEAC4",
    x"1E7E8744",
    x"1E7E23EB",
    x"1E7DC0B8",
    x"1E7D5DAC",
    x"1E7CFAC7",
    x"1E7C9808",
    x"1E7C3570",
    x"1E7BD2FE",
    x"1E7B70B3",
    x"1E7B0E8E",
    x"1E7AAC90",
    x"1E7A4AB8",
    x"1E79E905",
    x"1E798779",
    x"1E792614",
    x"1E78C4D4",
    x"1E7863BA",
    x"1E7802C6",
    x"1E77A1F8",
    x"1E77414F",
    x"1E76E0CD",
    x"1E768070",
    x"1E762038",
    x"1E75C026",
    x"1E75603A",
    x"1E750073",
    x"1E74A0D2",
    x"1E744156",
    x"1E73E1FF",
    x"1E7382CD",
    x"1E7323C0",
    x"1E72C4D9",
    x"1E726617",
    x"1E720779",
    x"1E71A901",
    x"1E714AAD",
    x"1E70EC7E",
    x"1E708E74",
    x"1E70308F",
    x"1E6FD2CE",
    x"1E6F7532",
    x"1E6F17BB",
    x"1E6EBA68",
    x"1E6E5D39",
    x"1E6E002F",
    x"1E6DA349",
    x"1E6D4687",
    x"1E6CE9EA",
    x"1E6C8D71",
    x"1E6C311B",
    x"1E6BD4EA",
    x"1E6B78DD",
    x"1E6B1CF4",
    x"1E6AC12E",
    x"1E6A658D",
    x"1E6A0A0F",
    x"1E69AEB5",
    x"1E69537F",
    x"1E68F86C",
    x"1E689D7C",
    x"1E6842B1",
    x"1E67E808",
    x"1E678D83",
    x"1E673322",
    x"1E66D8E3",
    x"1E667EC8",
    x"1E6624D0",
    x"1E65CAFC",
    x"1E65714A",
    x"1E6517BB",
    x"1E64BE4F",
    x"1E646506",
    x"1E640BE0",
    x"1E63B2DD",
    x"1E6359FD",
    x"1E63013F",
    x"1E62A8A4",
    x"1E62502B",
    x"1E61F7D5",
    x"1E619FA1",
    x"1E614790",
    x"1E60EFA1",
    x"1E6097D5",
    x"1E60402B",
    x"1E5FE8A3",
    x"1E5F913D",
    x"1E5F39F9",
    x"1E5EE2D8",
    x"1E5E8BD8",
    x"1E5E34FA",
    x"1E5DDE3F",
    x"1E5D87A5",
    x"1E5D312D",
    x"1E5CDAD6",
    x"1E5C84A2",
    x"1E5C2E8F",
    x"1E5BD89D",
    x"1E5B82CD",
    x"1E5B2D1F",
    x"1E5AD792",
    x"1E5A8227",
    x"1E5A2CDC",
    x"1E59D7B4",
    x"1E5982AC",
    x"1E592DC5",
    x"1E58D900",
    x"1E58845C",
    x"1E582FD9",
    x"1E57DB77",
    x"1E578735",
    x"1E573315",
    x"1E56DF15",
    x"1E568B37",
    x"1E563779",
    x"1E55E3DB",
    x"1E55905F",
    x"1E553D02",
    x"1E54E9C7",
    x"1E5496AC",
    x"1E5443B1",
    x"1E53F0D7",
    x"1E539E1D",
    x"1E534B83",
    x"1E52F90A",
    x"1E52A6B1",
    x"1E525478",
    x"1E52025F",
    x"1E51B066",
    x"1E515E8D",
    x"1E510CD4",
    x"1E50BB3B",
    x"1E5069C2",
    x"1E501868",
    x"1E4FC72F",
    x"1E4F7615",
    x"1E4F251A",
    x"1E4ED440",
    x"1E4E8384",
    x"1E4E32E9",
    x"1E4DE26D",
    x"1E4D9210",
    x"1E4D41D3",
    x"1E4CF1B4",
    x"1E4CA1B6",
    x"1E4C51D6",
    x"1E4C0216",
    x"1E4BB274",
    x"1E4B62F2",
    x"1E4B138F",
    x"1E4AC44B",
    x"1E4A7526",
    x"1E4A261F",
    x"1E49D738",
    x"1E49886F",
    x"1E4939C5",
    x"1E48EB3A",
    x"1E489CCE",
    x"1E484E80",
    x"1E480050",
    x"1E47B23F",
    x"1E47644D",
    x"1E471679",
    x"1E46C8C3",
    x"1E467B2C",
    x"1E462DB3",
    x"1E45E058",
    x"1E45931C",
    x"1E4545FD",
    x"1E44F8FD",
    x"1E44AC1B",
    x"1E445F57",
    x"1E4412B0",
    x"1E43C628",
    x"1E4379BE",
    x"1E432D71",
    x"1E42E142",
    x"1E429531",
    x"1E42493E",
    x"1E41FD68",
    x"1E41B1B0",
    x"1E416615",
    x"1E411A98",
    x"1E40CF38",
    x"1E4083F6",
    x"1E4038D1",
    x"1E3FEDC9",
    x"1E3FA2DF",
    x"1E3F5812",
    x"1E3F0D62",
    x"1E3EC2D0",
    x"1E3E785A",
    x"1E3E2E02",
    x"1E3DE3C6",
    x"1E3D99A8",
    x"1E3D4FA6",
    x"1E3D05C2",
    x"1E3CBBFA",
    x"1E3C724F",
    x"1E3C28C0",
    x"1E3BDF4F",
    x"1E3B95FA",
    x"1E3B4CC2",
    x"1E3B03A6",
    x"1E3ABAA7",
    x"1E3A71C4",
    x"1E3A28FE",
    x"1E39E054",
    x"1E3997C7",
    x"1E394F55",
    x"1E390701",
    x"1E38BEC8",
    x"1E3876AC",
    x"1E382EAB",
    x"1E37E6C7",
    x"1E379EFF",
    x"1E375753",
    x"1E370FC3",
    x"1E36C84E",
    x"1E3680F6",
    x"1E3639BA",
    x"1E35F299",
    x"1E35AB94",
    x"1E3564AB",
    x"1E351DDE",
    x"1E34D72C",
    x"1E349095",
    x"1E344A1B",
    x"1E3403BB",
    x"1E33BD78",
    x"1E33774F",
    x"1E333143",
    x"1E32EB51",
    x"1E32A57B",
    x"1E325FC0",
    x"1E321A20",
    x"1E31D49B",
    x"1E318F32",
    x"1E3149E3",
    x"1E3104B0",
    x"1E30BF98",
    x"1E307A9A",
    x"1E3035B8",
    x"1E2FF0F0",
    x"1E2FAC44",
    x"1E2F67B2",
    x"1E2F233B",
    x"1E2EDEDE",
    x"1E2E9A9C",
    x"1E2E5675",
    x"1E2E1269",
    x"1E2DCE77",
    x"1E2D8AA0",
    x"1E2D46E3",
    x"1E2D0340",
    x"1E2CBFB8",
    x"1E2C7C4A",
    x"1E2C38F7",
    x"1E2BF5BE",
    x"1E2BB29F",
    x"1E2B6F9A",
    x"1E2B2CB0",
    x"1E2AE9DF",
    x"1E2AA729",
    x"1E2A648D",
    x"1E2A220B",
    x"1E29DFA2",
    x"1E299D54",
    x"1E295B1F",
    x"1E291905",
    x"1E28D704",
    x"1E28951D",
    x"1E28534F",
    x"1E28119C",
    x"1E27D001",
    x"1E278E81",
    x"1E274D1A",
    x"1E270BCD",
    x"1E26CA99",
    x"1E26897E",
    x"1E26487D",
    x"1E260796",
    x"1E25C6C8",
    x"1E258612",
    x"1E254577",
    x"1E2504F4",
    x"1E24C48B",
    x"1E24843B",
    x"1E244404",
    x"1E2403E6",
    x"1E23C3E0",
    x"1E2383F4",
    x"1E234421",
    x"1E230467",
    x"1E22C4C6",
    x"1E22853D",
    x"1E2245CE",
    x"1E220677",
    x"1E21C739",
    x"1E218813",
    x"1E214906",
    x"1E210A12",
    x"1E20CB37",
    x"1E208C73",
    x"1E204DC9",
    x"1E200F37",
    x"1E1FD0BD",
    x"1E1F925C",
    x"1E1F5413",
    x"1E1F15E2",
    x"1E1ED7C9",
    x"1E1E99C9",
    x"1E1E5BE1",
    x"1E1E1E11",
    x"1E1DE05A",
    x"1E1DA2BA",
    x"1E1D6533",
    x"1E1D27C3",
    x"1E1CEA6C",
    x"1E1CAD2C",
    x"1E1C7004",
    x"1E1C32F4",
    x"1E1BF5FC",
    x"1E1BB91C",
    x"1E1B7C54",
    x"1E1B3FA3",
    x"1E1B030A",
    x"1E1AC689",
    x"1E1A8A1F",
    x"1E1A4DCD",
    x"1E1A1192",
    x"1E19D56F",
    x"1E199963",
    x"1E195D6F",
    x"1E192192",
    x"1E18E5CD",
    x"1E18AA1F",
    x"1E186E88",
    x"1E183309",
    x"1E17F7A0",
    x"1E17BC4F",
    x"1E178115",
    x"1E1745F2",
    x"1E170AE6",
    x"1E16CFF2",
    x"1E169514",
    x"1E165A4D",
    x"1E161F9D",
    x"1E15E504",
    x"1E15AA82",
    x"1E157017",
    x"1E1535C3",
    x"1E14FB85",
    x"1E14C15E",
    x"1E14874E",
    x"1E144D55",
    x"1E141372",
    x"1E13D9A5",
    x"1E139FF0",
    x"1E136650",
    x"1E132CC8",
    x"1E12F355",
    x"1E12B9FA",
    x"1E1280B4",
    x"1E124785",
    x"1E120E6C",
    x"1E11D56A",
    x"1E119C7E",
    x"1E1163A8",
    x"1E112AE8",
    x"1E10F23E",
    x"1E10B9AA",
    x"1E10812D",
    x"1E1048C5",
    x"1E101074",
    x"1E0FD839",
    x"1E0FA013",
    x"1E0F6804",
    x"1E0F300A",
    x"1E0EF826",
    x"1E0EC058",
    x"1E0E88A0",
    x"1E0E50FD",
    x"1E0E1970",
    x"1E0DE1F9",
    x"1E0DAA98",
    x"1E0D734C",
    x"1E0D3C16",
    x"1E0D04F5",
    x"1E0CCDEA",
    x"1E0C96F4",
    x"1E0C6014",
    x"1E0C2949",
    x"1E0BF294",
    x"1E0BBBF4",
    x"1E0B8569",
    x"1E0B4EF3",
    x"1E0B1893",
    x"1E0AE248",
    x"1E0AAC12",
    x"1E0A75F2",
    x"1E0A3FE6",
    x"1E0A09F0",
    x"1E09D40E",
    x"1E099E42",
    x"1E09688B",
    x"1E0932E8",
    x"1E08FD5B",
    x"1E08C7E2",
    x"1E08927F",
    x"1E085D30",
    x"1E0827F6",
    x"1E07F2D1",
    x"1E07BDC0",
    x"1E0788C5",
    x"1E0753DD",
    x"1E071F0B",
    x"1E06EA4D",
    x"1E06B5A4",
    x"1E06810F",
    x"1E064C8F",
    x"1E061823",
    x"1E05E3CC",
    x"1E05AF89",
    x"1E057B5B",
    x"1E054741",
    x"1E05133B",
    x"1E04DF4A",
    x"1E04AB6D",
    x"1E0477A4",
    x"1E0443EF",
    x"1E04104F",
    x"1E03DCC3",
    x"1E03A94B",
    x"1E0375E6",
    x"1E034296",
    x"1E030F5A",
    x"1E02DC32",
    x"1E02A91E",
    x"1E02761E",
    x"1E024332",
    x"1E02105A",
    x"1E01DD95",
    x"1E01AAE5",
    x"1E017848",
    x"1E0145BF",
    x"1E011349",
    x"1E00E0E8",
    x"1E00AE9A",
    x"1E007C5F",
    x"1E004A38",
    x"1E001825",
    x"1DFFCC4B",
    x"1DFF6873",
    x"1DFF04C1",
    x"1DFEA137",
    x"1DFE3DD3",
    x"1DFDDA97",
    x"1DFD7781",
    x"1DFD1491",
    x"1DFCB1C9",
    x"1DFC4F26",
    x"1DFBECAB",
    x"1DFB8A56",
    x"1DFB2827",
    x"1DFAC61E",
    x"1DFA643C",
    x"1DFA0280",
    x"1DF9A0EA",
    x"1DF93F7A",
    x"1DF8DE30",
    x"1DF87D0C",
    x"1DF81C0F",
    x"1DF7BB37",
    x"1DF75A84",
    x"1DF6F9F8",
    x"1DF69991",
    x"1DF63950",
    x"1DF5D934",
    x"1DF5793E",
    x"1DF5196D",
    x"1DF4B9C2",
    x"1DF45A3C",
    x"1DF3FADC",
    x"1DF39BA0",
    x"1DF33C8A",
    x"1DF2DD99",
    x"1DF27ECD",
    x"1DF22026",
    x"1DF1C1A4",
    x"1DF16347",
    x"1DF1050E",
    x"1DF0A6FB",
    x"1DF0490C",
    x"1DEFEB42",
    x"1DEF8D9C",
    x"1DEF301B",
    x"1DEED2BE",
    x"1DEE7586",
    x"1DEE1873",
    x"1DEDBB83",
    x"1DED5EB8",
    x"1DED0211",
    x"1DECA58E",
    x"1DEC4930",
    x"1DEBECF5",
    x"1DEB90DF",
    x"1DEB34EC",
    x"1DEAD91D",
    x"1DEA7D72",
    x"1DEA21EB",
    x"1DE9C688",
    x"1DE96B48",
    x"1DE9102C",
    x"1DE8B533",
    x"1DE85A5E",
    x"1DE7FFAD",
    x"1DE7A51F",
    x"1DE74AB4",
    x"1DE6F06C",
    x"1DE69648",
    x"1DE63C47",
    x"1DE5E269",
    x"1DE588AE",
    x"1DE52F16",
    x"1DE4D5A1",
    x"1DE47C4F",
    x"1DE42320",
    x"1DE3CA14",
    x"1DE3712A",
    x"1DE31863",
    x"1DE2BFBF",
    x"1DE2673D",
    x"1DE20EDE",
    x"1DE1B6A2",
    x"1DE15E88",
    x"1DE10690",
    x"1DE0AEBB",
    x"1DE05707",
    x"1DDFFF77",
    x"1DDFA808",
    x"1DDF50BB",
    x"1DDEF991",
    x"1DDEA288",
    x"1DDE4BA2",
    x"1DDDF4DD",
    x"1DDD9E3A",
    x"1DDD47B9",
    x"1DDCF15A",
    x"1DDC9B1D",
    x"1DDC4501",
    x"1DDBEF07",
    x"1DDB992E",
    x"1DDB4377",
    x"1DDAEDE2",
    x"1DDA986D",
    x"1DDA431B",
    x"1DD9EDE9",
    x"1DD998D9",
    x"1DD943EA",
    x"1DD8EF1C",
    x"1DD89A6F",
    x"1DD845E3",
    x"1DD7F178",
    x"1DD79D2E",
    x"1DD74905",
    x"1DD6F4FD",
    x"1DD6A116",
    x"1DD64D4F",
    x"1DD5F9A9",
    x"1DD5A624",
    x"1DD552C0",
    x"1DD4FF7C",
    x"1DD4AC58",
    x"1DD45955",
    x"1DD40672",
    x"1DD3B3B0",
    x"1DD3610E",
    x"1DD30E8C",
    x"1DD2BC2A",
    x"1DD269E9",
    x"1DD217C8",
    x"1DD1C5C6",
    x"1DD173E5",
    x"1DD12224",
    x"1DD0D083",
    x"1DD07F01",
    x"1DD02D9F",
    x"1DCFDC5D",
    x"1DCF8B3B",
    x"1DCF3A39",
    x"1DCEE956",
    x"1DCE9892",
    x"1DCE47EE",
    x"1DCDF76A",
    x"1DCDA705",
    x"1DCD56C0",
    x"1DCD0699",
    x"1DCCB692",
    x"1DCC66AB",
    x"1DCC16E2",
    x"1DCBC739",
    x"1DCB77AE",
    x"1DCB2843",
    x"1DCAD8F7",
    x"1DCA89CA",
    x"1DCA3ABB",
    x"1DC9EBCC",
    x"1DC99CFB",
    x"1DC94E49",
    x"1DC8FFB6",
    x"1DC8B141",
    x"1DC862EB",
    x"1DC814B4",
    x"1DC7C69B",
    x"1DC778A1",
    x"1DC72AC5",
    x"1DC6DD07",
    x"1DC68F68",
    x"1DC641E7",
    x"1DC5F485",
    x"1DC5A740",
    x"1DC55A1A",
    x"1DC50D12",
    x"1DC4C028",
    x"1DC4735C",
    x"1DC426AE",
    x"1DC3DA1E",
    x"1DC38DAB",
    x"1DC34157",
    x"1DC2F520",
    x"1DC2A907",
    x"1DC25D0C",
    x"1DC2112F",
    x"1DC1C56F",
    x"1DC179CC",
    x"1DC12E48",
    x"1DC0E2E0",
    x"1DC09796",
    x"1DC04C6A",
    x"1DC0015B",
    x"1DBFB669",
    x"1DBF6B94",
    x"1DBF20DD",
    x"1DBED642",
    x"1DBE8BC5",
    x"1DBE4165",
    x"1DBDF722",
    x"1DBDACFC",
    x"1DBD62F3",
    x"1DBD1907",
    x"1DBCCF37",
    x"1DBC8585",
    x"1DBC3BEF",
    x"1DBBF276",
    x"1DBBA91A",
    x"1DBB5FDA",
    x"1DBB16B7",
    x"1DBACDB0",
    x"1DBA84C6",
    x"1DBA3BF8",
    x"1DB9F347",
    x"1DB9AAB2",
    x"1DB9623A",
    x"1DB919DE",
    x"1DB8D19E",
    x"1DB8897A",
    x"1DB84172",
    x"1DB7F987",
    x"1DB7B1B7",
    x"1DB76A04",
    x"1DB7226C",
    x"1DB6DAF1",
    x"1DB69391",
    x"1DB64C4E",
    x"1DB60526",
    x"1DB5BE1A",
    x"1DB57729",
    x"1DB53054",
    x"1DB4E99B",
    x"1DB4A2FE",
    x"1DB45C7C",
    x"1DB41616",
    x"1DB3CFCB",
    x"1DB3899B",
    x"1DB34387",
    x"1DB2FD8F",
    x"1DB2B7B1",
    x"1DB271EF",
    x"1DB22C48",
    x"1DB1E6BC",
    x"1DB1A14C",
    x"1DB15BF6",
    x"1DB116BC",
    x"1DB0D19D",
    x"1DB08C98",
    x"1DB047AF",
    x"1DB002E0",
    x"1DAFBE2C",
    x"1DAF7994",
    x"1DAF3515",
    x"1DAEF0B2",
    x"1DAEAC69",
    x"1DAE683B",
    x"1DAE2428",
    x"1DADE02F",
    x"1DAD9C51",
    x"1DAD588D",
    x"1DAD14E4",
    x"1DACD155",
    x"1DAC8DE0",
    x"1DAC4A86",
    x"1DAC0746",
    x"1DABC420",
    x"1DAB8115",
    x"1DAB3E23",
    x"1DAAFB4C",
    x"1DAAB88F",
    x"1DAA75EC",
    x"1DAA3363",
    x"1DA9F0F4",
    x"1DA9AE9F",
    x"1DA96C63",
    x"1DA92A42",
    x"1DA8E83A",
    x"1DA8A64C",
    x"1DA86478",
    x"1DA822BE",
    x"1DA7E11D",
    x"1DA79F96",
    x"1DA75E28",
    x"1DA71CD4",
    x"1DA6DB9A",
    x"1DA69A79",
    x"1DA65971",
    x"1DA61883",
    x"1DA5D7AE",
    x"1DA596F2",
    x"1DA55650",
    x"1DA515C7",
    x"1DA4D557",
    x"1DA49500",
    x"1DA454C3",
    x"1DA4149E",
    x"1DA3D493",
    x"1DA394A0",
    x"1DA354C6",
    x"1DA31506",
    x"1DA2D55E",
    x"1DA295CF",
    x"1DA25659",
    x"1DA216FC",
    x"1DA1D7B7",
    x"1DA1988B",
    x"1DA15978",
    x"1DA11A7D",
    x"1DA0DB9B",
    x"1DA09CD2",
    x"1DA05E21",
    x"1DA01F88",
    x"1D9FE108",
    x"1D9FA2A0",
    x"1D9F6451",
    x"1D9F261A",
    x"1D9EE7FB",
    x"1D9EA9F5",
    x"1D9E6C06",
    x"1D9E2E30",
    x"1D9DF072",
    x"1D9DB2CC",
    x"1D9D753E",
    x"1D9D37C9",
    x"1D9CFA6B",
    x"1D9CBD25",
    x"1D9C7FF7",
    x"1D9C42E1",
    x"1D9C05E3",
    x"1D9BC8FC",
    x"1D9B8C2E",
    x"1D9B4F77",
    x"1D9B12D8",
    x"1D9AD650",
    x"1D9A99E0",
    x"1D9A5D88",
    x"1D9A2147",
    x"1D99E51E",
    x"1D99A90C",
    x"1D996D12",
    x"1D99312F",
    x"1D98F563",
    x"1D98B9AF",
    x"1D987E12",
    x"1D98428D",
    x"1D98071E",
    x"1D97CBC7",
    x"1D979087",
    x"1D97555E",
    x"1D971A4C",
    x"1D96DF52",
    x"1D96A46E",
    x"1D9669A1",
    x"1D962EEB",
    x"1D95F44D",
    x"1D95B9C5",
    x"1D957F53",
    x"1D9544F9",
    x"1D950AB6",
    x"1D94D089",
    x"1D949673",
    x"1D945C73",
    x"1D94228A",
    x"1D93E8B8",
    x"1D93AEFD",
    x"1D937557",
    x"1D933BC9",
    x"1D930251",
    x"1D92C8EF",
    x"1D928FA4",
    x"1D92566F",
    x"1D921D50",
    x"1D91E448",
    x"1D91AB56",
    x"1D91727A",
    x"1D9139B4",
    x"1D910105",
    x"1D90C86C",
    x"1D908FE8",
    x"1D90577B",
    x"1D901F24",
    x"1D8FE6E3",
    x"1D8FAEB8",
    x"1D8F76A2",
    x"1D8F3EA3",
    x"1D8F06B9",
    x"1D8ECEE6",
    x"1D8E9728",
    x"1D8E5F80",
    x"1D8E27ED",
    x"1D8DF070",
    x"1D8DB909",
    x"1D8D81B8",
    x"1D8D4A7C",
    x"1D8D1356",
    x"1D8CDC45",
    x"1D8CA549",
    x"1D8C6E64",
    x"1D8C3793",
    x"1D8C00D8",
    x"1D8BCA33",
    x"1D8B93A2",
    x"1D8B5D27",
    x"1D8B26C1",
    x"1D8AF071",
    x"1D8ABA36",
    x"1D8A840F",
    x"1D8A4DFE",
    x"1D8A1802",
    x"1D89E21C",
    x"1D89AC4A",
    x"1D89768D",
    x"1D8940E5",
    x"1D890B52",
    x"1D88D5D4",
    x"1D88A06B",
    x"1D886B17",
    x"1D8835D8",
    x"1D8800AD",
    x"1D87CB97",
    x"1D879696",
    x"1D8761A9",
    x"1D872CD2",
    x"1D86F80E",
    x"1D86C360",
    x"1D868EC6",
    x"1D865A40",
    x"1D8625CF",
    x"1D85F173",
    x"1D85BD2B",
    x"1D8588F7",
    x"1D8554D8",
    x"1D8520CD",
    x"1D84ECD6",
    x"1D84B8F3",
    x"1D848525",
    x"1D84516B",
    x"1D841DC6",
    x"1D83EA34",
    x"1D83B6B7",
    x"1D83834D",
    x"1D834FF8",
    x"1D831CB7",
    x"1D82E98A",
    x"1D82B670",
    x"1D82836B",
    x"1D82507A",
    x"1D821D9C",
    x"1D81EAD3",
    x"1D81B81D",
    x"1D81857B",
    x"1D8152ED",
    x"1D812072",
    x"1D80EE0B",
    x"1D80BBB8",
    x"1D808979",
    x"1D80574D",
    x"1D802534",
    x"1D7FE65F",
    x"1D7F827D",
    x"1D7F1EC1",
    x"1D7EBB2D",
    x"1D7E57BF",
    x"1D7DF478",
    x"1D7D9158",
    x"1D7D2E5E",
    x"1D7CCB8C",
    x"1D7C68DF",
    x"1D7C065A",
    x"1D7BA3FA",
    x"1D7B41C2",
    x"1D7ADFAF",
    x"1D7A7DC3",
    x"1D7A1BFD",
    x"1D79BA5D",
    x"1D7958E3",
    x"1D78F78F",
    x"1D789662",
    x"1D78355A",
    x"1D77D478",
    x"1D7773BC",
    x"1D771326",
    x"1D76B2B5",
    x"1D76526A",
    x"1D75F245",
    x"1D759245",
    x"1D75326A",
    x"1D74D2B5",
    x"1D747326",
    x"1D7413BB",
    x"1D73B476",
    x"1D735556",
    x"1D72F65B",
    x"1D729786",
    x"1D7238D5",
    x"1D71DA49",
    x"1D717BE3",
    x"1D711DA1",
    x"1D70BF83",
    x"1D70618B",
    x"1D7003B7",
    x"1D6FA608",
    x"1D6F487D",
    x"1D6EEB17",
    x"1D6E8DD6",
    x"1D6E30B9",
    x"1D6DD3C0",
    x"1D6D76EB",
    x"1D6D1A3B",
    x"1D6CBDAF",
    x"1D6C6147",
    x"1D6C0503",
    x"1D6BA8E3",
    x"1D6B4CE7",
    x"1D6AF10F",
    x"1D6A955A",
    x"1D6A39CA",
    x"1D69DE5D",
    x"1D698314",
    x"1D6927EF",
    x"1D68CCED",
    x"1D68720F",
    x"1D681754",
    x"1D67BCBC",
    x"1D676248",
    x"1D6707F8",
    x"1D66ADCA",
    x"1D6653C0",
    x"1D65F9D9",
    x"1D65A015",
    x"1D654673",
    x"1D64ECF5",
    x"1D64939A",
    x"1D643A62",
    x"1D63E14D",
    x"1D63885A",
    x"1D632F8A",
    x"1D62D6DD",
    x"1D627E52",
    x"1D6225EA",
    x"1D61CDA5",
    x"1D617582",
    x"1D611D81",
    x"1D60C5A2",
    x"1D606DE6",
    x"1D60164D",
    x"1D5FBED5",
    x"1D5F677F",
    x"1D5F104C",
    x"1D5EB93B",
    x"1D5E624B",
    x"1D5E0B7E",
    x"1D5DB4D2",
    x"1D5D5E49",
    x"1D5D07E1",
    x"1D5CB19A",
    x"1D5C5B76",
    x"1D5C0573",
    x"1D5BAF92",
    x"1D5B59D2",
    x"1D5B0433",
    x"1D5AAEB7",
    x"1D5A595B",
    x"1D5A0421",
    x"1D59AF08",
    x"1D595A10",
    x"1D590539",
    x"1D58B084",
    x"1D585BEF",
    x"1D58077C",
    x"1D57B32A",
    x"1D575EF8",
    x"1D570AE7",
    x"1D56B6F7",
    x"1D566328",
    x"1D560F7A",
    x"1D55BBEC",
    x"1D55687F",
    x"1D551533",
    x"1D54C207",
    x"1D546EFB",
    x"1D541C10",
    x"1D53C945",
    x"1D53769B",
    x"1D532410",
    x"1D52D1A6",
    x"1D527F5D",
    x"1D522D33",
    x"1D51DB29",
    x"1D518940",
    x"1D513776",
    x"1D50E5CC",
    x"1D509442",
    x"1D5042D8",
    x"1D4FF18E",
    x"1D4FA064",
    x"1D4F4F59",
    x"1D4EFE6E",
    x"1D4EADA2",
    x"1D4E5CF6",
    x"1D4E0C69",
    x"1D4DBBFC",
    x"1D4D6BAF",
    x"1D4D1B80",
    x"1D4CCB71",
    x"1D4C7B81",
    x"1D4C2BB1",
    x"1D4BDBFF",
    x"1D4B8C6D",
    x"1D4B3CF9",
    x"1D4AEDA5",
    x"1D4A9E70",
    x"1D4A4F59",
    x"1D4A0062",
    x"1D49B189",
    x"1D4962CF",
    x"1D491434",
    x"1D48C5B7",
    x"1D487759",
    x"1D48291A",
    x"1D47DAF9",
    x"1D478CF7",
    x"1D473F13",
    x"1D46F14E",
    x"1D46A3A6",
    x"1D46561E",
    x"1D4608B3",
    x"1D45BB67",
    x"1D456E39",
    x"1D452129",
    x"1D44D437",
    x"1D448763",
    x"1D443AAD",
    x"1D43EE15",
    x"1D43A19B",
    x"1D43553F",
    x"1D430900",
    x"1D42BCE0",
    x"1D4270DD",
    x"1D4224F8",
    x"1D41D930",
    x"1D418D86",
    x"1D4141F9",
    x"1D40F68A",
    x"1D40AB39",
    x"1D406005",
    x"1D4014EE",
    x"1D3FC9F4",
    x"1D3F7F18",
    x"1D3F3459",
    x"1D3EE9B7",
    x"1D3E9F32",
    x"1D3E54CB",
    x"1D3E0A80",
    x"1D3DC052",
    x"1D3D7642",
    x"1D3D2C4E",
    x"1D3CE277",
    x"1D3C98BD",
    x"1D3C4F20",
    x"1D3C059F",
    x"1D3BBC3B",
    x"1D3B72F4",
    x"1D3B29CA",
    x"1D3AE0BB",
    x"1D3A97CA",
    x"1D3A4EF5",
    x"1D3A063C",
    x"1D39BDA0",
    x"1D397520",
    x"1D392CBC",
    x"1D38E475",
    x"1D389C4A",
    x"1D38543B",
    x"1D380C48",
    x"1D37C471",
    x"1D377CB7",
    x"1D373518",
    x"1D36ED95",
    x"1D36A62E",
    x"1D365EE3",
    x"1D3617B4",
    x"1D35D0A1",
    x"1D3589A9",
    x"1D3542CD",
    x"1D34FC0D",
    x"1D34B568",
    x"1D346EDF",
    x"1D342872",
    x"1D33E220",
    x"1D339BE9",
    x"1D3355CE",
    x"1D330FCE",
    x"1D32C9E9",
    x"1D328420",
    x"1D323E72",
    x"1D31F8DF",
    x"1D31B368",
    x"1D316E0B",
    x"1D3128CA",
    x"1D30E3A3",
    x"1D309E98",
    x"1D3059A7",
    x"1D3014D2",
    x"1D2FD017",
    x"1D2F8B77",
    x"1D2F46F2",
    x"1D2F0288",
    x"1D2EBE38",
    x"1D2E7A03",
    x"1D2E35E9",
    x"1D2DF1E9",
    x"1D2DAE04",
    x"1D2D6A39",
    x"1D2D2689",
    x"1D2CE2F3",
    x"1D2C9F78",
    x"1D2C5C16",
    x"1D2C18D0",
    x"1D2BD5A3",
    x"1D2B9291",
    x"1D2B4F99",
    x"1D2B0CBA",
    x"1D2AC9F7",
    x"1D2A874D",
    x"1D2A44BD",
    x"1D2A0247",
    x"1D29BFEB",
    x"1D297DA9",
    x"1D293B81",
    x"1D28F973",
    x"1D28B77E",
    x"1D2875A3",
    x"1D2833E2",
    x"1D27F23B",
    x"1D27B0AD",
    x"1D276F39",
    x"1D272DDE",
    x"1D26EC9D",
    x"1D26AB75",
    x"1D266A67",
    x"1D262972",
    x"1D25E896",
    x"1D25A7D4",
    x"1D25672B",
    x"1D25269C",
    x"1D24E625",
    x"1D24A5C8",
    x"1D246584",
    x"1D242558",
    x"1D23E546",
    x"1D23A54D",
    x"1D23656D",
    x"1D2325A6",
    x"1D22E5F8",
    x"1D22A662",
    x"1D2266E6",
    x"1D222782",
    x"1D21E837",
    x"1D21A905",
    x"1D2169EB",
    x"1D212AEA",
    x"1D20EC01",
    x"1D20AD31",
    x"1D206E7A",
    x"1D202FDB",
    x"1D1FF155",
    x"1D1FB2E6",
    x"1D1F7491",
    x"1D1F3653",
    x"1D1EF82E",
    x"1D1EBA22",
    x"1D1E7C2D",
    x"1D1E3E50",
    x"1D1E008C",
    x"1D1DC2E0",
    x"1D1D854C",
    x"1D1D47D0",
    x"1D1D0A6C",
    x"1D1CCD20",
    x"1D1C8FEC",
    x"1D1C52CF",
    x"1D1C15CB",
    x"1D1BD8DE",
    x"1D1B9C09",
    x"1D1B5F4C",
    x"1D1B22A7",
    x"1D1AE619",
    x"1D1AA9A3",
    x"1D1A6D45",
    x"1D1A30FE",
    x"1D19F4CE",
    x"1D19B8B7",
    x"1D197CB6",
    x"1D1940CD",
    x"1D1904FB",
    x"1D18C941",
    x"1D188D9E",
    x"1D185213",
    x"1D18169E",
    x"1D17DB41",
    x"1D179FFB",
    x"1D1764CC",
    x"1D1729B4",
    x"1D16EEB3",
    x"1D16B3CA",
    x"1D1678F7",
    x"1D163E3B",
    x"1D160396",
    x"1D15C908",
    x"1D158E91",
    x"1D155431",
    x"1D1519E7",
    x"1D14DFB5",
    x"1D14A599",
    x"1D146B93",
    x"1D1431A4",
    x"1D13F7CC",
    x"1D13BE0B",
    x"1D138460",
    x"1D134ACB",
    x"1D13114D",
    x"1D12D7E6",
    x"1D129E95",
    x"1D12655A",
    x"1D122C36",
    x"1D11F327",
    x"1D11BA30",
    x"1D11814E",
    x"1D114883",
    x"1D110FCD",
    x"1D10D72E",
    x"1D109EA5",
    x"1D106632",
    x"1D102DD5",
    x"1D0FF58E",
    x"1D0FBD5E",
    x"1D0F8543",
    x"1D0F4D3D",
    x"1D0F154E",
    x"1D0EDD75",
    x"1D0EA5B1",
    x"1D0E6E03",
    x"1D0E366B",
    x"1D0DFEE9",
    x"1D0DC77C",
    x"1D0D9025",
    x"1D0D58E3",
    x"1D0D21B7",
    x"1D0CEAA1",
    x"1D0CB3A0",
    x"1D0C7CB5",
    x"1D0C45DF",
    x"1D0C0F1E",
    x"1D0BD873",
    x"1D0BA1DD",
    x"1D0B6B5C",
    x"1D0B34F1",
    x"1D0AFE9B",
    x"1D0AC85A",
    x"1D0A922E",
    x"1D0A5C18",
    x"1D0A2617",
    x"1D09F02A",
    x"1D09BA53",
    x"1D098491",
    x"1D094EE3",
    x"1D09194B",
    x"1D08E3C8",
    x"1D08AE59",
    x"1D0878FF",
    x"1D0843BA",
    x"1D080E8A",
    x"1D07D96F",
    x"1D07A469",
    x"1D076F77",
    x"1D073A99",
    x"1D0705D1",
    x"1D06D11D",
    x"1D069C7D",
    x"1D0667F3",
    x"1D06337C",
    x"1D05FF1A",
    x"1D05CACD",
    x"1D059694",
    x"1D05626F",
    x"1D052E5F",
    x"1D04FA63",
    x"1D04C67B",
    x"1D0492A8",
    x"1D045EE9",
    x"1D042B3E",
    x"1D03F7A7",
    x"1D03C424",
    x"1D0390B6",
    x"1D035D5B",
    x"1D032A15",
    x"1D02F6E2",
    x"1D02C3C4",
    x"1D0290B9",
    x"1D025DC3",
    x"1D022AE0",
    x"1D01F811",
    x"1D01C556",
    x"1D0192AF",
    x"1D01601C",
    x"1D012D9C",
    x"1D00FB30",
    x"1D00C8D8",
    x"1D009693",
    x"1D006462",
    x"1D003245",
    x"1D00003B",
    x"1CFF9C89",
    x"1CFF38C3",
    x"1CFED525",
    x"1CFE71AD",
    x"1CFE0E5C",
    x"1CFDAB32",
    x"1CFD482E",
    x"1CFCE551",
    x"1CFC829B",
    x"1CFC200B",
    x"1CFBBDA2",
    x"1CFB5B5F",
    x"1CFAF943",
    x"1CFA974C",
    x"1CFA357C",
    x"1CF9D3D3",
    x"1CF9724F",
    x"1CF910F1",
    x"1CF8AFBA",
    x"1CF84EA8",
    x"1CF7EDBC",
    x"1CF78CF6",
    x"1CF72C56",
    x"1CF6CBDB",
    x"1CF66B87",
    x"1CF60B57",
    x"1CF5AB4E",
    x"1CF54B6A",
    x"1CF4EBAB",
    x"1CF48C11",
    x"1CF42C9D",
    x"1CF3CD4F",
    x"1CF36E25",
    x"1CF30F21",
    x"1CF2B041",
    x"1CF25187",
    x"1CF1F2F1",
    x"1CF19481",
    x"1CF13635",
    x"1CF0D80F",
    x"1CF07A0D",
    x"1CF01C2F",
    x"1CEFBE77",
    x"1CEF60E2",
    x"1CEF0373",
    x"1CEEA628",
    x"1CEE4901",
    x"1CEDEBFF",
    x"1CED8F21",
    x"1CED3267",
    x"1CECD5D1",
    x"1CEC7960",
    x"1CEC1D12",
    x"1CEBC0E9",
    x"1CEB64E4",
    x"1CEB0902",
    x"1CEAAD45",
    x"1CEA51AB",
    x"1CE9F635",
    x"1CE99AE2",
    x"1CE93FB4",
    x"1CE8E4A9",
    x"1CE889C1",
    x"1CE82EFD",
    x"1CE7D45C",
    x"1CE779DF",
    x"1CE71F85",
    x"1CE6C54E",
    x"1CE66B3B",
    x"1CE6114B",
    x"1CE5B77D",
    x"1CE55DD3",
    x"1CE5044C",
    x"1CE4AAE8",
    x"1CE451A7",
    x"1CE3F888",
    x"1CE39F8C",
    x"1CE346B3",
    x"1CE2EDFD",
    x"1CE2956A",
    x"1CE23CF8",
    x"1CE1E4AA",
    x"1CE18C7E",
    x"1CE13474",
    x"1CE0DC8D",
    x"1CE084C8",
    x"1CE02D25",
    x"1CDFD5A4",
    x"1CDF7E46",
    x"1CDF270A",
    x"1CDECFF0",
    x"1CDE78F7",
    x"1CDE2221",
    x"1CDDCB6D",
    x"1CDD74DA",
    x"1CDD1E69",
    x"1CDCC81A",
    x"1CDC71ED",
    x"1CDC1BE1",
    x"1CDBC5F7",
    x"1CDB702F",
    x"1CDB1A88",
    x"1CDAC502",
    x"1CDA6F9E",
    x"1CDA1A5B",
    x"1CD9C539",
    x"1CD97039",
    x"1CD91B59",
    x"1CD8C69B",
    x"1CD871FE",
    x"1CD81D82",
    x"1CD7C927",
    x"1CD774ED",
    x"1CD720D4",
    x"1CD6CCDB",
    x"1CD67904",
    x"1CD6254D",
    x"1CD5D1B6",
    x"1CD57E41",
    x"1CD52AEC",
    x"1CD4D7B7",
    x"1CD484A3",
    x"1CD431B0",
    x"1CD3DEDC",
    x"1CD38C2A",
    x"1CD33997",
    x"1CD2E725",
    x"1CD294D2",
    x"1CD242A0",
    x"1CD1F08E",
    x"1CD19E9C",
    x"1CD14CCA",
    x"1CD0FB18",
    x"1CD0A986",
    x"1CD05814",
    x"1CD006C1",
    x"1CCFB58F",
    x"1CCF647B",
    x"1CCF1388",
    x"1CCEC2B4",
    x"1CCE7200",
    x"1CCE216B",
    x"1CCDD0F6",
    x"1CCD80A0",
    x"1CCD3069",
    x"1CCCE052",
    x"1CCC905A",
    x"1CCC4081",
    x"1CCBF0C8",
    x"1CCBA12D",
    x"1CCB51B2",
    x"1CCB0255",
    x"1CCAB318",
    x"1CCA63F9",
    x"1CCA14FA",
    x"1CC9C619",
    x"1CC97757",
    x"1CC928B4",
    x"1CC8DA2F",
    x"1CC88BC9",
    x"1CC83D82",
    x"1CC7EF59",
    x"1CC7A14F",
    x"1CC75363",
    x"1CC70596",
    x"1CC6B7E7",
    x"1CC66A56",
    x"1CC61CE4",
    x"1CC5CF8F",
    x"1CC58259",
    x"1CC53542",
    x"1CC4E848",
    x"1CC49B6C",
    x"1CC44EAE",
    x"1CC4020F",
    x"1CC3B58D",
    x"1CC36929",
    x"1CC31CE3",
    x"1CC2D0BA",
    x"1CC284B0",
    x"1CC238C3",
    x"1CC1ECF3",
    x"1CC1A141",
    x"1CC155AD",
    x"1CC10A36",
    x"1CC0BEDD",
    x"1CC073A1",
    x"1CC02883",
    x"1CBFDD82",
    x"1CBF929E",
    x"1CBF47D7",
    x"1CBEFD2E",
    x"1CBEB2A1",
    x"1CBE6832",
    x"1CBE1DE0",
    x"1CBDD3AB",
    x"1CBD8992",
    x"1CBD3F97",
    x"1CBCF5B9",
    x"1CBCABF7",
    x"1CBC6252",
    x"1CBC18CA",
    x"1CBBCF5F",
    x"1CBB8610",
    x"1CBB3CDE",
    x"1CBAF3C9",
    x"1CBAAAD0",
    x"1CBA61F3",
    x"1CBA1933",
    x"1CB9D090",
    x"1CB98808",
    x"1CB93F9D",
    x"1CB8F74F",
    x"1CB8AF1C",
    x"1CB86706",
    x"1CB81F0C",
    x"1CB7D72E",
    x"1CB78F6B",
    x"1CB747C5",
    x"1CB7003B",
    x"1CB6B8CD",
    x"1CB6717B",
    x"1CB62A45",
    x"1CB5E32A",
    x"1CB59C2B",
    x"1CB55548",
    x"1CB50E80",
    x"1CB4C7D5",
    x"1CB48144",
    x"1CB43AD0",
    x"1CB3F476",
    x"1CB3AE39",
    x"1CB36816",
    x"1CB3220F",
    x"1CB2DC24",
    x"1CB29653",
    x"1CB2509E",
    x"1CB20B04",
    x"1CB1C586",
    x"1CB18022",
    x"1CB13AD9",
    x"1CB0F5AC",
    x"1CB0B099",
    x"1CB06BA2",
    x"1CB026C5",
    x"1CAFE204",
    x"1CAF9D5D",
    x"1CAF58D1",
    x"1CAF145F",
    x"1CAED009",
    x"1CAE8BCD",
    x"1CAE47AC",
    x"1CAE03A5",
    x"1CADBFB9",
    x"1CAD7BE7",
    x"1CAD3830",
    x"1CACF493",
    x"1CACB111",
    x"1CAC6DA9",
    x"1CAC2A5B",
    x"1CABE728",
    x"1CABA40F",
    x"1CAB6110",
    x"1CAB1E2B",
    x"1CAADB60",
    x"1CAA98AF",
    x"1CAA5619",
    x"1CAA139C",
    x"1CA9D139",
    x"1CA98EF1",
    x"1CA94CC2",
    x"1CA90AAD",
    x"1CA8C8B1",
    x"1CA886D0",
    x"1CA84508",
    x"1CA8035A",
    x"1CA7C1C5",
    x"1CA7804A",
    x"1CA73EE9",
    x"1CA6FDA1",
    x"1CA6BC73",
    x"1CA67B5E",
    x"1CA63A63",
    x"1CA5F980",
    x"1CA5B8B8",
    x"1CA57808",
    x"1CA53772",
    x"1CA4F6F5",
    x"1CA4B691",
    x"1CA47646",
    x"1CA43614",
    x"1CA3F5FC",
    x"1CA3B5FC",
    x"1CA37616",
    x"1CA33648",
    x"1CA2F693",
    x"1CA2B6F7",
    x"1CA27774",
    x"1CA2380A",
    x"1CA1F8B8",
    x"1CA1B980",
    x"1CA17A60",
    x"1CA13B58",
    x"1CA0FC69",
    x"1CA0BD93",
    x"1CA07ED5",
    x"1CA04030",
    x"1CA001A3",
    x"1C9FC32E",
    x"1C9F84D2",
    x"1C9F468F",
    x"1C9F0863",
    x"1C9ECA50",
    x"1C9E8C55",
    x"1C9E4E72",
    x"1C9E10A8",
    x"1C9DD2F5",
    x"1C9D955B",
    x"1C9D57D9",
    x"1C9D1A6E",
    x"1C9CDD1C",
    x"1C9C9FE2",
    x"1C9C62BF",
    x"1C9C25B5",
    x"1C9BE8C2",
    x"1C9BABE7",
    x"1C9B6F23",
    x"1C9B3278",
    x"1C9AF5E4",
    x"1C9AB968",
    x"1C9A7D03",
    x"1C9A40B6",
    x"1C9A0481",
    x"1C99C862",
    x"1C998C5C",
    x"1C99506D",
    x"1C991495",
    x"1C98D8D5",
    x"1C989D2C",
    x"1C98619A",
    x"1C98261F",
    x"1C97EABC",
    x"1C97AF70",
    x"1C97743B",
    x"1C97391D",
    x"1C96FE16",
    x"1C96C327",
    x"1C96884E",
    x"1C964D8C",
    x"1C9612E1",
    x"1C95D84D",
    x"1C959DD0",
    x"1C95636A",
    x"1C95291B",
    x"1C94EEE2",
    x"1C94B4C0",
    x"1C947AB5",
    x"1C9440C0",
    x"1C9406E2",
    x"1C93CD1B",
    x"1C93936A",
    x"1C9359D0",
    x"1C93204C",
    x"1C92E6DE",
    x"1C92AD87",
    x"1C927447",
    x"1C923B1D",
    x"1C920209",
    x"1C91C90B",
    x"1C919024",
    x"1C915752",
    x"1C911E97",
    x"1C90E5F2",
    x"1C90AD64",
    x"1C9074EB",
    x"1C903C88",
    x"1C90043C",
    x"1C8FCC05",
    x"1C8F93E4",
    x"1C8F5BD9",
    x"1C8F23E4",
    x"1C8EEC05",
    x"1C8EB43C",
    x"1C8E7C89",
    x"1C8E44EB",
    x"1C8E0D63",
    x"1C8DD5F0",
    x"1C8D9E94",
    x"1C8D674C",
    x"1C8D301B",
    x"1C8CF8FF",
    x"1C8CC1F8",
    x"1C8C8B07",
    x"1C8C542C",
    x"1C8C1D65",
    x"1C8BE6B5",
    x"1C8BB019",
    x"1C8B7993",
    x"1C8B4322",
    x"1C8B0CC7",
    x"1C8AD680",
    x"1C8AA04F",
    x"1C8A6A33",
    x"1C8A342C",
    x"1C89FE3A",
    x"1C89C85D",
    x"1C899296",
    x"1C895CE3",
    x"1C892745",
    x"1C88F1BC",
    x"1C88BC48",
    x"1C8886E9",
    x"1C88519F",
    x"1C881C69",
    x"1C87E749",
    x"1C87B23D",
    x"1C877D45",
    x"1C874863",
    x"1C871395",
    x"1C86DEDB",
    x"1C86AA37",
    x"1C8675A6",
    x"1C86412B",
    x"1C860CC4",
    x"1C85D871",
    x"1C85A432",
    x"1C857008",
    x"1C853BF3",
    x"1C8507F2",
    x"1C84D405",
    x"1C84A02C",
    x"1C846C68",
    x"1C8438B7",
    x"1C84051B",
    x"1C83D193",
    x"1C839E1F",
    x"1C836AC0",
    x"1C833774",
    x"1C83043C",
    x"1C82D119",
    x"1C829E09",
    x"1C826B0D",
    x"1C823825",
    x"1C820551",
    x"1C81D291",
    x"1C819FE5",
    x"1C816D4C",
    x"1C813AC7",
    x"1C810856",
    x"1C80D5F9",
    x"1C80A3AF",
    x"1C807179",
    x"1C803F57",
    x"1C800D48",
    x"1C7FB698",
    x"1C7F52C8",
    x"1C7EEF20",
    x"1C7E8B9E",
    x"1C7E2843",
    x"1C7DC50E",
    x"1C7D6201",
    x"1C7CFF1A",
    x"1C7C9C59",
    x"1C7C39BF",
    x"1C7BD74C",
    x"1C7B74FF",
    x"1C7B12D9",
    x"1C7AB0D8",
    x"1C7A4EFE",
    x"1C79ED4B",
    x"1C798BBD",
    x"1C792A56",
    x"1C78C914",
    x"1C7867F8",
    x"1C780703",
    x"1C77A633",
    x"1C774589",
    x"1C76E505",
    x"1C7684A6",
    x"1C76246D",
    x"1C75C459",
    x"1C75646C",
    x"1C7504A3",
    x"1C74A500",
    x"1C744582",
    x"1C73E62A",
    x"1C7386F6",
    x"1C7327E8",
    x"1C72C8FF",
    x"1C726A3B",
    x"1C720B9C",
    x"1C71AD22",
    x"1C714ECD",
    x"1C70F09C",
    x"1C709291",
    x"1C7034AA",
    x"1C6FD6E8",
    x"1C6F794A",
    x"1C6F1BD1",
    x"1C6EBE7C",
    x"1C6E614C",
    x"1C6E0440",
    x"1C6DA759",
    x"1C6D4A95",
    x"1C6CEDF6",
    x"1C6C917B",
    x"1C6C3525",
    x"1C6BD8F2",
    x"1C6B7CE3",
    x"1C6B20F8",
    x"1C6AC531",
    x"1C6A698E",
    x"1C6A0E0F",
    x"1C69B2B3",
    x"1C69577B",
    x"1C68FC67",
    x"1C68A176",
    x"1C6846A9",
    x"1C67EBFF",
    x"1C679178",
    x"1C673715",
    x"1C66DCD5",
    x"1C6682B9",
    x"1C6628BF",
    x"1C65CEE9",
    x"1C657535",
    x"1C651BA5",
    x"1C64C238",
    x"1C6468ED",
    x"1C640FC6",
    x"1C63B6C1",
    x"1C635DDF",
    x"1C630520",
    x"1C62AC83",
    x"1C625409",
    x"1C61FBB1",
    x"1C61A37C",
    x"1C614B6A",
    x"1C60F379",
    x"1C609BAB",
    x"1C604400",
    x"1C5FEC76",
    x"1C5F950F",
    x"1C5F3DCA",
    x"1C5EE6A7",
    x"1C5E8FA6",
    x"1C5E38C6",
    x"1C5DE209",
    x"1C5D8B6E",
    x"1C5D34F4",
    x"1C5CDE9C",
    x"1C5C8866",
    x"1C5C3252",
    x"1C5BDC5F",
    x"1C5B868E",
    x"1C5B30DE",
    x"1C5ADB50",
    x"1C5A85E3",
    x"1C5A3097",
    x"1C59DB6D",
    x"1C598663",
    x"1C59317C",
    x"1C58DCB5",
    x"1C58880F",
    x"1C58338A",
    x"1C57DF27",
    x"1C578AE4",
    x"1C5736C2",
    x"1C56E2C1",
    x"1C568EE1",
    x"1C563B22",
    x"1C55E783",
    x"1C559405",
    x"1C5540A7",
    x"1C54ED6A",
    x"1C549A4E",
    x"1C544752",
    x"1C53F476",
    x"1C53A1BB",
    x"1C534F20",
    x"1C52FCA5",
    x"1C52AA4A",
    x"1C525810",
    x"1C5205F5",
    x"1C51B3FB",
    x"1C516221",
    x"1C511066",
    x"1C50BECC",
    x"1C506D51",
    x"1C501BF7",
    x"1C4FCABC",
    x"1C4F79A0",
    x"1C4F28A4",
    x"1C4ED7C8",
    x"1C4E870C",
    x"1C4E366F",
    x"1C4DE5F1",
    x"1C4D9593",
    x"1C4D4554",
    x"1C4CF535",
    x"1C4CA535",
    x"1C4C5554",
    x"1C4C0592",
    x"1C4BB5F0",
    x"1C4B666C",
    x"1C4B1708",
    x"1C4AC7C2",
    x"1C4A789B",
    x"1C4A2994",
    x"1C49DAAB",
    x"1C498BE1",
    x"1C493D36",
    x"1C48EEA9",
    x"1C48A03B",
    x"1C4851EC",
    x"1C4803BB",
    x"1C47B5A9",
    x"1C4767B5",
    x"1C4719E0",
    x"1C46CC29",
    x"1C467E90",
    x"1C463116",
    x"1C45E3BA",
    x"1C45967C",
    x"1C45495C",
    x"1C44FC5B",
    x"1C44AF77",
    x"1C4462B2",
    x"1C44160A",
    x"1C43C981",
    x"1C437D15",
    x"1C4330C7",
    x"1C42E497",
    x"1C429884",
    x"1C424C8F",
    x"1C4200B8",
    x"1C41B4FF",
    x"1C416963",
    x"1C411DE5",
    x"1C40D284",
    x"1C408740",
    x"1C403C1A",
    x"1C3FF111",
    x"1C3FA626",
    x"1C3F5B57",
    x"1C3F10A6",
    x"1C3EC612",
    x"1C3E7B9B",
    x"1C3E3142",
    x"1C3DE705",
    x"1C3D9CE5",
    x"1C3D52E2",
    x"1C3D08FC",
    x"1C3CBF33",
    x"1C3C7587",
    x"1C3C2BF7",
    x"1C3BE285",
    x"1C3B992F",
    x"1C3B4FF5",
    x"1C3B06D8",
    x"1C3ABDD8",
    x"1C3A74F4",
    x"1C3A2C2C",
    x"1C39E381",
    x"1C399AF2",
    x"1C395280",
    x"1C390A2A",
    x"1C38C1F0",
    x"1C3879D2",
    x"1C3831D1",
    x"1C37E9EC",
    x"1C37A222",
    x"1C375A75",
    x"1C3712E4",
    x"1C36CB6E",
    x"1C368415",
    x"1C363CD7",
    x"1C35F5B5",
    x"1C35AEAF",
    x"1C3567C5",
    x"1C3520F6",
    x"1C34DA43",
    x"1C3493AB",
    x"1C344D2F",
    x"1C3406CF",
    x"1C33C08A",
    x"1C337A61",
    x"1C333452",
    x"1C32EE60",
    x"1C32A888",
    x"1C3262CC",
    x"1C321D2B",
    x"1C31D7A5",
    x"1C31923B",
    x"1C314CEB",
    x"1C3107B6",
    x"1C30C29D",
    x"1C307D9E",
    x"1C3038BB",
    x"1C2FF3F2",
    x"1C2FAF44",
    x"1C2F6AB1",
    x"1C2F2639",
    x"1C2EE1DB",
    x"1C2E9D98",
    x"1C2E5970",
    x"1C2E1562",
    x"1C2DD16F",
    x"1C2D8D97",
    x"1C2D49D9",
    x"1C2D0635",
    x"1C2CC2AC",
    x"1C2C7F3D",
    x"1C2C3BE8",
    x"1C2BF8AE",
    x"1C2BB58E",
    x"1C2B7288",
    x"1C2B2F9D",
    x"1C2AECCB",
    x"1C2AAA14",
    x"1C2A6776",
    x"1C2A24F3",
    x"1C29E289",
    x"1C29A03A",
    x"1C295E04",
    x"1C291BE8",
    x"1C28D9E6",
    x"1C2897FE",
    x"1C285630",
    x"1C28147B",
    x"1C27D2E0",
    x"1C27915E",
    x"1C274FF6",
    x"1C270EA8",
    x"1C26CD73",
    x"1C268C57",
    x"1C264B55",
    x"1C260A6C",
    x"1C25C99D",
    x"1C2588E7",
    x"1C25484A",
    x"1C2507C6",
    x"1C24C75C",
    x"1C24870A",
    x"1C2446D2",
    x"1C2406B3",
    x"1C23C6AD",
    x"1C2386C0",
    x"1C2346EC",
    x"1C230730",
    x"1C22C78E",
    x"1C228804",
    x"1C224894",
    x"1C22093C",
    x"1C21C9FC",
    x"1C218AD6",
    x"1C214BC8",
    x"1C210CD3",
    x"1C20CDF6",
    x"1C208F32",
    x"1C205086",
    x"1C2011F3",
    x"1C1FD378",
    x"1C1F9516",
    x"1C1F56CC",
    x"1C1F189A",
    x"1C1EDA80",
    x"1C1E9C7F",
    x"1C1E5E96",
    x"1C1E20C5",
    x"1C1DE30C",
    x"1C1DA56C",
    x"1C1D67E3",
    x"1C1D2A73",
    x"1C1CED1A",
    x"1C1CAFD9",
    x"1C1C72B1",
    x"1C1C35A0",
    x"1C1BF8A7",
    x"1C1BBBC5",
    x"1C1B7EFC",
    x"1C1B424A",
    x"1C1B05B0",
    x"1C1AC92E",
    x"1C1A8CC3",
    x"1C1A5070",
    x"1C1A1434",
    x"1C19D810",
    x"1C199C03",
    x"1C19600E",
    x"1C192430",
    x"1C18E86A",
    x"1C18ACBB",
    x"1C187123",
    x"1C1835A2",
    x"1C17FA39",
    x"1C17BEE7",
    x"1C1783AC",
    x"1C174888",
    x"1C170D7B",
    x"1C16D285",
    x"1C1697A7",
    x"1C165CDF",
    x"1C16222E",
    x"1C15E794",
    x"1C15AD11",
    x"1C1572A5",
    x"1C153850",
    x"1C14FE11",
    x"1C14C3E9",
    x"1C1489D8",
    x"1C144FDD",
    x"1C1415FA",
    x"1C13DC2C",
    x"1C13A275",
    x"1C1368D5",
    x"1C132F4C",
    x"1C12F5D8",
    x"1C12BC7B",
    x"1C128335",
    x"1C124A05",
    x"1C1210EB",
    x"1C11D7E8",
    x"1C119EFB",
    x"1C116624",
    x"1C112D63",
    x"1C10F4B8",
    x"1C10BC24",
    x"1C1083A5",
    x"1C104B3D",
    x"1C1012EA",
    x"1C0FDAAE",
    x"1C0FA287",
    x"1C0F6A77",
    x"1C0F327C",
    x"1C0EFA97",
    x"1C0EC2C8",
    x"1C0E8B0F",
    x"1C0E536C",
    x"1C0E1BDE",
    x"1C0DE466",
    x"1C0DAD04",
    x"1C0D75B7",
    x"1C0D3E80",
    x"1C0D075E",
    x"1C0CD052",
    x"1C0C995B",
    x"1C0C627A",
    x"1C0C2BAE",
    x"1C0BF4F8",
    x"1C0BBE57",
    x"1C0B87CB",
    x"1C0B5155",
    x"1C0B1AF4",
    x"1C0AE4A8",
    x"1C0AAE71",
    x"1C0A784F",
    x"1C0A4243",
    x"1C0A0C4C",
    x"1C09D669",
    x"1C09A09C",
    x"1C096AE4",
    x"1C093541",
    x"1C08FFB2",
    x"1C08CA39",
    x"1C0894D4",
    x"1C085F85",
    x"1C082A4A",
    x"1C07F524",
    x"1C07C012",
    x"1C078B15",
    x"1C07562D",
    x"1C07215A",
    x"1C06EC9B",
    x"1C06B7F1",
    x"1C06835C",
    x"1C064EDB",
    x"1C061A6E",
    x"1C05E616",
    x"1C05B1D2",
    x"1C057DA3",
    x"1C054988",
    x"1C051582",
    x"1C04E18F",
    x"1C04ADB1",
    x"1C0479E8",
    x"1C044632",
    x"1C041291",
    x"1C03DF04",
    x"1C03AB8B",
    x"1C037826",
    x"1C0344D5",
    x"1C031198",
    x"1C02DE6F",
    x"1C02AB5A",
    x"1C027859",
    x"1C02456C",
    x"1C021293",
    x"1C01DFCD",
    x"1C01AD1C",
    x"1C017A7E",
    x"1C0147F4",
    x"1C01157E",
    x"1C00E31B",
    x"1C00B0CD",
    x"1C007E91",
    x"1C004C6A",
    x"1C001A56",
    x"1BFFD0AA",
    x"1BFF6CD0",
    x"1BFF091D",
    x"1BFEA591",
    x"1BFE422C",
    x"1BFDDEED",
    x"1BFD7BD6",
    x"1BFD18E4",
    x"1BFCB61A",
    x"1BFC5376",
    x"1BFBF0F9",
    x"1BFB8EA2",
    x"1BFB2C71",
    x"1BFACA67",
    x"1BFA6883",
    x"1BFA06C6",
    x"1BF9A52E",
    x"1BF943BC",
    x"1BF8E271",
    x"1BF8814C",
    x"1BF8204C",
    x"1BF7BF72",
    x"1BF75EBE",
    x"1BF6FE30",
    x"1BF69DC8",
    x"1BF63D85",
    x"1BF5DD68",
    x"1BF57D70",
    x"1BF51D9E",
    x"1BF4BDF1",
    x"1BF45E69",
    x"1BF3FF07",
    x"1BF39FCA",
    x"1BF340B2",
    x"1BF2E1BF",
    x"1BF282F2",
    x"1BF22449",
    x"1BF1C5C5",
    x"1BF16767",
    x"1BF1092D",
    x"1BF0AB17",
    x"1BF04D27",
    x"1BEFEF5B",
    x"1BEF91B4",
    x"1BEF3431",
    x"1BEED6D3",
    x"1BEE7999",
    x"1BEE1C84",
    x"1BEDBF93",
    x"1BED62C6",
    x"1BED061E",
    x"1BECA99A",
    x"1BEC4D39",
    x"1BEBF0FD",
    x"1BEB94E5",
    x"1BEB38F1",
    x"1BEADD21",
    x"1BEA8174",
    x"1BEA25EB",
    x"1BE9CA87",
    x"1BE96F45",
    x"1BE91428",
    x"1BE8B92D",
    x"1BE85E57",
    x"1BE803A4",
    x"1BE7A914",
    x"1BE74EA8",
    x"1BE6F45F",
    x"1BE69A39",
    x"1BE64036",
    x"1BE5E657",
    x"1BE58C9A",
    x"1BE53301",
    x"1BE4D98A",
    x"1BE48037",
    x"1BE42706",
    x"1BE3CDF8",
    x"1BE3750D",
    x"1BE31C45",
    x"1BE2C39F",
    x"1BE26B1C",
    x"1BE212BB",
    x"1BE1BA7D",
    x"1BE16262",
    x"1BE10A68",
    x"1BE0B291",
    x"1BE05ADD",
    x"1BE0034A",
    x"1BDFABDA",
    x"1BDF548C",
    x"1BDEFD60",
    x"1BDEA656",
    x"1BDE4F6E",
    x"1BDDF8A8",
    x"1BDDA204",
    x"1BDD4B82",
    x"1BDCF521",
    x"1BDC9EE2",
    x"1BDC48C5",
    x"1BDBF2C9",
    x"1BDB9CEF",
    x"1BDB4737",
    x"1BDAF19F",
    x"1BDA9C2A",
    x"1BDA46D5",
    x"1BD9F1A2",
    x"1BD99C91",
    x"1BD947A0",
    x"1BD8F2D1",
    x"1BD89E22",
    x"1BD84995",
    x"1BD7F529",
    x"1BD7A0DE",
    x"1BD74CB3",
    x"1BD6F8AA",
    x"1BD6A4C1",
    x"1BD650F9",
    x"1BD5FD52",
    x"1BD5A9CB",
    x"1BD55665",
    x"1BD5031F",
    x"1BD4AFFA",
    x"1BD45CF6",
    x"1BD40A12",
    x"1BD3B74E",
    x"1BD364AB",
    x"1BD31227",
    x"1BD2BFC4",
    x"1BD26D82",
    x"1BD21B5F",
    x"1BD1C95C",
    x"1BD17779",
    x"1BD125B7",
    x"1BD0D414",
    x"1BD08291",
    x"1BD0312E",
    x"1BCFDFEB",
    x"1BCF8EC7",
    x"1BCF3DC3",
    x"1BCEECDF",
    x"1BCE9C1A",
    x"1BCE4B75",
    x"1BCDFAEF",
    x"1BCDAA89",
    x"1BCD5A42",
    x"1BCD0A1A",
    x"1BCCBA12",
    x"1BCC6A29",
    x"1BCC1A5F",
    x"1BCBCAB4",
    x"1BCB7B29",
    x"1BCB2BBC",
    x"1BCADC6E",
    x"1BCA8D40",
    x"1BCA3E30",
    x"1BC9EF3F",
    x"1BC9A06D",
    x"1BC951BA",
    x"1BC90325",
    x"1BC8B4AF",
    x"1BC86658",
    x"1BC8181F",
    x"1BC7CA05",
    x"1BC77C0A",
    x"1BC72E2C",
    x"1BC6E06D",
    x"1BC692CD",
    x"1BC6454B",
    x"1BC5F7E7",
    x"1BC5AAA1",
    x"1BC55D79",
    x"1BC51070",
    x"1BC4C385",
    x"1BC476B7",
    x"1BC42A08",
    x"1BC3DD76",
    x"1BC39103",
    x"1BC344AD",
    x"1BC2F875",
    x"1BC2AC5B",
    x"1BC2605E",
    x"1BC21480",
    x"1BC1C8BE",
    x"1BC17D1B",
    x"1BC13195",
    x"1BC0E62C",
    x"1BC09AE1",
    x"1BC04FB3",
    x"1BC004A3",
    x"1BBFB9AF",
    x"1BBF6ED9",
    x"1BBF2421",
    x"1BBED985",
    x"1BBE8F07",
    x"1BBE44A5",
    x"1BBDFA61",
    x"1BBDB03A",
    x"1BBD662F",
    x"1BBD1C42",
    x"1BBCD271",
    x"1BBC88BE",
    x"1BBC3F27",
    x"1BBBF5AC",
    x"1BBBAC4F",
    x"1BBB630E",
    x"1BBB19E9",
    x"1BBAD0E1",
    x"1BBA87F6",
    x"1BBA3F27",
    x"1BB9F675",
    x"1BB9ADDF",
    x"1BB96565",
    x"1BB91D07",
    x"1BB8D4C6",
    x"1BB88CA1",
    x"1BB84498",
    x"1BB7FCAB",
    x"1BB7B4DB",
    x"1BB76D26",
    x"1BB7258E",
    x"1BB6DE11",
    x"1BB696B0",
    x"1BB64F6B",
    x"1BB60842",
    x"1BB5C135",
    x"1BB57A43",
    x"1BB5336D",
    x"1BB4ECB3",
    x"1BB4A614",
    x"1BB45F91",
    x"1BB41929",
    x"1BB3D2DD",
    x"1BB38CAD",
    x"1BB34697",
    x"1BB3009E",
    x"1BB2BABF",
    x"1BB274FC",
    x"1BB22F54",
    x"1BB1E9C7",
    x"1BB1A455",
    x"1BB15EFE",
    x"1BB119C3",
    x"1BB0D4A2",
    x"1BB08F9D",
    x"1BB04AB2",
    x"1BB005E2",
    x"1BAFC12D",
    x"1BAF7C93",
    x"1BAF3814",
    x"1BAEF3AF",
    x"1BAEAF66",
    x"1BAE6B36",
    x"1BAE2722",
    x"1BADE328",
    x"1BAD9F48",
    x"1BAD5B83",
    x"1BAD17D9",
    x"1BACD449",
    x"1BAC90D3",
    x"1BAC4D78",
    x"1BAC0A36",
    x"1BABC710",
    x"1BAB8403",
    x"1BAB4110",
    x"1BAAFE38",
    x"1BAABB7A",
    x"1BAA78D6",
    x"1BAA364B",
    x"1BA9F3DB",
    x"1BA9B185",
    x"1BA96F48",
    x"1BA92D26",
    x"1BA8EB1D",
    x"1BA8A92E",
    x"1BA86759",
    x"1BA8259D",
    x"1BA7E3FC",
    x"1BA7A273",
    x"1BA76105",
    x"1BA71FB0",
    x"1BA6DE74",
    x"1BA69D52",
    x"1BA65C49",
    x"1BA61B5A",
    x"1BA5DA84",
    x"1BA599C7",
    x"1BA55923",
    x"1BA51899",
    x"1BA4D828",
    x"1BA497D0",
    x"1BA45792",
    x"1BA4176C",
    x"1BA3D75F",
    x"1BA3976C",
    x"1BA35791",
    x"1BA317CF",
    x"1BA2D826",
    x"1BA29896",
    x"1BA2591F",
    x"1BA219C1",
    x"1BA1DA7B",
    x"1BA19B4E",
    x"1BA15C3A",
    x"1BA11D3E",
    x"1BA0DE5B",
    x"1BA09F90",
    x"1BA060DE",
    x"1BA02245",
    x"1B9FE3C3",
    x"1B9FA55B",
    x"1B9F670A",
    x"1B9F28D2",
    x"1B9EEAB2",
    x"1B9EACAB",
    x"1B9E6EBB",
    x"1B9E30E4",
    x"1B9DF325",
    x"1B9DB57E",
    x"1B9D77EF",
    x"1B9D3A78",
    x"1B9CFD1A",
    x"1B9CBFD3",
    x"1B9C82A4",
    x"1B9C458D",
    x"1B9C088D",
    x"1B9BCBA6",
    x"1B9B8ED6",
    x"1B9B521E",
    x"1B9B157E",
    x"1B9AD8F6",
    x"1B9A9C85",
    x"1B9A602B",
    x"1B9A23E9",
    x"1B99E7BF",
    x"1B99ABAC",
    x"1B996FB1",
    x"1B9933CD",
    x"1B98F801",
    x"1B98BC4B",
    x"1B9880AD",
    x"1B984527",
    x"1B9809B7",
    x"1B97CE5F",
    x"1B97931E",
    x"1B9757F4",
    x"1B971CE1",
    x"1B96E1E6",
    x"1B96A701",
    x"1B966C33",
    x"1B96317C",
    x"1B95F6DD",
    x"1B95BC54",
    x"1B9581E1",
    x"1B954786",
    x"1B950D42",
    x"1B94D314",
    x"1B9498FD",
    x"1B945EFC",
    x"1B942512",
    x"1B93EB3F",
    x"1B93B183",
    x"1B9377DD",
    x"1B933E4D",
    x"1B9304D4",
    x"1B92CB71",
    x"1B929225",
    x"1B9258EF",
    x"1B921FCF",
    x"1B91E6C6",
    x"1B91ADD3",
    x"1B9174F6",
    x"1B913C30",
    x"1B91037F",
    x"1B90CAE5",
    x"1B909261",
    x"1B9059F3",
    x"1B90219A",
    x"1B8FE958",
    x"1B8FB12C",
    x"1B8F7916",
    x"1B8F4116",
    x"1B8F092B",
    x"1B8ED156",
    x"1B8E9997",
    x"1B8E61EE",
    x"1B8E2A5B",
    x"1B8DF2DD",
    x"1B8DBB75",
    x"1B8D8423",
    x"1B8D4CE6",
    x"1B8D15BF",
    x"1B8CDEAD",
    x"1B8CA7B1",
    x"1B8C70CA",
    x"1B8C39F9",
    x"1B8C033D",
    x"1B8BCC96",
    x"1B8B9605",
    x"1B8B5F89",
    x"1B8B2922",
    x"1B8AF2D1",
    x"1B8ABC94",
    x"1B8A866D",
    x"1B8A505B",
    x"1B8A1A5F",
    x"1B89E477",
    x"1B89AEA4",
    x"1B8978E6",
    x"1B89433E",
    x"1B890DAA",
    x"1B88D82B",
    x"1B88A2C1",
    x"1B886D6C",
    x"1B88382B",
    x"1B880300",
    x"1B87CDE9",
    x"1B8798E7",
    x"1B8763FA",
    x"1B872F21",
    x"1B86FA5D",
    x"1B86C5AD",
    x"1B869112",
    x"1B865C8C",
    x"1B86281A",
    x"1B85F3BD",
    x"1B85BF74",
    x"1B858B3F",
    x"1B85571F",
    x"1B852313",
    x"1B84EF1B",
    x"1B84BB38",
    x"1B848769",
    x"1B8453AE",
    x"1B842008",
    x"1B83EC75",
    x"1B83B8F7",
    x"1B83858D",
    x"1B835237",
    x"1B831EF5",
    x"1B82EBC6",
    x"1B82B8AC",
    x"1B8285A6",
    x"1B8252B4",
    x"1B821FD6",
    x"1B81ED0B",
    x"1B81BA54",
    x"1B8187B1",
    x"1B815522",
    x"1B8122A7",
    x"1B80F03F",
    x"1B80BDEB",
    x"1B808BAB",
    x"1B80597E",
    x"1B802765",
    x"1B7FEABF",
    x"1B7F86DA",
    x"1B7F231D",
    x"1B7EBF87",
    x"1B7E5C18",
    x"1B7DF8CF",
    x"1B7D95AD",
    x"1B7D32B2",
    x"1B7CCFDE",
    x"1B7C6D30",
    x"1B7C0AA8",
    x"1B7BA847",
    x"1B7B460D",
    x"1B7AE3F9",
    x"1B7A820B",
    x"1B7A2043",
    x"1B79BEA1",
    x"1B795D26",
    x"1B78FBD1",
    x"1B789AA1",
    x"1B783998",
    x"1B77D8B4",
    x"1B7777F6",
    x"1B77175E",
    x"1B76B6EC",
    x"1B7656A0",
    x"1B75F678",
    x"1B759677",
    x"1B75369B",
    x"1B74D6E4",
    x"1B747753",
    x"1B7417E7",
    x"1B73B8A0",
    x"1B73597F",
    x"1B72FA82",
    x"1B729BAB",
    x"1B723CF9",
    x"1B71DE6B",
    x"1B718003",
    x"1B7121BF",
    x"1B70C3A1",
    x"1B7065A7",
    x"1B7007D1",
    x"1B6FAA20",
    x"1B6F4C94",
    x"1B6EEF2D",
    x"1B6E91E9",
    x"1B6E34CB",
    x"1B6DD7D0",
    x"1B6D7AFA",
    x"1B6D1E48",
    x"1B6CC1BA",
    x"1B6C6551",
    x"1B6C090B",
    x"1B6BACEA",
    x"1B6B50EC",
    x"1B6AF512",
    x"1B6A995C",
    x"1B6A3DCA",
    x"1B69E25C",
    x"1B698712",
    x"1B692BEB",
    x"1B68D0E7",
    x"1B687607",
    x"1B681B4B",
    x"1B67C0B2",
    x"1B67663C",
    x"1B670BEA",
    x"1B66B1BB",
    x"1B6657AF",
    x"1B65FDC7",
    x"1B65A401",
    x"1B654A5E",
    x"1B64F0DF",
    x"1B649782",
    x"1B643E49",
    x"1B63E532",
    x"1B638C3D",
    x"1B63336C",
    x"1B62DABD",
    x"1B628231",
    x"1B6229C8",
    x"1B61D180",
    x"1B61795C",
    x"1B61215A",
    x"1B60C97A",
    x"1B6071BC",
    x"1B601A21",
    x"1B5FC2A8",
    x"1B5F6B51",
    x"1B5F141C",
    x"1B5EBD09",
    x"1B5E6618",
    x"1B5E0F49",
    x"1B5DB89C",
    x"1B5D6211",
    x"1B5D0BA8",
    x"1B5CB560",
    x"1B5C5F3A",
    x"1B5C0936",
    x"1B5BB353",
    x"1B5B5D91",
    x"1B5B07F2",
    x"1B5AB273",
    x"1B5A5D16",
    x"1B5A07DA",
    x"1B59B2C0",
    x"1B595DC7",
    x"1B5908EF",
    x"1B58B438",
    x"1B585FA2",
    x"1B580B2D",
    x"1B57B6D9",
    x"1B5762A6",
    x"1B570E94",
    x"1B56BAA3",
    x"1B5666D2",
    x"1B561322",
    x"1B55BF93",
    x"1B556C25",
    x"1B5518D7",
    x"1B54C5A9",
    x"1B54729C",
    x"1B541FB0",
    x"1B53CCE4",
    x"1B537A38",
    x"1B5327AC",
    x"1B52D541",
    x"1B5282F5",
    x"1B5230CA",
    x"1B51DEBF",
    x"1B518CD4",
    x"1B513B09",
    x"1B50E95E",
    x"1B5097D3",
    x"1B504668",
    x"1B4FF51C",
    x"1B4FA3F0",
    x"1B4F52E4",
    x"1B4F01F7",
    x"1B4EB12A",
    x"1B4E607D",
    x"1B4E0FEF",
    x"1B4DBF80",
    x"1B4D6F31",
    x"1B4D1F01",
    x"1B4CCEF1",
    x"1B4C7F00",
    x"1B4C2F2E",
    x"1B4BDF7B",
    x"1B4B8FE7",
    x"1B4B4072",
    x"1B4AF11D",
    x"1B4AA1E6",
    x"1B4A52CE",
    x"1B4A03D5",
    x"1B49B4FB",
    x"1B496640",
    x"1B4917A3",
    x"1B48C926",
    x"1B487AC6",
    x"1B482C86",
    x"1B47DE63",
    x"1B479060",
    x"1B47427B",
    x"1B46F4B4",
    x"1B46A70B",
    x"1B465981",
    x"1B460C16",
    x"1B45BEC8",
    x"1B457198",
    x"1B452487",
    x"1B44D794",
    x"1B448ABF",
    x"1B443E07",
    x"1B43F16E",
    x"1B43A4F3",
    x"1B435895",
    x"1B430C56",
    x"1B42C034",
    x"1B42742F",
    x"1B422849",
    x"1B41DC80",
    x"1B4190D5",
    x"1B414547",
    x"1B40F9D6",
    x"1B40AE84",
    x"1B40634E",
    x"1B401836",
    x"1B3FCD3B",
    x"1B3F825E",
    x"1B3F379D",
    x"1B3EECFA",
    x"1B3EA274",
    x"1B3E580B",
    x"1B3E0DBF",
    x"1B3DC390",
    x"1B3D797F",
    x"1B3D2F8A",
    x"1B3CE5B1",
    x"1B3C9BF6",
    x"1B3C5258",
    x"1B3C08D6",
    x"1B3BBF71",
    x"1B3B7628",
    x"1B3B2CFC",
    x"1B3AE3ED",
    x"1B3A9AFA",
    x"1B3A5224",
    x"1B3A096A",
    x"1B39C0CD",
    x"1B39784B",
    x"1B392FE7",
    x"1B38E79E",
    x"1B389F72",
    x"1B385761",
    x"1B380F6D",
    x"1B37C795",
    x"1B377FD9",
    x"1B373839",
    x"1B36F0B5",
    x"1B36A94D",
    x"1B366201",
    x"1B361AD1",
    x"1B35D3BC",
    x"1B358CC3",
    x"1B3545E6",
    x"1B34FF25",
    x"1B34B87F",
    x"1B3471F5",
    x"1B342B86",
    x"1B33E533",
    x"1B339EFB",
    x"1B3358DE",
    x"1B3312DD",
    x"1B32CCF8",
    x"1B32872D",
    x"1B32417E",
    x"1B31FBEA",
    x"1B31B671",
    x"1B317113",
    x"1B312BD1",
    x"1B30E6A9",
    x"1B30A19D",
    x"1B305CAB",
    x"1B3017D4",
    x"1B2FD318",
    x"1B2F8E77",
    x"1B2F49F1",
    x"1B2F0585",
    x"1B2EC135",
    x"1B2E7CFF",
    x"1B2E38E3",
    x"1B2DF4E2",
    x"1B2DB0FC",
    x"1B2D6D30",
    x"1B2D297E",
    x"1B2CE5E7",
    x"1B2CA26B",
    x"1B2C5F08",
    x"1B2C1BC0",
    x"1B2BD893",
    x"1B2B957F",
    x"1B2B5286",
    x"1B2B0FA7",
    x"1B2ACCE2",
    x"1B2A8A37",
    x"1B2A47A6",
    x"1B2A052F",
    x"1B29C2D2",
    x"1B29808E",
    x"1B293E65",
    x"1B28FC56",
    x"1B28BA60",
    x"1B287884",
    x"1B2836C2",
    x"1B27F519",
    x"1B27B38A",
    x"1B277215",
    x"1B2730B9",
    x"1B26EF77",
    x"1B26AE4E",
    x"1B266D3F",
    x"1B262C49",
    x"1B25EB6C",
    x"1B25AAA9",
    x"1B2569FF",
    x"1B25296E",
    x"1B24E8F6",
    x"1B24A898",
    x"1B246853",
    x"1B242826",
    x"1B23E813",
    x"1B23A819",
    x"1B236838",
    x"1B232870",
    x"1B22E8C0",
    x"1B22A92A",
    x"1B2269AC",
    x"1B222A47",
    x"1B21EAFB",
    x"1B21ABC8",
    x"1B216CAD",
    x"1B212DAB",
    x"1B20EEC1",
    x"1B20AFF0",
    x"1B207138",
    x"1B203298",
    x"1B1FF410",
    x"1B1FB5A1",
    x"1B1F774A",
    x"1B1F390C",
    x"1B1EFAE6",
    x"1B1EBCD8",
    x"1B1E7EE2",
    x"1B1E4105",
    x"1B1E033F",
    x"1B1DC592",
    x"1B1D87FD",
    x"1B1D4A80",
    x"1B1D0D1B",
    x"1B1CCFCE",
    x"1B1C9298",
    x"1B1C557B",
    x"1B1C1876",
    x"1B1BDB88",
    x"1B1B9EB2",
    x"1B1B61F4",
    x"1B1B254E",
    x"1B1AE8BF",
    x"1B1AAC48",
    x"1B1A6FE8",
    x"1B1A33A0",
    x"1B19F770",
    x"1B19BB57",
    x"1B197F56",
    x"1B19436C",
    x"1B190799",
    x"1B18CBDE",
    x"1B18903A",
    x"1B1854AD",
    x"1B181937",
    x"1B17DDD9",
    x"1B17A292",
    x"1B176762",
    x"1B172C49",
    x"1B16F148",
    x"1B16B65D",
    x"1B167B89",
    x"1B1640CC",
    x"1B160626",
    x"1B15CB97",
    x"1B15911F",
    x"1B1556BE",
    x"1B151C74",
    x"1B14E240",
    x"1B14A823",
    x"1B146E1C",
    x"1B14342D",
    x"1B13FA54",
    x"1B13C091",
    x"1B1386E5",
    x"1B134D50",
    x"1B1313D1",
    x"1B12DA68",
    x"1B12A116",
    x"1B1267DA",
    x"1B122EB5",
    x"1B11F5A6",
    x"1B11BCAD",
    x"1B1183CB",
    x"1B114AFE",
    x"1B111248",
    x"1B10D9A8",
    x"1B10A11E",
    x"1B1068AA",
    x"1B10304C",
    x"1B0FF804",
    x"1B0FBFD2",
    x"1B0F87B6",
    x"1B0F4FB0",
    x"1B0F17C0",
    x"1B0EDFE6",
    x"1B0EA821",
    x"1B0E7072",
    x"1B0E38D9",
    x"1B0E0156",
    x"1B0DC9E8",
    x"1B0D9290",
    x"1B0D5B4E",
    x"1B0D2421",
    x"1B0CED09",
    x"1B0CB608",
    x"1B0C7F1B",
    x"1B0C4844",
    x"1B0C1183",
    x"1B0BDAD7",
    x"1B0BA440",
    x"1B0B6DBE",
    x"1B0B3752",
    x"1B0B00FB",
    x"1B0ACAB9",
    x"1B0A948D",
    x"1B0A5E75",
    x"1B0A2873",
    x"1B09F286",
    x"1B09BCAD",
    x"1B0986EA",
    x"1B09513C",
    x"1B091BA3",
    x"1B08E61E",
    x"1B08B0AF",
    x"1B087B54",
    x"1B08460F",
    x"1B0810DE",
    x"1B07DBC1",
    x"1B07A6BA",
    x"1B0771C7",
    x"1B073CE9",
    x"1B070820",
    x"1B06D36B",
    x"1B069ECA",
    x"1B066A3F",
    x"1B0635C7",
    x"1B060165",
    x"1B05CD16",
    x"1B0598DC",
    x"1B0564B7",
    x"1B0530A6",
    x"1B04FCA9",
    x"1B04C8C0",
    x"1B0494EC",
    x"1B04612C",
    x"1B042D80",
    x"1B03F9E8",
    x"1B03C665",
    x"1B0392F5",
    x"1B035F9A",
    x"1B032C53",
    x"1B02F91F",
    x"1B02C600",
    x"1B0292F5",
    x"1B025FFD",
    x"1B022D1A",
    x"1B01FA4A",
    x"1B01C78E",
    x"1B0194E6",
    x"1B016252",
    x"1B012FD1",
    x"1B00FD64",
    x"1B00CB0B",
    x"1B0098C6",
    x"1B006694",
    x"1B003476",
    x"1B00026B",
    x"1AFFA0E7",
    x"1AFF3D20",
    x"1AFED980",
    x"1AFE7606",
    x"1AFE12B3",
    x"1AFDAF87",
    x"1AFD4C82",
    x"1AFCE9A4",
    x"1AFC86EC",
    x"1AFC245A",
    x"1AFBC1EF",
    x"1AFB5FAB",
    x"1AFAFD8C",
    x"1AFA9B95",
    x"1AFA39C3",
    x"1AF9D817",
    x"1AF97692",
    x"1AF91533",
    x"1AF8B3F9",
    x"1AF852E6",
    x"1AF7F1F9",
    x"1AF79131",
    x"1AF7308F",
    x"1AF6D013",
    x"1AF66FBD",
    x"1AF60F8C",
    x"1AF5AF81",
    x"1AF54F9B",
    x"1AF4EFDA",
    x"1AF4903F",
    x"1AF430CA",
    x"1AF3D179",
    x"1AF3724E",
    x"1AF31348",
    x"1AF2B467",
    x"1AF255AB",
    x"1AF1F714",
    x"1AF198A2",
    x"1AF13A55",
    x"1AF0DC2C",
    x"1AF07E29",
    x"1AF0204A",
    x"1AEFC28F",
    x"1AEF64FA",
    x"1AEF0788",
    x"1AEEAA3C",
    x"1AEE4D13",
    x"1AEDF00F",
    x"1AED9330",
    x"1AED3674",
    x"1AECD9DD",
    x"1AEC7D6A",
    x"1AEC211B",
    x"1AEBC4F0",
    x"1AEB68E9",
    x"1AEB0D06",
    x"1AEAB147",
    x"1AEA55AC",
    x"1AE9FA34",
    x"1AE99EE0",
    x"1AE943B0",
    x"1AE8E8A3",
    x"1AE88DBA",
    x"1AE832F5",
    x"1AE7D853",
    x"1AE77DD4",
    x"1AE72378",
    x"1AE6C940",
    x"1AE66F2B",
    x"1AE61539",
    x"1AE5BB6A",
    x"1AE561BF",
    x"1AE50836",
    x"1AE4AED0",
    x"1AE4558D",
    x"1AE3FC6D",
    x"1AE3A370",
    x"1AE34A96",
    x"1AE2F1DE",
    x"1AE29949",
    x"1AE240D6",
    x"1AE1E886",
    x"1AE19058",
    x"1AE1384D",
    x"1AE0E064",
    x"1AE0889E",
    x"1AE030FA",
    x"1ADFD978",
    x"1ADF8218",
    x"1ADF2ADA",
    x"1ADED3BE",
    x"1ADE7CC5",
    x"1ADE25ED",
    x"1ADDCF37",
    x"1ADD78A3",
    x"1ADD2231",
    x"1ADCCBE0",
    x"1ADC75B1",
    x"1ADC1FA4",
    x"1ADBC9B9",
    x"1ADB73EF",
    x"1ADB1E46",
    x"1ADAC8BF",
    x"1ADA7359",
    x"1ADA1E15",
    x"1AD9C8F2",
    x"1AD973F0",
    x"1AD91F0F",
    x"1AD8CA50",
    x"1AD875B1",
    x"1AD82134",
    x"1AD7CCD7",
    x"1AD7789B",
    x"1AD72481",
    x"1AD6D087",
    x"1AD67CAE",
    x"1AD628F6",
    x"1AD5D55E",
    x"1AD581E7",
    x"1AD52E90",
    x"1AD4DB5A",
    x"1AD48845",
    x"1AD43550",
    x"1AD3E27B",
    x"1AD38FC7",
    x"1AD33D33",
    x"1AD2EABF",
    x"1AD2986C",
    x"1AD24638",
    x"1AD1F425",
    x"1AD1A231",
    x"1AD1505E",
    x"1AD0FEAB",
    x"1AD0AD17",
    x"1AD05BA3",
    x"1AD00A4F",
    x"1ACFB91B",
    x"1ACF6807",
    x"1ACF1712",
    x"1ACEC63D",
    x"1ACE7587",
    x"1ACE24F1",
    x"1ACDD47A",
    x"1ACD8423",
    x"1ACD33EB",
    x"1ACCE3D2",
    x"1ACC93D9",
    x"1ACC43FF",
    x"1ACBF444",
    x"1ACBA4A8",
    x"1ACB552B",
    x"1ACB05CD",
    x"1ACAB68F",
    x"1ACA676F",
    x"1ACA186E",
    x"1AC9C98C",
    x"1AC97AC8",
    x"1AC92C24",
    x"1AC8DD9E",
    x"1AC88F37",
    x"1AC840EE",
    x"1AC7F2C4",
    x"1AC7A4B8",
    x"1AC756CB",
    x"1AC708FC",
    x"1AC6BB4C",
    x"1AC66DBA",
    x"1AC62046",
    x"1AC5D2F1",
    x"1AC585B9",
    x"1AC538A0",
    x"1AC4EBA5",
    x"1AC49EC8",
    x"1AC45209",
    x"1AC40568",
    x"1AC3B8E5",
    x"1AC36C80",
    x"1AC32038",
    x"1AC2D40E",
    x"1AC28802",
    x"1AC23C14",
    x"1AC1F044",
    x"1AC1A490",
    x"1AC158FB",
    x"1AC10D83",
    x"1AC0C228",
    x"1AC076EB",
    x"1AC02BCB",
    x"1ABFE0C9",
    x"1ABF95E4",
    x"1ABF4B1C",
    x"1ABF0071",
    x"1ABEB5E4",
    x"1ABE6B73",
    x"1ABE2120",
    x"1ABDD6E9",
    x"1ABD8CD0",
    x"1ABD42D3",
    x"1ABCF8F3",
    x"1ABCAF31",
    x"1ABC658B",
    x"1ABC1C01",
    x"1ABBD295",
    x"1ABB8945",
    x"1ABB4011",
    x"1ABAF6FB",
    x"1ABAAE00",
    x"1ABA6523",
    x"1ABA1C61",
    x"1AB9D3BD",
    x"1AB98B34",
    x"1AB942C8",
    x"1AB8FA78",
    x"1AB8B244",
    x"1AB86A2C",
    x"1AB82231",
    x"1AB7DA52",
    x"1AB7928F",
    x"1AB74AE7",
    x"1AB7035C",
    x"1AB6BBED",
    x"1AB67499",
    x"1AB62D62",
    x"1AB5E646",
    x"1AB59F46",
    x"1AB55861",
    x"1AB51199",
    x"1AB4CAEB",
    x"1AB4845A",
    x"1AB43DE4",
    x"1AB3F78A",
    x"1AB3B14B",
    x"1AB36B27",
    x"1AB3251F",
    x"1AB2DF32",
    x"1AB29961",
    x"1AB253AA",
    x"1AB20E0F",
    x"1AB1C88F",
    x"1AB1832A",
    x"1AB13DE1",
    x"1AB0F8B2",
    x"1AB0B39E",
    x"1AB06EA6",
    x"1AB029C8",
    x"1AAFE505",
    x"1AAFA05D",
    x"1AAF5BD0",
    x"1AAF175D",
    x"1AAED306",
    x"1AAE8EC8",
    x"1AAE4AA6",
    x"1AAE069E",
    x"1AADC2B1",
    x"1AAD7EDE",
    x"1AAD3B26",
    x"1AACF788",
    x"1AACB404",
    x"1AAC709B",
    x"1AAC2D4C",
    x"1AABEA18",
    x"1AABA6FD",
    x"1AAB63FD",
    x"1AAB2117",
    x"1AAADE4B",
    x"1AAA9B9A",
    x"1AAA5902",
    x"1AAA1684",
    x"1AA9D420",
    x"1AA991D6",
    x"1AA94FA6",
    x"1AA90D90",
    x"1AA8CB94",
    x"1AA889B1",
    x"1AA847E8",
    x"1AA80639",
    x"1AA7C4A3",
    x"1AA78327",
    x"1AA741C5",
    x"1AA7007C",
    x"1AA6BF4C",
    x"1AA67E36",
    x"1AA63D3A",
    x"1AA5FC56",
    x"1AA5BB8D",
    x"1AA57ADC",
    x"1AA53A45",
    x"1AA4F9C6",
    x"1AA4B961",
    x"1AA47916",
    x"1AA438E3",
    x"1AA3F8C9",
    x"1AA3B8C8",
    x"1AA378E1",
    x"1AA33912",
    x"1AA2F95C",
    x"1AA2B9BF",
    x"1AA27A3B",
    x"1AA23AD0",
    x"1AA1FB7D",
    x"1AA1BC43",
    x"1AA17D22",
    x"1AA13E19",
    x"1AA0FF29",
    x"1AA0C052",
    x"1AA08193",
    x"1AA042ED",
    x"1AA0045F",
    x"1A9FC5E9",
    x"1A9F878C",
    x"1A9F4947",
    x"1A9F0B1B",
    x"1A9ECD07",
    x"1A9E8F0B",
    x"1A9E5127",
    x"1A9E135B",
    x"1A9DD5A8",
    x"1A9D980C",
    x"1A9D5A89",
    x"1A9D1D1E",
    x"1A9CDFCA",
    x"1A9CA28F",
    x"1A9C656B",
    x"1A9C2860",
    x"1A9BEB6C",
    x"1A9BAE90",
    x"1A9B71CB",
    x"1A9B351F",
    x"1A9AF88A",
    x"1A9ABC0D",
    x"1A9A7FA7",
    x"1A9A4359",
    x"1A9A0722",
    x"1A99CB03",
    x"1A998EFC",
    x"1A99530C",
    x"1A991733",
    x"1A98DB71",
    x"1A989FC7",
    x"1A986435",
    x"1A9828B9",
    x"1A97ED55",
    x"1A97B208",
    x"1A9776D2",
    x"1A973BB3",
    x"1A9700AB",
    x"1A96C5BA",
    x"1A968AE0",
    x"1A96501E",
    x"1A961572",
    x"1A95DADD",
    x"1A95A05F",
    x"1A9565F8",
    x"1A952BA7",
    x"1A94F16E",
    x"1A94B74B",
    x"1A947D3E",
    x"1A944349",
    x"1A94096A",
    x"1A93CFA1",
    x"1A9395F0",
    x"1A935C54",
    x"1A9322CF",
    x"1A92E961",
    x"1A92B009",
    x"1A9276C7",
    x"1A923D9C",
    x"1A920487",
    x"1A91CB89",
    x"1A9192A0",
    x"1A9159CE",
    x"1A912112",
    x"1A90E86C",
    x"1A90AFDD",
    x"1A907763",
    x"1A903EFF",
    x"1A9006B2",
    x"1A8FCE7A",
    x"1A8F9658",
    x"1A8F5E4D",
    x"1A8F2657",
    x"1A8EEE77",
    x"1A8EB6AC",
    x"1A8E7EF8",
    x"1A8E4759",
    x"1A8E0FD0",
    x"1A8DD85D",
    x"1A8DA0FF",
    x"1A8D69B7",
    x"1A8D3284",
    x"1A8CFB67",
    x"1A8CC460",
    x"1A8C8D6E",
    x"1A8C5692",
    x"1A8C1FCA",
    x"1A8BE919",
    x"1A8BB27C",
    x"1A8B7BF5",
    x"1A8B4583",
    x"1A8B0F27",
    x"1A8AD8E0",
    x"1A8AA2AD",
    x"1A8A6C91",
    x"1A8A3689",
    x"1A8A0096",
    x"1A89CAB8",
    x"1A8994F0",
    x"1A895F3C",
    x"1A89299D",
    x"1A88F413",
    x"1A88BE9E",
    x"1A88893E",
    x"1A8853F3",
    x"1A881EBD",
    x"1A87E99B",
    x"1A87B48E",
    x"1A877F96",
    x"1A874AB3",
    x"1A8715E4",
    x"1A86E129",
    x"1A86AC84",
    x"1A8677F3",
    x"1A864376",
    x"1A860F0E",
    x"1A85DABA",
    x"1A85A67B",
    x"1A857250",
    x"1A853E3A",
    x"1A850A38",
    x"1A84D64A",
    x"1A84A270",
    x"1A846EAB",
    x"1A843AFA",
    x"1A84075D",
    x"1A83D3D4",
    x"1A83A05F",
    x"1A836CFF",
    x"1A8339B2",
    x"1A83067A",
    x"1A82D355",
    x"1A82A044",
    x"1A826D48",
    x"1A823A5F",
    x"1A82078A",
    x"1A81D4C9",
    x"1A81A21C",
    x"1A816F82",
    x"1A813CFD",
    x"1A810A8B",
    x"1A80D82D",
    x"1A80A5E2",
    x"1A8073AB",
    x"1A804188",
    x"1A800F78",
    x"1A7FBAF7",
    x"1A7F5725",
    x"1A7EF37B",
    x"1A7E8FF7",
    x"1A7E2C9A",
    x"1A7DC964",
    x"1A7D6655",
    x"1A7D036C",
    x"1A7CA0AA",
    x"1A7C3E0F",
    x"1A7BDB9A",
    x"1A7B794B",
    x"1A7B1723",
    x"1A7AB521",
    x"1A7A5345",
    x"1A79F190",
    x"1A799001",
    x"1A792E98",
    x"1A78CD54",
    x"1A786C37",
    x"1A780B40",
    x"1A77AA6E",
    x"1A7749C3",
    x"1A76E93D",
    x"1A7688DC",
    x"1A7628A2",
    x"1A75C88D",
    x"1A75689D",
    x"1A7508D3",
    x"1A74A92E",
    x"1A7449AF",
    x"1A73EA55",
    x"1A738B20",
    x"1A732C10",
    x"1A72CD25",
    x"1A726E60",
    x"1A720FBF",
    x"1A71B143",
    x"1A7152EC",
    x"1A70F4BA",
    x"1A7096AD",
    x"1A7038C5",
    x"1A6FDB01",
    x"1A6F7D62",
    x"1A6F1FE7",
    x"1A6EC291",
    x"1A6E655F",
    x"1A6E0851",
    x"1A6DAB68",
    x"1A6D4EA3",
    x"1A6CF203",
    x"1A6C9586",
    x"1A6C392E",
    x"1A6BDCFA",
    x"1A6B80E9",
    x"1A6B24FD",
    x"1A6AC934",
    x"1A6A6D90",
    x"1A6A120F",
    x"1A69B6B2",
    x"1A695B78",
    x"1A690062",
    x"1A68A570",
    x"1A684AA1",
    x"1A67EFF5",
    x"1A67956D",
    x"1A673B09",
    x"1A66E0C7",
    x"1A6686A9",
    x"1A662CAE",
    x"1A65D2D6",
    x"1A657921",
    x"1A651F8F",
    x"1A64C621",
    x"1A646CD5",
    x"1A6413AC",
    x"1A63BAA5",
    x"1A6361C2",
    x"1A630901",
    x"1A62B063",
    x"1A6257E7",
    x"1A61FF8E",
    x"1A61A757",
    x"1A614F43",
    x"1A60F751",
    x"1A609F82",
    x"1A6047D5",
    x"1A5FF04A",
    x"1A5F98E1",
    x"1A5F419A",
    x"1A5EEA76",
    x"1A5E9373",
    x"1A5E3C93",
    x"1A5DE5D4",
    x"1A5D8F37",
    x"1A5D38BC",
    x"1A5CE263",
    x"1A5C8C2B",
    x"1A5C3615",
    x"1A5BE021",
    x"1A5B8A4E",
    x"1A5B349D",
    x"1A5ADF0D",
    x"1A5A899E",
    x"1A5A3451",
    x"1A59DF26",
    x"1A598A1B",
    x"1A593532",
    x"1A58E069",
    x"1A588BC2",
    x"1A58373C",
    x"1A57E2D7",
    x"1A578E93",
    x"1A573A70",
    x"1A56E66D",
    x"1A56928C",
    x"1A563ECB",
    x"1A55EB2B",
    x"1A5597AB",
    x"1A55444C",
    x"1A54F10E",
    x"1A549DF0",
    x"1A544AF2",
    x"1A53F815",
    x"1A53A559",
    x"1A5352BC",
    x"1A530040",
    x"1A52ADE4",
    x"1A525BA8",
    x"1A52098C",
    x"1A51B791",
    x"1A5165B5",
    x"1A5113F9",
    x"1A50C25D",
    x"1A5070E1",
    x"1A501F85",
    x"1A4FCE49",
    x"1A4F7D2C",
    x"1A4F2C2F",
    x"1A4EDB51",
    x"1A4E8A93",
    x"1A4E39F5",
    x"1A4DE976",
    x"1A4D9917",
    x"1A4D48D6",
    x"1A4CF8B6",
    x"1A4CA8B4",
    x"1A4C58D2",
    x"1A4C090F",
    x"1A4BB96B",
    x"1A4B69E6",
    x"1A4B1A80",
    x"1A4ACB39",
    x"1A4A7C11",
    x"1A4A2D08",
    x"1A49DE1E",
    x"1A498F53",
    x"1A4940A6",
    x"1A48F218",
    x"1A48A3A9",
    x"1A485558",
    x"1A480726",
    x"1A47B913",
    x"1A476B1E",
    x"1A471D47",
    x"1A46CF8F",
    x"1A4681F5",
    x"1A463479",
    x"1A45E71C",
    x"1A4599DD",
    x"1A454CBC",
    x"1A44FFB9",
    x"1A44B2D4",
    x"1A44660D",
    x"1A441964",
    x"1A43CCD9",
    x"1A43806C",
    x"1A43341D",
    x"1A42E7EB",
    x"1A429BD8",
    x"1A424FE1",
    x"1A420409",
    x"1A41B84E",
    x"1A416CB1",
    x"1A412131",
    x"1A40D5CF",
    x"1A408A8A",
    x"1A403F63",
    x"1A3FF459",
    x"1A3FA96C",
    x"1A3F5E9C",
    x"1A3F13EA",
    x"1A3EC955",
    x"1A3E7EDD",
    x"1A3E3482",
    x"1A3DEA44",
    x"1A3DA023",
    x"1A3D561F",
    x"1A3D0C37",
    x"1A3CC26D",
    x"1A3C78BF",
    x"1A3C2F2F",
    x"1A3BE5BB",
    x"1A3B9C63",
    x"1A3B5328",
    x"1A3B0A0A",
    x"1A3AC109",
    x"1A3A7823",
    x"1A3A2F5B",
    x"1A39E6AE",
    x"1A399E1E",
    x"1A3955AB",
    x"1A390D53",
    x"1A38C518",
    x"1A387CF9",
    x"1A3834F7",
    x"1A37ED10",
    x"1A37A546",
    x"1A375D97",
    x"1A371604",
    x"1A36CE8E",
    x"1A368733",
    x"1A363FF4",
    x"1A35F8D1",
    x"1A35B1CA",
    x"1A356ADE",
    x"1A35240E",
    x"1A34DD5A",
    x"1A3496C1",
    x"1A345044",
    x"1A3409E3",
    x"1A33C39C",
    x"1A337D72",
    x"1A333762",
    x"1A32F16E",
    x"1A32AB96",
    x"1A3265D8",
    x"1A322036",
    x"1A31DAAF",
    x"1A319543",
    x"1A314FF3",
    x"1A310ABD",
    x"1A30C5A2",
    x"1A3080A2",
    x"1A303BBE",
    x"1A2FF6F4",
    x"1A2FB245",
    x"1A2F6DB0",
    x"1A2F2937",
    x"1A2EE4D8",
    x"1A2EA094",
    x"1A2E5C6B",
    x"1A2E185C",
    x"1A2DD468",
    x"1A2D908E",
    x"1A2D4CCF",
    x"1A2D092A",
    x"1A2CC5A0",
    x"1A2C8230",
    x"1A2C3EDA",
    x"1A2BFB9E",
    x"1A2BB87D",
    x"1A2B7576",
    x"1A2B328A",
    x"1A2AEFB7",
    x"1A2AACFE",
    x"1A2A6A60",
    x"1A2A27DB",
    x"1A29E571",
    x"1A29A320",
    x"1A2960E9",
    x"1A291ECC",
    x"1A28DCC9",
    x"1A289AE0",
    x"1A285910",
    x"1A28175A",
    x"1A27D5BE",
    x"1A27943B",
    x"1A2752D2",
    x"1A271182",
    x"1A26D04C",
    x"1A268F30",
    x"1A264E2C",
    x"1A260D42",
    x"1A25CC72",
    x"1A258BBB",
    x"1A254B1D",
    x"1A250A98",
    x"1A24CA2D",
    x"1A2489DA",
    x"1A2449A1",
    x"1A240981",
    x"1A23C979",
    x"1A23898B",
    x"1A2349B6",
    x"1A2309FA",
    x"1A22CA56",
    x"1A228ACB",
    x"1A224B5A",
    x"1A220C01",
    x"1A21CCC0",
    x"1A218D99",
    x"1A214E8A",
    x"1A210F93",
    x"1A20D0B5",
    x"1A2091F0",
    x"1A205343",
    x"1A2014AF",
    x"1A1FD633",
    x"1A1F97D0",
    x"1A1F5985",
    x"1A1F1B52",
    x"1A1EDD37",
    x"1A1E9F35",
    x"1A1E614B",
    x"1A1E2379",
    x"1A1DE5BF",
    x"1A1DA81D",
    x"1A1D6A94",
    x"1A1D2D22",
    x"1A1CEFC9",
    x"1A1CB287",
    x"1A1C755D",
    x"1A1C384B",
    x"1A1BFB51",
    x"1A1BBE6F",
    x"1A1B81A4",
    x"1A1B44F1",
    x"1A1B0856",
    x"1A1ACBD3",
    x"1A1A8F67",
    x"1A1A5313",
    x"1A1A16D6",
    x"1A19DAB1",
    x"1A199EA3",
    x"1A1962AD",
    x"1A1926CE",
    x"1A18EB07",
    x"1A18AF57",
    x"1A1873BE",
    x"1A18383C",
    x"1A17FCD2",
    x"1A17C17F",
    x"1A178643",
    x"1A174B1E",
    x"1A171010",
    x"1A16D519",
    x"1A169A39",
    x"1A165F71",
    x"1A1624BF",
    x"1A15EA24",
    x"1A15AFA0",
    x"1A157533",
    x"1A153ADC",
    x"1A15009D",
    x"1A14C674",
    x"1A148C62",
    x"1A145266",
    x"1A141881",
    x"1A13DEB3",
    x"1A13A4FB",
    x"1A136B5A",
    x"1A1331CF",
    x"1A12F85B",
    x"1A12BEFD",
    x"1A1285B6",
    x"1A124C85",
    x"1A12136A",
    x"1A11DA66",
    x"1A11A178",
    x"1A1168A0",
    x"1A112FDE",
    x"1A10F732",
    x"1A10BE9D",
    x"1A10861D",
    x"1A104DB4",
    x"1A101561",
    x"1A0FDD23",
    x"1A0FA4FC",
    x"1A0F6CEA",
    x"1A0F34EF",
    x"1A0EFD09",
    x"1A0EC539",
    x"1A0E8D7F",
    x"1A0E55DA",
    x"1A0E1E4C",
    x"1A0DE6D3",
    x"1A0DAF6F",
    x"1A0D7822",
    x"1A0D40EA",
    x"1A0D09C7",
    x"1A0CD2BA",
    x"1A0C9BC2",
    x"1A0C64E0",
    x"1A0C2E13",
    x"1A0BF75C",
    x"1A0BC0BA",
    x"1A0B8A2E",
    x"1A0B53B6",
    x"1A0B1D54",
    x"1A0AE707",
    x"1A0AB0D0",
    x"1A0A7AAD",
    x"1A0A44A0",
    x"1A0A0EA8",
    x"1A09D8C4",
    x"1A09A2F6",
    x"1A096D3D",
    x"1A093799",
    x"1A09020A",
    x"1A08CC8F",
    x"1A08972A",
    x"1A0861D9",
    x"1A082C9D",
    x"1A07F776",
    x"1A07C264",
    x"1A078D66",
    x"1A07587E",
    x"1A0723A9",
    x"1A06EEEA",
    x"1A06BA3F",
    x"1A0685A8",
    x"1A065126",
    x"1A061CB9",
    x"1A05E860",
    x"1A05B41B",
    x"1A057FEB",
    x"1A054BCF",
    x"1A0517C8",
    x"1A04E3D5",
    x"1A04AFF6",
    x"1A047C2B",
    x"1A044875",
    x"1A0414D3",
    x"1A03E144",
    x"1A03ADCB",
    x"1A037A65",
    x"1A034713",
    x"1A0313D5",
    x"1A02E0AB",
    x"1A02AD96",
    x"1A027A94",
    x"1A0247A6",
    x"1A0214CC",
    x"1A01E206",
    x"1A01AF53",
    x"1A017CB5",
    x"1A014A2A",
    x"1A0117B3",
    x"1A00E54F",
    x"1A00B300",
    x"1A0080C3",
    x"1A004E9B",
    x"1A001C86",
    x"19FFD509",
    x"19FF712E",
    x"19FF0D79",
    x"19FEA9EB",
    x"19FE4684",
    x"19FDE344",
    x"19FD802A",
    x"19FD1D38",
    x"19FCBA6C",
    x"19FC57C6",
    x"19FBF547",
    x"19FB92EE",
    x"19FB30BC",
    x"19FACEB0",
    x"19FA6CCB",
    x"19FA0B0B",
    x"19F9A972",
    x"19F947FF",
    x"19F8E6B2",
    x"19F8858B",
    x"19F82489",
    x"19F7C3AE",
    x"19F762F9",
    x"19F70269",
    x"19F6A1FF",
    x"19F641BA",
    x"19F5E19B",
    x"19F581A2",
    x"19F521CE",
    x"19F4C21F",
    x"19F46296",
    x"19F40332",
    x"19F3A3F4",
    x"19F344DA",
    x"19F2E5E6",
    x"19F28717",
    x"19F2286C",
    x"19F1C9E7",
    x"19F16B87",
    x"19F10D4B",
    x"19F0AF34",
    x"19F05142",
    x"19EFF375",
    x"19EF95CC",
    x"19EF3848",
    x"19EEDAE8",
    x"19EE7DAD",
    x"19EE2096",
    x"19EDC3A3",
    x"19ED66D5",
    x"19ED0A2B",
    x"19ECADA5",
    x"19EC5143",
    x"19EBF505",
    x"19EB98EC",
    x"19EB3CF6",
    x"19EAE124",
    x"19EA8576",
    x"19EA29EC",
    x"19E9CE85",
    x"19E97342",
    x"19E91823",
    x"19E8BD28",
    x"19E8624F",
    x"19E8079B",
    x"19E7AD09",
    x"19E7529C",
    x"19E6F851",
    x"19E69E2A",
    x"19E64425",
    x"19E5EA44",
    x"19E59086",
    x"19E536EB",
    x"19E4DD73",
    x"19E4841E",
    x"19E42AEC",
    x"19E3D1DD",
    x"19E378F0",
    x"19E32026",
    x"19E2C77F",
    x"19E26EFA",
    x"19E21698",
    x"19E1BE59",
    x"19E1663C",
    x"19E10E41",
    x"19E0B668",
    x"19E05EB2",
    x"19E0071E",
    x"19DFAFAD",
    x"19DF585D",
    x"19DF0130",
    x"19DEAA24",
    x"19DE533B",
    x"19DDFC73",
    x"19DDA5CD",
    x"19DD4F4A",
    x"19DCF8E8",
    x"19DCA2A7",
    x"19DC4C88",
    x"19DBF68B",
    x"19DBA0B0",
    x"19DB4AF6",
    x"19DAF55D",
    x"19DA9FE6",
    x"19DA4A90",
    x"19D9F55C",
    x"19D9A049",
    x"19D94B57",
    x"19D8F686",
    x"19D8A1D6",
    x"19D84D47",
    x"19D7F8DA",
    x"19D7A48D",
    x"19D75061",
    x"19D6FC56",
    x"19D6A86C",
    x"19D654A2",
    x"19D600FA",
    x"19D5AD72",
    x"19D55A0A",
    x"19D506C3",
    x"19D4B39D",
    x"19D46097",
    x"19D40DB1",
    x"19D3BAEC",
    x"19D36847",
    x"19D315C3",
    x"19D2C35E",
    x"19D2711A",
    x"19D21EF6",
    x"19D1CCF2",
    x"19D17B0E",
    x"19D1294A",
    x"19D0D7A6",
    x"19D08621",
    x"19D034BD",
    x"19CFE378",
    x"19CF9253",
    x"19CF414E",
    x"19CEF068",
    x"19CE9FA2",
    x"19CE4EFB",
    x"19CDFE74",
    x"19CDAE0C",
    x"19CD5DC4",
    x"19CD0D9B",
    x"19CCBD91",
    x"19CC6DA7",
    x"19CC1DDC",
    x"19CBCE30",
    x"19CB7EA3",
    x"19CB2F35",
    x"19CADFE6",
    x"19CA90B6",
    x"19CA41A5",
    x"19C9F2B3",
    x"19C9A3DF",
    x"19C9552A",
    x"19C90695",
    x"19C8B81D",
    x"19C869C5",
    x"19C81B8B",
    x"19C7CD6F",
    x"19C77F72",
    x"19C73194",
    x"19C6E3D3",
    x"19C69632",
    x"19C648AE",
    x"19C5FB49",
    x"19C5AE02",
    x"19C560D9",
    x"19C513CE",
    x"19C4C6E1",
    x"19C47A13",
    x"19C42D62",
    x"19C3E0CF",
    x"19C3945A",
    x"19C34803",
    x"19C2FBCA",
    x"19C2AFAF",
    x"19C263B1",
    x"19C217D1",
    x"19C1CC0E",
    x"19C18069",
    x"19C134E2",
    x"19C0E978",
    x"19C09E2B",
    x"19C052FC",
    x"19C007EB",
    x"19BFBCF6",
    x"19BF721F",
    x"19BF2765",
    x"19BEDCC8",
    x"19BE9248",
    x"19BE47E6",
    x"19BDFDA0",
    x"19BDB378",
    x"19BD696C",
    x"19BD1F7D",
    x"19BCD5AB",
    x"19BC8BF6",
    x"19BC425E",
    x"19BBF8E2",
    x"19BBAF84",
    x"19BB6641",
    x"19BB1D1C",
    x"19BAD413",
    x"19BA8B26",
    x"19BA4256",
    x"19B9F9A2",
    x"19B9B10B",
    x"19B96890",
    x"19B92031",
    x"19B8D7EF",
    x"19B88FC8",
    x"19B847BE",
    x"19B7FFD0",
    x"19B7B7FE",
    x"19B77049",
    x"19B728AF",
    x"19B6E131",
    x"19B699CF",
    x"19B65289",
    x"19B60B5E",
    x"19B5C450",
    x"19B57D5D",
    x"19B53686",
    x"19B4EFCA",
    x"19B4A92A",
    x"19B462A6",
    x"19B41C3D",
    x"19B3D5F0",
    x"19B38FBE",
    x"19B349A8",
    x"19B303AD",
    x"19B2BDCD",
    x"19B27808",
    x"19B2325F",
    x"19B1ECD1",
    x"19B1A75E",
    x"19B16206",
    x"19B11CC9",
    x"19B0D7A8",
    x"19B092A1",
    x"19B04DB5",
    x"19B008E4",
    x"19AFC42E",
    x"19AF7F93",
    x"19AF3B12",
    x"19AEF6AD",
    x"19AEB262",
    x"19AE6E31",
    x"19AE2A1C",
    x"19ADE620",
    x"19ADA240",
    x"19AD5E7A",
    x"19AD1ACE",
    x"19ACD73D",
    x"19AC93C6",
    x"19AC5069",
    x"19AC0D27",
    x"19ABC9FF",
    x"19AB86F1",
    x"19AB43FE",
    x"19AB0124",
    x"19AABE65",
    x"19AA7BBF",
    x"19AA3934",
    x"19A9F6C3",
    x"19A9B46B",
    x"19A9722E",
    x"19A9300A",
    x"19A8EE00",
    x"19A8AC10",
    x"19A86A3A",
    x"19A8287D",
    x"19A7E6DA",
    x"19A7A551",
    x"19A763E1",
    x"19A7228B",
    x"19A6E14E",
    x"19A6A02B",
    x"19A65F21",
    x"19A61E30",
    x"19A5DD59",
    x"19A59C9B",
    x"19A55BF7",
    x"19A51B6B",
    x"19A4DAF9",
    x"19A49AA0",
    x"19A45A61",
    x"19A41A3A",
    x"19A3DA2C",
    x"19A39A37",
    x"19A35A5C",
    x"19A31A99",
    x"19A2DAEF",
    x"19A29B5E",
    x"19A25BE5",
    x"19A21C86",
    x"19A1DD3F",
    x"19A19E11",
    x"19A15EFC",
    x"19A11FFF",
    x"19A0E11B",
    x"19A0A24F",
    x"19A0639C",
    x"19A02501",
    x"199FE67F",
    x"199FA815",
    x"199F69C3",
    x"199F2B8A",
    x"199EED69",
    x"199EAF61",
    x"199E7170",
    x"199E3398",
    x"199DF5D8",
    x"199DB830",
    x"199D7AA0",
    x"199D3D28",
    x"199CFFC8",
    x"199CC280",
    x"199C8550",
    x"199C4838",
    x"199C0B38",
    x"199BCE50",
    x"199B917F",
    x"199B54C6",
    x"199B1825",
    x"199ADB9B",
    x"199A9F29",
    x"199A62CF",
    x"199A268C",
    x"1999EA60",
    x"1999AE4D",
    x"19997250",
    x"1999366B",
    x"1998FA9E",
    x"1998BEE8",
    x"19988349",
    x"199847C1",
    x"19980C51",
    x"1997D0F7",
    x"199795B5",
    x"19975A8A",
    x"19971F77",
    x"1996E47A",
    x"1996A994",
    x"19966EC5",
    x"1996340D",
    x"1995F96D",
    x"1995BEE3",
    x"1995846F",
    x"19954A13",
    x"19950FCE",
    x"1994D59F",
    x"19949B87",
    x"19946185",
    x"1994279A",
    x"1993EDC6",
    x"1993B409",
    x"19937A62",
    x"199340D1",
    x"19930757",
    x"1992CDF3",
    x"199294A6",
    x"19925B6F",
    x"1992224F",
    x"1991E944",
    x"1991B050",
    x"19917773",
    x"19913EAB",
    x"199105FA",
    x"1990CD5E",
    x"199094D9",
    x"19905C6A",
    x"19902411",
    x"198FEBCE",
    x"198FB3A1",
    x"198F7B8A",
    x"198F4388",
    x"198F0B9D",
    x"198ED3C7",
    x"198E9C07",
    x"198E645D",
    x"198E2CC9",
    x"198DF54A",
    x"198DBDE1",
    x"198D868E",
    x"198D4F50",
    x"198D1828",
    x"198CE115",
    x"198CAA18",
    x"198C7330",
    x"198C3C5E",
    x"198C05A1",
    x"198BCEFA",
    x"198B9867",
    x"198B61EB",
    x"198B2B83",
    x"198AF531",
    x"198ABEF3",
    x"198A88CB",
    x"198A52B8",
    x"198A1CBB",
    x"1989E6D2",
    x"1989B0FE",
    x"19897B40",
    x"19894596",
    x"19891001",
    x"1988DA82",
    x"1988A517",
    x"19886FC1",
    x"19883A7F",
    x"19880553",
    x"1987D03B",
    x"19879B38",
    x"1987664A",
    x"19873170",
    x"1986FCAB",
    x"1986C7FB",
    x"1986935F",
    x"19865ED8",
    x"19862A65",
    x"1985F607",
    x"1985C1BD",
    x"19858D87",
    x"19855966",
    x"19852559",
    x"1984F161",
    x"1984BD7D",
    x"198489AD",
    x"198455F1",
    x"1984224A",
    x"1983EEB6",
    x"1983BB37",
    x"198387CC",
    x"19835475",
    x"19832132",
    x"1982EE03",
    x"1982BAE8",
    x"198287E1",
    x"198254EE",
    x"1982220F",
    x"1981EF43",
    x"1981BC8C",
    x"198189E8",
    x"19815758",
    x"198124DC",
    x"1980F273",
    x"1980C01E",
    x"19808DDD",
    x"19805BB0",
    x"19802996",
    x"197FEF1E",
    x"197F8B38",
    x"197F2779",
    x"197EC3E1",
    x"197E6070",
    x"197DFD26",
    x"197D9A02",
    x"197D3706",
    x"197CD42F",
    x"197C7180",
    x"197C0EF7",
    x"197BAC94",
    x"197B4A58",
    x"197AE842",
    x"197A8652",
    x"197A2489",
    x"1979C2E6",
    x"19796169",
    x"19790012",
    x"19789EE1",
    x"19783DD6",
    x"1977DCF0",
    x"19777C31",
    x"19771B97",
    x"1976BB23",
    x"19765AD5",
    x"1975FAAC",
    x"19759AA9",
    x"19753ACC",
    x"1974DB13",
    x"19747B80",
    x"19741C13",
    x"1973BCCB",
    x"19735DA7",
    x"1972FEA9",
    x"19729FD0",
    x"1972411C",
    x"1971E28D",
    x"19718423",
    x"197125DE",
    x"1970C7BE",
    x"197069C2",
    x"19700BEB",
    x"196FAE39",
    x"196F50AB",
    x"196EF342",
    x"196E95FD",
    x"196E38DD",
    x"196DDBE1",
    x"196D7F09",
    x"196D2255",
    x"196CC5C6",
    x"196C695B",
    x"196C0D14",
    x"196BB0F1",
    x"196B54F1",
    x"196AF916",
    x"196A9D5F",
    x"196A41CB",
    x"1969E65B",
    x"19698B0F",
    x"19692FE7",
    x"1968D4E2",
    x"19687A00",
    x"19681F42",
    x"1967C4A8",
    x"19676A31",
    x"19670FDD",
    x"1966B5AC",
    x"19665B9F",
    x"196601B5",
    x"1965A7EE",
    x"19654E4A",
    x"1964F4C8",
    x"19649B6A",
    x"1964422F",
    x"1963E917",
    x"19639021",
    x"1963374E",
    x"1962DE9E",
    x"19628610",
    x"19622DA5",
    x"1961D55C",
    x"19617D36",
    x"19612532",
    x"1960CD51",
    x"19607592",
    x"19601DF5",
    x"195FC67B",
    x"195F6F22",
    x"195F17EC",
    x"195EC0D7",
    x"195E69E5",
    x"195E1315",
    x"195DBC66",
    x"195D65DA",
    x"195D0F6F",
    x"195CB925",
    x"195C62FE",
    x"195C0CF8",
    x"195BB714",
    x"195B6151",
    x"195B0BB0",
    x"195AB630",
    x"195A60D1",
    x"195A0B94",
    x"1959B678",
    x"1959617E",
    x"19590CA4",
    x"1958B7EC",
    x"19586354",
    x"19580EDE",
    x"1957BA89",
    x"19576654",
    x"19571241",
    x"1956BE4E",
    x"19566A7C",
    x"195616CB",
    x"1955C33A",
    x"19556FCA",
    x"19551C7B",
    x"1954C94C",
    x"1954763E",
    x"19542350",
    x"1953D082",
    x"19537DD5",
    x"19532B48",
    x"1952D8DB",
    x"1952868E",
    x"19523462",
    x"1951E255",
    x"19519069",
    x"19513E9D",
    x"1950ECF0",
    x"19509B63",
    x"195049F7",
    x"194FF8AA",
    x"194FA77C",
    x"194F566F",
    x"194F0581",
    x"194EB4B2",
    x"194E6404",
    x"194E1374",
    x"194DC304",
    x"194D72B4",
    x"194D2283",
    x"194CD271",
    x"194C827E",
    x"194C32AB",
    x"194BE2F7",
    x"194B9362",
    x"194B43EC",
    x"194AF495",
    x"194AA55D",
    x"194A5643",
    x"194A0749",
    x"1949B86E",
    x"194969B1",
    x"19491B13",
    x"1948CC94",
    x"19487E33",
    x"19482FF1",
    x"1947E1CE",
    x"194793C9",
    x"194745E2",
    x"1946F81A",
    x"1946AA70",
    x"19465CE5",
    x"19460F78",
    x"1945C229",
    x"194574F8",
    x"194527E6",
    x"1944DAF1",
    x"19448E1A",
    x"19444162",
    x"1943F4C7",
    x"1943A84B",
    x"19435BEC",
    x"19430FAB",
    x"1942C388",
    x"19427782",
    x"19422B9A",
    x"1941DFD0",
    x"19419423",
    x"19414894",
    x"1940FD23",
    x"1940B1CF",
    x"19406698",
    x"19401B7E",
    x"193FD082",
    x"193F85A3",
    x"193F3AE2",
    x"193EF03D",
    x"193EA5B6",
    x"193E5B4C",
    x"193E10FF",
    x"193DC6CF",
    x"193D7CBB",
    x"193D32C5",
    x"193CE8EC",
    x"193C9F2F",
    x"193C558F",
    x"193C0C0C",
    x"193BC2A6",
    x"193B795C",
    x"193B302F",
    x"193AE71F",
    x"193A9E2B",
    x"193A5553",
    x"193A0C98",
    x"1939C3F9",
    x"19397B77",
    x"19393311",
    x"1938EAC7",
    x"1938A299",
    x"19385A88",
    x"19381293",
    x"1937CAB9",
    x"193782FC",
    x"19373B5B",
    x"1936F3D6",
    x"1936AC6C",
    x"1936651F",
    x"19361DED",
    x"1935D6D8",
    x"19358FDE",
    x"193548FF",
    x"1935023D",
    x"1934BB95",
    x"1934750A",
    x"19342E9A",
    x"1933E846",
    x"1933A20D",
    x"19335BEF",
    x"193315ED",
    x"1932D006",
    x"19328A3A",
    x"1932448A",
    x"1931FEF5",
    x"1931B97B",
    x"1931741C",
    x"19312ED8",
    x"1930E9AF",
    x"1930A4A1",
    x"19305FAE",
    x"19301AD7",
    x"192FD619",
    x"192F9177",
    x"192F4CF0",
    x"192F0883",
    x"192EC431",
    x"192E7FFA",
    x"192E3BDD",
    x"192DF7DB",
    x"192DB3F3",
    x"192D7026",
    x"192D2C74",
    x"192CE8DC",
    x"192CA55E",
    x"192C61FB",
    x"192C1EB1",
    x"192BDB83",
    x"192B986E",
    x"192B5573",
    x"192B1293",
    x"192ACFCD",
    x"192A8D21",
    x"192A4A8F",
    x"192A0816",
    x"1929C5B8",
    x"19298374",
    x"1929414A",
    x"1928FF39",
    x"1928BD42",
    x"19287B65",
    x"192839A2",
    x"1927F7F8",
    x"1927B668",
    x"192774F2",
    x"19273395",
    x"1926F251",
    x"1926B127",
    x"19267017",
    x"19262F20",
    x"1925EE42",
    x"1925AD7E",
    x"19256CD2",
    x"19252C41",
    x"1924EBC8",
    x"1924AB68",
    x"19246B22",
    x"19242AF5",
    x"1923EAE0",
    x"1923AAE5",
    x"19236B03",
    x"19232B39",
    x"1922EB89",
    x"1922ABF1",
    x"19226C73",
    x"19222D0D",
    x"1921EDC0",
    x"1921AE8B",
    x"19216F6F",
    x"1921306C",
    x"1920F181",
    x"1920B2AF",
    x"192073F6",
    x"19203555",
    x"191FF6CC",
    x"191FB85C",
    x"191F7A04",
    x"191F3BC4",
    x"191EFD9D",
    x"191EBF8E",
    x"191E8198",
    x"191E43B9",
    x"191E05F3",
    x"191DC844",
    x"191D8AAE",
    x"191D4D30",
    x"191D0FCA",
    x"191CD27C",
    x"191C9545",
    x"191C5827",
    x"191C1B21",
    x"191BDE32",
    x"191BA15B",
    x"191B649C",
    x"191B27F4",
    x"191AEB65",
    x"191AAEEC",
    x"191A728C",
    x"191A3643",
    x"1919FA11",
    x"1919BDF8",
    x"191981F5",
    x"1919460A",
    x"19190A36",
    x"1918CE7A",
    x"191892D5",
    x"19185747",
    x"19181BD1",
    x"1917E072",
    x"1917A529",
    x"191769F8",
    x"19172EDF",
    x"1916F3DC",
    x"1916B8F0",
    x"19167E1B",
    x"1916435E",
    x"191608B7",
    x"1915CE27",
    x"191593AE",
    x"1915594B",
    x"19151F00",
    x"1914E4CB",
    x"1914AAAD",
    x"191470A6",
    x"191436B5",
    x"1913FCDB",
    x"1913C318",
    x"1913896B",
    x"19134FD4",
    x"19131654",
    x"1912DCEB",
    x"1912A398",
    x"19126A5B",
    x"19123135",
    x"1911F824",
    x"1911BF2B",
    x"19118647",
    x"19114D7A",
    x"191114C3",
    x"1910DC22",
    x"1910A397",
    x"19106B22",
    x"191032C3",
    x"190FFA7A",
    x"190FC247",
    x"190F8A2A",
    x"190F5223",
    x"190F1A32",
    x"190EE257",
    x"190EAA91",
    x"190E72E1",
    x"190E3B47",
    x"190E03C3",
    x"190DCC55",
    x"190D94FC",
    x"190D5DB8",
    x"190D268A",
    x"190CEF72",
    x"190CB86F",
    x"190C8182",
    x"190C4AAA",
    x"190C13E8",
    x"190BDD3A",
    x"190BA6A3",
    x"190B7020",
    x"190B39B3",
    x"190B035B",
    x"190ACD18",
    x"190A96EB",
    x"190A60D3",
    x"190A2ACF",
    x"1909F4E1",
    x"1909BF08",
    x"19098944",
    x"19095395",
    x"19091DFB",
    x"1908E875",
    x"1908B305",
    x"19087DA9",
    x"19084863",
    x"19081331",
    x"1907DE14",
    x"1907A90B",
    x"19077418",
    x"19073F39",
    x"19070A6E",
    x"1906D5B8",
    x"1906A117",
    x"19066C8B",
    x"19063812",
    x"190603AF",
    x"1905CF60",
    x"19059B25",
    x"190566FE",
    x"190532EC",
    x"1904FEEF",
    x"1904CB05",
    x"19049730",
    x"1904636F",
    x"19042FC2",
    x"1903FC2A",
    x"1903C8A5",
    x"19039535",
    x"190361D9",
    x"19032E90",
    x"1902FB5C",
    x"1902C83C",
    x"19029530",
    x"19026238",
    x"19022F53",
    x"1901FC83",
    x"1901C9C6",
    x"1901971D",
    x"19016488",
    x"19013206",
    x"1900FF99",
    x"1900CD3F",
    x"19009AF8",
    x"190068C6",
    x"190036A6",
    x"1900049B",
    x"18FFA546",
    x"18FF417D",
    x"18FEDDDA",
    x"18FE7A5F",
    x"18FE170B",
    x"18FDB3DD",
    x"18FD50D6",
    x"18FCEDF6",
    x"18FC8B3C",
    x"18FC28A9",
    x"18FBC63D",
    x"18FB63F6",
    x"18FB01D6",
    x"18FA9FDD",
    x"18FA3E0A",
    x"18F9DC5C",
    x"18F97AD5",
    x"18F91974",
    x"18F8B839",
    x"18F85724",
    x"18F7F635",
    x"18F7956C",
    x"18F734C9",
    x"18F6D44B",
    x"18F673F3",
    x"18F613C0",
    x"18F5B3B3",
    x"18F553CC",
    x"18F4F40A",
    x"18F4946D",
    x"18F434F6",
    x"18F3D5A4",
    x"18F37677",
    x"18F3176F",
    x"18F2B88D",
    x"18F259CF",
    x"18F1FB36",
    x"18F19CC3",
    x"18F13E74",
    x"18F0E04A",
    x"18F08245",
    x"18F02464",
    x"18EFC6A8",
    x"18EF6911",
    x"18EF0B9E",
    x"18EEAE50",
    x"18EE5126",
    x"18EDF420",
    x"18ED973F",
    x"18ED3A82",
    x"18ECDDE9",
    x"18EC8175",
    x"18EC2524",
    x"18EBC8F8",
    x"18EB6CEF",
    x"18EB110B",
    x"18EAB54A",
    x"18EA59AD",
    x"18E9FE34",
    x"18E9A2DE",
    x"18E947AD",
    x"18E8EC9E",
    x"18E891B4",
    x"18E836ED",
    x"18E7DC49",
    x"18E781C8",
    x"18E7276B",
    x"18E6CD32",
    x"18E6731B",
    x"18E61928",
    x"18E5BF57",
    x"18E565AA",
    x"18E50C20",
    x"18E4B2B9",
    x"18E45974",
    x"18E40053",
    x"18E3A754",
    x"18E34E78",
    x"18E2F5BF",
    x"18E29D28",
    x"18E244B4",
    x"18E1EC62",
    x"18E19433",
    x"18E13C27",
    x"18E0E43C",
    x"18E08C74",
    x"18E034CE",
    x"18DFDD4B",
    x"18DF85EA",
    x"18DF2EAA",
    x"18DED78D",
    x"18DE8092",
    x"18DE29B9",
    x"18DDD301",
    x"18DD7C6C",
    x"18DD25F8",
    x"18DCCFA6",
    x"18DC7976",
    x"18DC2367",
    x"18DBCD7A",
    x"18DB77AF",
    x"18DB2205",
    x"18DACC7C",
    x"18DA7715",
    x"18DA21CF",
    x"18D9CCAA",
    x"18D977A7",
    x"18D922C5",
    x"18D8CE04",
    x"18D87964",
    x"18D824E5",
    x"18D7D087",
    x"18D77C4A",
    x"18D7282E",
    x"18D6D433",
    x"18D68058",
    x"18D62C9E",
    x"18D5D905",
    x"18D5858D",
    x"18D53235",
    x"18D4DEFE",
    x"18D48BE7",
    x"18D438F0",
    x"18D3E61A",
    x"18D39365",
    x"18D340CF",
    x"18D2EE5A",
    x"18D29C05",
    x"18D249D0",
    x"18D1F7BB",
    x"18D1A5C6",
    x"18D153F2",
    x"18D1023D",
    x"18D0B0A8",
    x"18D05F33",
    x"18D00DDD",
    x"18CFBCA8",
    x"18CF6B92",
    x"18CF1A9C",
    x"18CEC9C5",
    x"18CE790E",
    x"18CE2877",
    x"18CDD7FF",
    x"18CD87A6",
    x"18CD376D",
    x"18CCE753",
    x"18CC9758",
    x"18CC477C",
    x"18CBF7C0",
    x"18CBA823",
    x"18CB58A5",
    x"18CB0946",
    x"18CABA05",
    x"18CA6AE4",
    x"18CA1BE2",
    x"18C9CCFE",
    x"18C97E3A",
    x"18C92F94",
    x"18C8E10C",
    x"18C892A4",
    x"18C8445A",
    x"18C7F62E",
    x"18C7A822",
    x"18C75A33",
    x"18C70C63",
    x"18C6BEB1",
    x"18C6711E",
    x"18C623A9",
    x"18C5D652",
    x"18C5891A",
    x"18C53BFF",
    x"18C4EF03",
    x"18C4A224",
    x"18C45564",
    x"18C408C2",
    x"18C3BC3D",
    x"18C36FD7",
    x"18C3238E",
    x"18C2D763",
    x"18C28B55",
    x"18C23F66",
    x"18C1F394",
    x"18C1A7E0",
    x"18C15C49",
    x"18C110CF",
    x"18C0C574",
    x"18C07A35",
    x"18C02F14",
    x"18BFE410",
    x"18BF992A",
    x"18BF4E61",
    x"18BF03B5",
    x"18BEB926",
    x"18BE6EB4",
    x"18BE245F",
    x"18BDDA28",
    x"18BD900D",
    x"18BD460F",
    x"18BCFC2E",
    x"18BCB26A",
    x"18BC68C3",
    x"18BC1F38",
    x"18BBD5CA",
    x"18BB8C79",
    x"18BB4345",
    x"18BAFA2D",
    x"18BAB131",
    x"18BA6852",
    x"18BA1F90",
    x"18B9D6E9",
    x"18B98E60",
    x"18B945F2",
    x"18B8FDA1",
    x"18B8B56C",
    x"18B86D53",
    x"18B82557",
    x"18B7DD76",
    x"18B795B2",
    x"18B74E09",
    x"18B7067D",
    x"18B6BF0C",
    x"18B677B7",
    x"18B6307E",
    x"18B5E961",
    x"18B5A260",
    x"18B55B7B",
    x"18B514B1",
    x"18B4CE02",
    x"18B48770",
    x"18B440F9",
    x"18B3FA9D",
    x"18B3B45D",
    x"18B36E38",
    x"18B3282F",
    x"18B2E241",
    x"18B29C6E",
    x"18B256B6",
    x"18B2111A",
    x"18B1CB99",
    x"18B18633",
    x"18B140E8",
    x"18B0FBB8",
    x"18B0B6A3",
    x"18B071AA",
    x"18B02CCB",
    x"18AFE807",
    x"18AFA35D",
    x"18AF5ECF",
    x"18AF1A5B",
    x"18AED602",
    x"18AE91C4",
    x"18AE4DA0",
    x"18AE0997",
    x"18ADC5A9",
    x"18AD81D5",
    x"18AD3E1B",
    x"18ACFA7C",
    x"18ACB6F8",
    x"18AC738D",
    x"18AC303D",
    x"18ABED08",
    x"18ABA9EC",
    x"18AB66EB",
    x"18AB2404",
    x"18AAE137",
    x"18AA9E84",
    x"18AA5BEB",
    x"18AA196C",
    x"18A9D707",
    x"18A994BC",
    x"18A9528B",
    x"18A91074",
    x"18A8CE76",
    x"18A88C92",
    x"18A84AC8",
    x"18A80918",
    x"18A7C781",
    x"18A78604",
    x"18A744A0",
    x"18A70356",
    x"18A6C226",
    x"18A6810F",
    x"18A64011",
    x"18A5FF2D",
    x"18A5BE62",
    x"18A57DB0",
    x"18A53D17",
    x"18A4FC98",
    x"18A4BC32",
    x"18A47BE5",
    x"18A43BB1",
    x"18A3FB96",
    x"18A3BB95",
    x"18A37BAC",
    x"18A33BDC",
    x"18A2FC25",
    x"18A2BC87",
    x"18A27D02",
    x"18A23D95",
    x"18A1FE42",
    x"18A1BF07",
    x"18A17FE4",
    x"18A140DB",
    x"18A101EA",
    x"18A0C311",
    x"18A08451",
    x"18A045AA",
    x"18A0071B",
    x"189FC8A4",
    x"189F8A46",
    x"189F4C00",
    x"189F0DD3",
    x"189ECFBD",
    x"189E91C0",
    x"189E53DC",
    x"189E160F",
    x"189DD85A",
    x"189D9ABE",
    x"189D5D39",
    x"189D1FCD",
    x"189CE279",
    x"189CA53C",
    x"189C6817",
    x"189C2B0B",
    x"189BEE16",
    x"189BB139",
    x"189B7473",
    x"189B37C6",
    x"189AFB30",
    x"189ABEB1",
    x"189A824B",
    x"189A45FC",
    x"189A09C4",
    x"1899CDA4",
    x"1899919B",
    x"189955AA",
    x"189919D0",
    x"1898DE0E",
    x"1898A263",
    x"189866CF",
    x"18982B53",
    x"1897EFED",
    x"1897B49F",
    x"18977968",
    x"18973E48",
    x"18970340",
    x"1896C84E",
    x"18968D73",
    x"189652AF",
    x"18961802",
    x"1895DD6D",
    x"1895A2ED",
    x"18956885",
    x"18952E34",
    x"1894F3F9",
    x"1894B9D5",
    x"18947FC8",
    x"189445D1",
    x"18940BF1",
    x"1893D228",
    x"18939875",
    x"18935ED9",
    x"18932553",
    x"1892EBE4",
    x"1892B28B",
    x"18927948",
    x"1892401C",
    x"18920706",
    x"1891CE06",
    x"1891951D",
    x"18915C4A",
    x"1891238D",
    x"1890EAE6",
    x"1890B255",
    x"189079DB",
    x"18904176",
    x"18900928",
    x"188FD0EF",
    x"188F98CC",
    x"188F60C0",
    x"188F28C9",
    x"188EF0E8",
    x"188EB91D",
    x"188E8167",
    x"188E49C8",
    x"188E123E",
    x"188DDAC9",
    x"188DA36B",
    x"188D6C22",
    x"188D34EE",
    x"188CFDD0",
    x"188CC6C8",
    x"188C8FD5",
    x"188C58F7",
    x"188C222F",
    x"188BEB7D",
    x"188BB4DF",
    x"188B7E57",
    x"188B47E5",
    x"188B1187",
    x"188ADB3F",
    x"188AA50C",
    x"188A6EEE",
    x"188A38E5",
    x"188A02F2",
    x"1889CD13",
    x"18899749",
    x"18896195",
    x"18892BF5",
    x"1888F66A",
    x"1888C0F5",
    x"18888B94",
    x"18885648",
    x"18882110",
    x"1887EBEE",
    x"1887B6E0",
    x"188781E7",
    x"18874D02",
    x"18871833",
    x"1886E378",
    x"1886AED1",
    x"18867A3F",
    x"188645C1",
    x"18861158",
    x"1885DD04",
    x"1885A8C4",
    x"18857498",
    x"18854081",
    x"18850C7E",
    x"1884D88F",
    x"1884A4B4",
    x"188470EE",
    x"18843D3C",
    x"1884099E",
    x"1883D615",
    x"1883A29F",
    x"18836F3E",
    x"18833BF0",
    x"188308B7",
    x"1882D591",
    x"1882A280",
    x"18826F82",
    x"18823C99",
    x"188209C3",
    x"1881D701",
    x"1881A453",
    x"188171B9",
    x"18813F32",
    x"18810CBF",
    x"1880DA60",
    x"1880A815",
    x"188075DD",
    x"188043B9",
    x"188011A8",
    x"187FBF56",
    x"187F5B82",
    x"187EF7D6",
    x"187E9451",
    x"187E30F2",
    x"187DCDBB",
    x"187D6AAA",
    x"187D07BF",
    x"187CA4FB",
    x"187C425E",
    x"187BDFE8",
    x"187B7D97",
    x"187B1B6D",
    x"187AB96A",
    x"187A578D",
    x"1879F5D5",
    x"18799445",
    x"187932DA",
    x"1878D195",
    x"18787076",
    x"18780F7D",
    x"1877AEAA",
    x"18774DFC",
    x"1876ED75",
    x"18768D13",
    x"18762CD7",
    x"1875CCC0",
    x"18756CCF",
    x"18750D03",
    x"1874AD5C",
    x"18744DDB",
    x"1873EE80",
    x"18738F49",
    x"18733038",
    x"1872D14B",
    x"18727284",
    x"187213E2",
    x"1871B565",
    x"1871570C",
    x"1870F8D8",
    x"18709ACA",
    x"18703CE0",
    x"186FDF1A",
    x"186F8179",
    x"186F23FD",
    x"186EC6A5",
    x"186E6972",
    x"186E0C63",
    x"186DAF78",
    x"186D52B2",
    x"186CF60F",
    x"186C9991",
    x"186C3D37",
    x"186BE101",
    x"186B84F0",
    x"186B2902",
    x"186ACD38",
    x"186A7191",
    x"186A160F",
    x"1869BAB0",
    x"18695F75",
    x"1869045D",
    x"1868A969",
    x"18684E99",
    x"1867F3EC",
    x"18679962",
    x"18673EFC",
    x"1866E4B9",
    x"18668A9A",
    x"1866309D",
    x"1865D6C4",
    x"18657D0D",
    x"1865237A",
    x"1864CA09",
    x"186470BC",
    x"18641791",
    x"1863BE8A",
    x"186365A4",
    x"18630CE2",
    x"1862B442",
    x"18625BC5",
    x"1862036B",
    x"1861AB33",
    x"1861531D",
    x"1860FB2A",
    x"1860A359",
    x"18604BAA",
    x"185FF41E",
    x"185F9CB3",
    x"185F456B",
    x"185EEE45",
    x"185E9741",
    x"185E405F",
    x"185DE99F",
    x"185D9300",
    x"185D3C84",
    x"185CE629",
    x"185C8FF0",
    x"185C39D9",
    x"185BE3E3",
    x"185B8E0E",
    x"185B385C",
    x"185AE2CA",
    x"185A8D5B",
    x"185A380C",
    x"1859E2DF",
    x"18598DD3",
    x"185938E8",
    x"1858E41E",
    x"18588F76",
    x"18583AEE",
    x"1857E688",
    x"18579242",
    x"18573E1D",
    x"1856EA19",
    x"18569636",
    x"18564274",
    x"1855EED2",
    x"18559B52",
    x"185547F1",
    x"1854F4B1",
    x"1854A192",
    x"18544E93",
    x"1853FBB5",
    x"1853A8F6",
    x"18535659",
    x"185303DB",
    x"1852B17D",
    x"18525F40",
    x"18520D23",
    x"1851BB26",
    x"18516949",
    x"1851178C",
    x"1850C5EE",
    x"18507471",
    x"18502313",
    x"184FD1D6",
    x"184F80B7",
    x"184F2FB9",
    x"184EDEDA",
    x"184E8E1B",
    x"184E3D7B",
    x"184DECFB",
    x"184D9C9A",
    x"184D4C59",
    x"184CFC36",
    x"184CAC33",
    x"184C5C50",
    x"184C0C8B",
    x"184BBCE6",
    x"184B6D60",
    x"184B1DF9",
    x"184ACEB0",
    x"184A7F87",
    x"184A307D",
    x"1849E191",
    x"184992C4",
    x"18494416",
    x"1848F587",
    x"1848A717",
    x"184858C5",
    x"18480A91",
    x"1847BC7C",
    x"18476E86",
    x"184720AE",
    x"1846D2F4",
    x"18468559",
    x"184637DC",
    x"1845EA7E",
    x"18459D3D",
    x"1845501B",
    x"18450316",
    x"1844B630",
    x"18446968",
    x"18441CBE",
    x"1843D032",
    x"184383C3",
    x"18433773",
    x"1842EB40",
    x"18429F2B",
    x"18425334",
    x"1842075A",
    x"1841BB9E",
    x"18416FFF",
    x"1841247E",
    x"1840D91B",
    x"18408DD5",
    x"184042AC",
    x"183FF7A1",
    x"183FACB2",
    x"183F61E2",
    x"183F172E",
    x"183ECC97",
    x"183E821E",
    x"183E37C2",
    x"183DED83",
    x"183DA360",
    x"183D595B",
    x"183D0F72",
    x"183CC5A7",
    x"183C7BF8",
    x"183C3266",
    x"183BE8F1",
    x"183B9F98",
    x"183B565C",
    x"183B0D3C",
    x"183AC43A",
    x"183A7B53",
    x"183A3289",
    x"1839E9DC",
    x"1839A14A",
    x"183958D6",
    x"1839107D",
    x"1838C841",
    x"18388021",
    x"1838381D",
    x"1837F035",
    x"1837A869",
    x"183760B9",
    x"18371925",
    x"1836D1AD",
    x"18368A52",
    x"18364311",
    x"1835FBED",
    x"1835B4E5",
    x"18356DF8",
    x"18352727",
    x"1834E071",
    x"183499D7",
    x"18345359",
    x"18340CF6",
    x"1833C6AF",
    x"18338083",
    x"18333A72",
    x"1832F47D",
    x"1832AEA3",
    x"183268E5",
    x"18322341",
    x"1831DDB9",
    x"1831984C",
    x"183152FA",
    x"18310DC3",
    x"1830C8A7",
    x"183083A7",
    x"18303EC1",
    x"182FF9F6",
    x"182FB545",
    x"182F70B0",
    x"182F2C35",
    x"182EE7D5",
    x"182EA390",
    x"182E5F66",
    x"182E1B56",
    x"182DD760",
    x"182D9385",
    x"182D4FC5",
    x"182D0C1F",
    x"182CC893",
    x"182C8522",
    x"182C41CB",
    x"182BFE8F",
    x"182BBB6D",
    x"182B7864",
    x"182B3576",
    x"182AF2A3",
    x"182AAFE9",
    x"182A6D49",
    x"182A2AC3",
    x"1829E858",
    x"1829A606",
    x"182963CE",
    x"182921B0",
    x"1828DFAC",
    x"18289DC1",
    x"18285BF0",
    x"18281A39",
    x"1827D89C",
    x"18279718",
    x"182755AE",
    x"1827145D",
    x"1826D326",
    x"18269208",
    x"18265104",
    x"18261019",
    x"1825CF47",
    x"18258E8F",
    x"18254DF0",
    x"18250D6A",
    x"1824CCFD",
    x"18248CAA",
    x"18244C70",
    x"18240C4E",
    x"1823CC46",
    x"18238C57",
    x"18234C80",
    x"18230CC3",
    x"1822CD1E",
    x"18228D93",
    x"18224E20",
    x"18220EC5",
    x"1821CF84",
    x"1821905B",
    x"1821514B",
    x"18211254",
    x"1820D375",
    x"182094AF",
    x"18205601",
    x"1820176B",
    x"181FD8EE",
    x"181F9A8A",
    x"181F5C3E",
    x"181F1E0A",
    x"181EDFEE",
    x"181EA1EB",
    x"181E6400",
    x"181E262D",
    x"181DE872",
    x"181DAACF",
    x"181D6D44",
    x"181D2FD2",
    x"181CF277",
    x"181CB534",
    x"181C7809",
    x"181C3AF7",
    x"181BFDFB",
    x"181BC118",
    x"181B844D",
    x"181B4799",
    x"181B0AFD",
    x"181ACE78",
    x"181A920B",
    x"181A55B6",
    x"181A1978",
    x"1819DD52",
    x"1819A143",
    x"1819654C",
    x"1819296C",
    x"1818EDA4",
    x"1818B1F3",
    x"18187659",
    x"18183AD6",
    x"1817FF6B",
    x"1817C417",
    x"181788DA",
    x"18174DB4",
    x"181712A5",
    x"1816D7AD",
    x"18169CCC",
    x"18166203",
    x"18162750",
    x"1815ECB4",
    x"1815B22F",
    x"181577C1",
    x"18153D69",
    x"18150329",
    x"1814C8FF",
    x"18148EEC",
    x"181454EF",
    x"18141B09",
    x"1813E13A",
    x"1813A781",
    x"18136DDF",
    x"18133453",
    x"1812FADE",
    x"1812C17F",
    x"18128837",
    x"18124F05",
    x"181215E9",
    x"1811DCE4",
    x"1811A3F5",
    x"18116B1C",
    x"18113259",
    x"1810F9AC",
    x"1810C116",
    x"18108896",
    x"1810502B",
    x"181017D7",
    x"180FDF99",
    x"180FA770",
    x"180F6F5E",
    x"180F3761",
    x"180EFF7A",
    x"180EC7AA",
    x"180E8FEE",
    x"180E5849",
    x"180E20B9",
    x"180DE940",
    x"180DB1DB",
    x"180D7A8D",
    x"180D4353",
    x"180D0C30",
    x"180CD522",
    x"180C9E29",
    x"180C6746",
    x"180C3079",
    x"180BF9C0",
    x"180BC31E",
    x"180B8C90",
    x"180B5618",
    x"180B1FB5",
    x"180AE967",
    x"180AB32E",
    x"180A7D0B",
    x"180A46FD",
    x"180A1104",
    x"1809DB1F",
    x"1809A550",
    x"18096F96",
    x"180939F1",
    x"18090461",
    x"1808CEE6",
    x"1808997F",
    x"1808642E",
    x"18082EF1",
    x"1807F9C9",
    x"1807C4B6",
    x"18078FB7",
    x"18075ACE",
    x"180725F8",
    x"1806F138",
    x"1806BC8C",
    x"180687F5",
    x"18065372",
    x"18061F03",
    x"1805EAAA",
    x"1805B664",
    x"18058233",
    x"18054E16",
    x"18051A0E",
    x"1804E61A",
    x"1804B23A",
    x"18047E6F",
    x"18044AB7",
    x"18041714",
    x"1803E385",
    x"1803B00B",
    x"18037CA4",
    x"18034951",
    x"18031613",
    x"1802E2E8",
    x"1802AFD1",
    x"18027CCF",
    x"180249E0",
    x"18021705",
    x"1801E43E",
    x"1801B18B",
    x"18017EEB",
    x"18014C5F",
    x"180119E7",
    x"1800E783",
    x"1800B533",
    x"180082F6",
    x"180050CC",
    x"18001EB6",
    x"17FFD968",
    x"17FF758B",
    x"17FF11D5",
    x"17FEAE45",
    x"17FE4ADC",
    x"17FDE79B",
    x"17FD847F",
    x"17FD218B",
    x"17FCBEBD",
    x"17FC5C16",
    x"17FBF995",
    x"17FB973B",
    x"17FB3507",
    x"17FAD2F9",
    x"17FA7112",
    x"17FA0F51",
    x"17F9ADB6",
    x"17F94C41",
    x"17F8EAF3",
    x"17F889CA",
    x"17F828C7",
    x"17F7C7EA",
    x"17F76733",
    x"17F706A1",
    x"17F6A636",
    x"17F645EF",
    x"17F5E5CF",
    x"17F585D4",
    x"17F525FE",
    x"17F4C64E",
    x"17F466C3",
    x"17F4075E",
    x"17F3A81E",
    x"17F34903",
    x"17F2EA0D",
    x"17F28B3C",
    x"17F22C90",
    x"17F1CE09",
    x"17F16FA7",
    x"17F1116A",
    x"17F0B351",
    x"17F0555D",
    x"17EFF78E",
    x"17EF99E4",
    x"17EF3C5E",
    x"17EEDEFD",
    x"17EE81C0",
    x"17EE24A7",
    x"17EDC7B3",
    x"17ED6AE3",
    x"17ED0E38",
    x"17ECB1B0",
    x"17EC554D",
    x"17EBF90E",
    x"17EB9CF2",
    x"17EB40FB",
    x"17EAE528",
    x"17EA8978",
    x"17EA2DEC",
    x"17E9D284",
    x"17E97740",
    x"17E91C1F",
    x"17E8C122",
    x"17E86648",
    x"17E80B92",
    x"17E7B0FF",
    x"17E7568F",
    x"17E6FC43",
    x"17E6A21A",
    x"17E64815",
    x"17E5EE32",
    x"17E59473",
    x"17E53AD6",
    x"17E4E15D",
    x"17E48806",
    x"17E42ED2",
    x"17E3D5C1",
    x"17E37CD3",
    x"17E32408",
    x"17E2CB5F",
    x"17E272D9",
    x"17E21A75",
    x"17E1C234",
    x"17E16A16",
    x"17E11219",
    x"17E0BA3F",
    x"17E06288",
    x"17E00AF2",
    x"17DFB37F",
    x"17DF5C2E",
    x"17DF04FF",
    x"17DEADF2",
    x"17DE5707",
    x"17DE003E",
    x"17DDA997",
    x"17DD5312",
    x"17DCFCAE",
    x"17DCA66C",
    x"17DC504C",
    x"17DBFA4E",
    x"17DBA471",
    x"17DB4EB5",
    x"17DAF91B",
    x"17DAA3A2",
    x"17DA4E4B",
    x"17D9F915",
    x"17D9A401",
    x"17D94F0D",
    x"17D8FA3B",
    x"17D8A58A",
    x"17D850F9",
    x"17D7FC8A",
    x"17D7A83C",
    x"17D7540F",
    x"17D70002",
    x"17D6AC17",
    x"17D6584C",
    x"17D604A2",
    x"17D5B118",
    x"17D55DB0",
    x"17D50A67",
    x"17D4B73F",
    x"17D46438",
    x"17D41151",
    x"17D3BE8A",
    x"17D36BE4",
    x"17D3195E",
    x"17D2C6F8",
    x"17D274B3",
    x"17D2228D",
    x"17D1D088",
    x"17D17EA2",
    x"17D12CDD",
    x"17D0DB37",
    x"17D089B1",
    x"17D0384C",
    x"17CFE705",
    x"17CF95DF",
    x"17CF44D8",
    x"17CEF3F1",
    x"17CEA32A",
    x"17CE5282",
    x"17CE01F9",
    x"17CDB190",
    x"17CD6147",
    x"17CD111C",
    x"17CCC111",
    x"17CC7125",
    x"17CC2159",
    x"17CBD1AB",
    x"17CB821D",
    x"17CB32AE",
    x"17CAE35D",
    x"17CA942C",
    x"17CA451A",
    x"17C9F626",
    x"17C9A751",
    x"17C9589B",
    x"17C90A04",
    x"17C8BB8B",
    x"17C86D31",
    x"17C81EF6",
    x"17C7D0D9",
    x"17C782DB",
    x"17C734FB",
    x"17C6E73A",
    x"17C69996",
    x"17C64C11",
    x"17C5FEAB",
    x"17C5B163",
    x"17C56438",
    x"17C5172C",
    x"17C4CA3E",
    x"17C47D6E",
    x"17C430BC",
    x"17C3E428",
    x"17C397B2",
    x"17C34B5A",
    x"17C2FF1F",
    x"17C2B302",
    x"17C26703",
    x"17C21B22",
    x"17C1CF5E",
    x"17C183B8",
    x"17C1382F",
    x"17C0ECC4",
    x"17C0A176",
    x"17C05646",
    x"17C00B33",
    x"17BFC03D",
    x"17BF7564",
    x"17BF2AA9",
    x"17BEE00B",
    x"17BE958A",
    x"17BE4B26",
    x"17BE00DF",
    x"17BDB6B6",
    x"17BD6CA9",
    x"17BD22B9",
    x"17BCD8E6",
    x"17BC8F2F",
    x"17BC4596",
    x"17BBFC19",
    x"17BBB2B9",
    x"17BB6975",
    x"17BB204E",
    x"17BAD744",
    x"17BA8E56",
    x"17BA4585",
    x"17B9FCD0",
    x"17B9B437",
    x"17B96BBB",
    x"17B9235B",
    x"17B8DB17",
    x"17B892F0",
    x"17B84AE4",
    x"17B802F5",
    x"17B7BB22",
    x"17B7736B",
    x"17B72BD0",
    x"17B6E451",
    x"17B69CEE",
    x"17B655A6",
    x"17B60E7B",
    x"17B5C76B",
    x"17B58077",
    x"17B5399F",
    x"17B4F2E2",
    x"17B4AC41",
    x"17B465BB",
    x"17B41F51",
    x"17B3D903",
    x"17B392D0",
    x"17B34CB8",
    x"17B306BC",
    x"17B2C0DB",
    x"17B27B15",
    x"17B2356B",
    x"17B1EFDB",
    x"17B1AA67",
    x"17B1650E",
    x"17B11FD0",
    x"17B0DAAD",
    x"17B095A5",
    x"17B050B8",
    x"17B00BE6",
    x"17AFC72F",
    x"17AF8293",
    x"17AF3E11",
    x"17AEF9AA",
    x"17AEB55E",
    x"17AE712C",
    x"17AE2D16",
    x"17ADE919",
    x"17ADA537",
    x"17AD6170",
    x"17AD1DC3",
    x"17ACDA31",
    x"17AC96B9",
    x"17AC535B",
    x"17AC1018",
    x"17ABCCEF",
    x"17AB89E0",
    x"17AB46EB",
    x"17AB0410",
    x"17AAC150",
    x"17AA7EA9",
    x"17AA3C1D",
    x"17A9F9AA",
    x"17A9B752",
    x"17A97513",
    x"17A932EE",
    x"17A8F0E3",
    x"17A8AEF2",
    x"17A86D1A",
    x"17A82B5D",
    x"17A7E9B9",
    x"17A7A82E",
    x"17A766BD",
    x"17A72566",
    x"17A6E428",
    x"17A6A304",
    x"17A661F9",
    x"17A62107",
    x"17A5E02F",
    x"17A59F70",
    x"17A55ECA",
    x"17A51E3E",
    x"17A4DDCB",
    x"17A49D70",
    x"17A45D30",
    x"17A41D08",
    x"17A3DCF9",
    x"17A39D03",
    x"17A35D26",
    x"17A31D62",
    x"17A2DDB7",
    x"17A29E25",
    x"17A25EAC",
    x"17A21F4B",
    x"17A1E003",
    x"17A1A0D4",
    x"17A161BD",
    x"17A122C0",
    x"17A0E3DA",
    x"17A0A50E",
    x"17A06659",
    x"17A027BE",
    x"179FE93A",
    x"179FAACF",
    x"179F6C7D",
    x"179F2E43",
    x"179EF021",
    x"179EB217",
    x"179E7426",
    x"179E364C",
    x"179DF88B",
    x"179DBAE2",
    x"179D7D51",
    x"179D3FD8",
    x"179D0277",
    x"179CC52E",
    x"179C87FD",
    x"179C4AE4",
    x"179C0DE3",
    x"179BD0F9",
    x"179B9427",
    x"179B576D",
    x"179B1ACB",
    x"179ADE40",
    x"179AA1CD",
    x"179A6572",
    x"179A292E",
    x"1799ED02",
    x"1799B0ED",
    x"179974F0",
    x"1799390A",
    x"1798FD3B",
    x"1798C184",
    x"179885E4",
    x"17984A5B",
    x"17980EEA",
    x"1797D38F",
    x"1797984C",
    x"17975D20",
    x"1797220C",
    x"1796E70E",
    x"1796AC27",
    x"17967157",
    x"1796369F",
    x"1795FBFD",
    x"1795C172",
    x"179586FE",
    x"17954CA0",
    x"1795125A",
    x"1794D82A",
    x"17949E11",
    x"1794640E",
    x"17942A23",
    x"1793F04D",
    x"1793B68F",
    x"17937CE7",
    x"17934355",
    x"179309DA",
    x"1792D076",
    x"17929727",
    x"17925DEF",
    x"179224CE",
    x"1791EBC3",
    x"1791B2CE",
    x"179179EF",
    x"17914126",
    x"17910874",
    x"1790CFD8",
    x"17909752",
    x"17905EE2",
    x"17902688",
    x"178FEE43",
    x"178FB615",
    x"178F7DFD",
    x"178F45FB",
    x"178F0E0F",
    x"178ED638",
    x"178E9E77",
    x"178E66CC",
    x"178E2F37",
    x"178DF7B7",
    x"178DC04D",
    x"178D88F9",
    x"178D51BA",
    x"178D1A91",
    x"178CE37E",
    x"178CAC7F",
    x"178C7597",
    x"178C3EC4",
    x"178C0806",
    x"178BD15D",
    x"178B9ACA",
    x"178B644C",
    x"178B2DE4",
    x"178AF790",
    x"178AC152",
    x"178A8B29",
    x"178A5516",
    x"178A1F17",
    x"1789E92D",
    x"1789B359",
    x"17897D99",
    x"178947EF",
    x"17891259",
    x"1788DCD8",
    x"1788A76C",
    x"17887215",
    x"17883CD3",
    x"178807A6",
    x"1787D28D",
    x"17879D89",
    x"1787689A",
    x"178733C0",
    x"1786FEFA",
    x"1786CA48",
    x"178695AC",
    x"17866124",
    x"17862CB0",
    x"1785F851",
    x"1785C406",
    x"17858FCF",
    x"17855BAD",
    x"178527A0",
    x"1784F3A6",
    x"1784BFC1",
    x"17848BF1",
    x"17845834",
    x"1784248C",
    x"1783F0F8",
    x"1783BD77",
    x"17838A0C",
    x"178356B4",
    x"17832370",
    x"1782F040",
    x"1782BD24",
    x"17828A1C",
    x"17825728",
    x"17822448",
    x"1781F17C",
    x"1781BEC3",
    x"17818C1F",
    x"1781598E",
    x"17812711",
    x"1780F4A7",
    x"1780C252",
    x"17809010",
    x"17805DE1",
    x"17802BC6",
    x"177FF37E",
    x"177F8F96",
    x"177F2BD6",
    x"177EC83C",
    x"177E64C9",
    x"177E017D",
    x"177D9E58",
    x"177D3B59",
    x"177CD882",
    x"177C75D0",
    x"177C1345",
    x"177BB0E1",
    x"177B4EA3",
    x"177AEC8C",
    x"177A8A9A",
    x"177A28CF",
    x"1779C72B",
    x"177965AC",
    x"17790453",
    x"1778A320",
    x"17784214",
    x"1777E12D",
    x"1777806C",
    x"17771FD0",
    x"1776BF5B",
    x"17765F0B",
    x"1775FEE1",
    x"17759EDC",
    x"17753EFC",
    x"1774DF43",
    x"17747FAE",
    x"1774203F",
    x"1773C0F5",
    x"177361D0",
    x"177302D0",
    x"1772A3F6",
    x"17724540",
    x"1771E6B0",
    x"17718844",
    x"177129FD",
    x"1770CBDB",
    x"17706DDE",
    x"17701005",
    x"176FB251",
    x"176F54C2",
    x"176EF757",
    x"176E9A11",
    x"176E3CEF",
    x"176DDFF1",
    x"176D8318",
    x"176D2663",
    x"176CC9D2",
    x"176C6D65",
    x"176C111C",
    x"176BB4F8",
    x"176B58F7",
    x"176AFD1A",
    x"176AA161",
    x"176A45CC",
    x"1769EA5B",
    x"17698F0D",
    x"176933E3",
    x"1768D8DC",
    x"17687DF9",
    x"1768233A",
    x"1767C89E",
    x"17676E25",
    x"176713D0",
    x"1766B99E",
    x"17665F8F",
    x"176605A3",
    x"1765ABDA",
    x"17655235",
    x"1764F8B2",
    x"17649F52",
    x"17644616",
    x"1763ECFC",
    x"17639404",
    x"17633B30",
    x"1762E27E",
    x"176289EF",
    x"17623182",
    x"1761D938",
    x"17618111",
    x"1761290B",
    x"1760D129",
    x"17607968",
    x"176021CA",
    x"175FCA4E",
    x"175F72F4",
    x"175F1BBC",
    x"175EC4A6",
    x"175E6DB2",
    x"175E16E0",
    x"175DC030",
    x"175D69A2",
    x"175D1336",
    x"175CBCEB",
    x"175C66C2",
    x"175C10BB",
    x"175BBAD5",
    x"175B6511",
    x"175B0F6E",
    x"175AB9ED",
    x"175A648D",
    x"175A0F4E",
    x"1759BA31",
    x"17596535",
    x"1759105A",
    x"1758BBA0",
    x"17586707",
    x"1758128F",
    x"1757BE39",
    x"17576A03",
    x"175715EE",
    x"1756C1FA",
    x"17566E26",
    x"17561A74",
    x"1755C6E1",
    x"17557370",
    x"1755201F",
    x"1754CCEF",
    x"175479DF",
    x"175426F0",
    x"1753D421",
    x"17538172",
    x"17532EE4",
    x"1752DC75",
    x"17528A27",
    x"175237F9",
    x"1751E5EC",
    x"175193FE",
    x"17514230",
    x"1750F082",
    x"17509EF4",
    x"17504D86",
    x"174FFC37",
    x"174FAB09",
    x"174F59FA",
    x"174F090A",
    x"174EB83B",
    x"174E678B",
    x"174E16FA",
    x"174DC689",
    x"174D7637",
    x"174D2604",
    x"174CD5F1",
    x"174C85FD",
    x"174C3628",
    x"174BE673",
    x"174B96DC",
    x"174B4765",
    x"174AF80C",
    x"174AA8D3",
    x"174A59B9",
    x"174A0ABD",
    x"1749BBE0",
    x"17496D22",
    x"17491E83",
    x"1748D002",
    x"174881A0",
    x"1748335D",
    x"1747E538",
    x"17479732",
    x"1747494A",
    x"1746FB81",
    x"1746ADD6",
    x"17466049",
    x"174612DA",
    x"1745C58A",
    x"17457858",
    x"17452B44",
    x"1744DE4E",
    x"17449176",
    x"174444BD",
    x"1743F821",
    x"1743ABA3",
    x"17435F43",
    x"17431300",
    x"1742C6DC",
    x"17427AD5",
    x"17422EEC",
    x"1741E320",
    x"17419772",
    x"17414BE2",
    x"1741006F",
    x"1740B519",
    x"174069E1",
    x"17401EC7",
    x"173FD3C9",
    x"173F88E9",
    x"173F3E26",
    x"173EF381",
    x"173EA8F8",
    x"173E5E8D",
    x"173E143E",
    x"173DCA0D",
    x"173D7FF8",
    x"173D3601",
    x"173CEC26",
    x"173CA268",
    x"173C58C7",
    x"173C0F43",
    x"173BC5DB",
    x"173B7C90",
    x"173B3362",
    x"173AEA50",
    x"173AA15B",
    x"173A5882",
    x"173A0FC6",
    x"1739C726",
    x"17397EA2",
    x"1739363B",
    x"1738EDF0",
    x"1738A5C1",
    x"17385DAE",
    x"173815B8",
    x"1737CDDD",
    x"1737861F",
    x"17373E7D",
    x"1736F6F6",
    x"1736AF8C",
    x"1736683D",
    x"1736210A",
    x"1735D9F3",
    x"173592F8",
    x"17354C18",
    x"17350554",
    x"1734BEAC",
    x"1734781F",
    x"173431AE",
    x"1733EB59",
    x"1733A51E",
    x"17335F00",
    x"173318FC",
    x"1732D314",
    x"17328D47",
    x"17324796",
    x"173201FF",
    x"1731BC84",
    x"17317724",
    x"173131DF",
    x"1730ECB5",
    x"1730A7A6",
    x"173062B2",
    x"17301DD9",
    x"172FD91B",
    x"172F9477",
    x"172F4FEF",
    x"172F0B81",
    x"172EC72E",
    x"172E82F5",
    x"172E3ED7",
    x"172DFAD4",
    x"172DB6EB",
    x"172D731D",
    x"172D2F69",
    x"172CEBD0",
    x"172CA851",
    x"172C64ED",
    x"172C21A2",
    x"172BDE72",
    x"172B9B5D",
    x"172B5861",
    x"172B157F",
    x"172AD2B8",
    x"172A900B",
    x"172A4D78",
    x"172A0AFE",
    x"1729C89F",
    x"1729865A",
    x"1729442E",
    x"1729021C",
    x"1728C024",
    x"17287E46",
    x"17283C82",
    x"1727FAD7",
    x"1727B946",
    x"172777CE",
    x"17273670",
    x"1726F52C",
    x"1726B401",
    x"172672EF",
    x"172631F7",
    x"1725F118",
    x"1725B052",
    x"17256FA6",
    x"17252F13",
    x"1724EE99",
    x"1724AE39",
    x"17246DF1",
    x"17242DC3",
    x"1723EDAD",
    x"1723ADB1",
    x"17236DCE",
    x"17232E03",
    x"1722EE52",
    x"1722AEB9",
    x"17226F39",
    x"17222FD2",
    x"1721F084",
    x"1721B14E",
    x"17217231",
    x"1721332D",
    x"1720F441",
    x"1720B56E",
    x"172076B4",
    x"17203811",
    x"171FF988",
    x"171FBB17",
    x"171F7CBE",
    x"171F3E7D",
    x"171F0055",
    x"171EC245",
    x"171E844D",
    x"171E466D",
    x"171E08A6",
    x"171DCAF7",
    x"171D8D5F",
    x"171D4FE0",
    x"171D1279",
    x"171CD52A",
    x"171C97F2",
    x"171C5AD3",
    x"171C1DCB",
    x"171BE0DC",
    x"171BA404",
    x"171B6744",
    x"171B2A9B",
    x"171AEE0A",
    x"171AB191",
    x"171A7530",
    x"171A38E6",
    x"1719FCB3",
    x"1719C098",
    x"17198495",
    x"171948A9",
    x"17190CD4",
    x"1718D116",
    x"17189570",
    x"171859E2",
    x"17181E6A",
    x"1717E30A",
    x"1717A7C1",
    x"17176C8F",
    x"17173174",
    x"1716F670",
    x"1716BB83",
    x"171680AE",
    x"171645EF",
    x"17160B47",
    x"1715D0B6",
    x"1715963C",
    x"17155BD9",
    x"1715218C",
    x"1714E757",
    x"1714AD38",
    x"1714732F",
    x"1714393E",
    x"1713FF62",
    x"1713C59E",
    x"17138BF0",
    x"17135259",
    x"171318D8",
    x"1712DF6D",
    x"1712A619",
    x"17126CDB",
    x"171233B4",
    x"1711FAA3",
    x"1711C1A8",
    x"171188C4",
    x"17114FF5",
    x"1711173D",
    x"1710DE9B",
    x"1710A60F",
    x"17106D99",
    x"1710353A",
    x"170FFCF0",
    x"170FC4BC",
    x"170F8C9E",
    x"170F5496",
    x"170F1CA4",
    x"170EE4C8",
    x"170EAD01",
    x"170E7551",
    x"170E3DB6",
    x"170E0630",
    x"170DCEC1",
    x"170D9767",
    x"170D6023",
    x"170D28F4",
    x"170CF1DB",
    x"170CBAD7",
    x"170C83E9",
    x"170C4D10",
    x"170C164C",
    x"170BDF9E",
    x"170BA906",
    x"170B7282",
    x"170B3C14",
    x"170B05BB",
    x"170ACF78",
    x"170A9949",
    x"170A6330",
    x"170A2D2C",
    x"1709F73D",
    x"1709C163",
    x"17098B9E",
    x"170955ED",
    x"17092052",
    x"1708EACC",
    x"1708B55B",
    x"17087FFF",
    x"17084AB7",
    x"17081584",
    x"1707E066",
    x"1707AB5D",
    x"17077668",
    x"17074188",
    x"17070CBD",
    x"1706D806",
    x"1706A364",
    x"17066ED7",
    x"17063A5E",
    x"170605F9",
    x"1705D1A9",
    x"17059D6D",
    x"17056946",
    x"17053533",
    x"17050134",
    x"1704CD4A",
    x"17049974",
    x"170465B2",
    x"17043205",
    x"1703FE6B",
    x"1703CAE6",
    x"17039775",
    x"17036417",
    x"170330CE",
    x"1702FD99",
    x"1702CA78",
    x"1702976B",
    x"17026472",
    x"1702318D",
    x"1701FEBB",
    x"1701CBFE",
    x"17019954",
    x"170166BE",
    x"1701343C",
    x"170101CD",
    x"1700CF72",
    x"17009D2B",
    x"17006AF7",
    x"170038D7",
    x"170006CB",
    x"16FFA9A4",
    x"16FF45D9",
    x"16FEE235",
    x"16FE7EB8",
    x"16FE1B62",
    x"16FDB833",
    x"16FD552A",
    x"16FCF249",
    x"16FC8F8D",
    x"16FC2CF8",
    x"16FBCA8A",
    x"16FB6842",
    x"16FB0621",
    x"16FAA425",
    x"16FA4250",
    x"16F9E0A1",
    x"16F97F19",
    x"16F91DB6",
    x"16F8BC7A",
    x"16F85B63",
    x"16F7FA72",
    x"16F799A7",
    x"16F73902",
    x"16F6D883",
    x"16F67829",
    x"16F617F5",
    x"16F5B7E6",
    x"16F557FD",
    x"16F4F839",
    x"16F4989B",
    x"16F43922",
    x"16F3D9CE",
    x"16F37AA0",
    x"16F31B97",
    x"16F2BCB2",
    x"16F25DF3",
    x"16F1FF59",
    x"16F1A0E4",
    x"16F14293",
    x"16F0E468",
    x"16F08661",
    x"16F0287F",
    x"16EFCAC1",
    x"16EF6D28",
    x"16EF0FB4",
    x"16EEB264",
    x"16EE5538",
    x"16EDF831",
    x"16ED9B4F",
    x"16ED3E90",
    x"16ECE1F6",
    x"16EC857F",
    x"16EC292D",
    x"16EBCCFF",
    x"16EB70F5",
    x"16EB150F",
    x"16EAB94D",
    x"16EA5DAE",
    x"16EA0233",
    x"16E9A6DC",
    x"16E94BA9",
    x"16E8F099",
    x"16E895AD",
    x"16E83AE4",
    x"16E7E03F",
    x"16E785BD",
    x"16E72B5F",
    x"16E6D123",
    x"16E6770B",
    x"16E61D16",
    x"16E5C344",
    x"16E56996",
    x"16E5100A",
    x"16E4B6A1",
    x"16E45D5B",
    x"16E40438",
    x"16E3AB38",
    x"16E3525A",
    x"16E2F9A0",
    x"16E2A107",
    x"16E24892",
    x"16E1F03F",
    x"16E1980E",
    x"16E14000",
    x"16E0E814",
    x"16E0904B",
    x"16E038A3",
    x"16DFE11E",
    x"16DF89BB",
    x"16DF327B",
    x"16DEDB5C",
    x"16DE845F",
    x"16DE2D85",
    x"16DDD6CC",
    x"16DD8035",
    x"16DD29BF",
    x"16DCD36C",
    x"16DC7D3A",
    x"16DC272A",
    x"16DBD13C",
    x"16DB7B6F",
    x"16DB25C3",
    x"16DAD039",
    x"16DA7AD1",
    x"16DA2589",
    x"16D9D063",
    x"16D97B5E",
    x"16D9267B",
    x"16D8D1B8",
    x"16D87D17",
    x"16D82897",
    x"16D7D437",
    x"16D77FF9",
    x"16D72BDB",
    x"16D6D7DE",
    x"16D68403",
    x"16D63047",
    x"16D5DCAD",
    x"16D58933",
    x"16D535DA",
    x"16D4E2A1",
    x"16D48F89",
    x"16D43C91",
    x"16D3E9B9",
    x"16D39702",
    x"16D3446B",
    x"16D2F1F5",
    x"16D29F9E",
    x"16D24D68",
    x"16D1FB52",
    x"16D1A95C",
    x"16D15785",
    x"16D105CF",
    x"16D0B439",
    x"16D062C2",
    x"16D0116C",
    x"16CFC035",
    x"16CF6F1D",
    x"16CF1E26",
    x"16CECD4E",
    x"16CE7C95",
    x"16CE2BFD",
    x"16CDDB83",
    x"16CD8B29",
    x"16CD3AEE",
    x"16CCEAD3",
    x"16CC9AD7",
    x"16CC4AFA",
    x"16CBFB3C",
    x"16CBAB9E",
    x"16CB5C1E",
    x"16CB0CBE",
    x"16CABD7C",
    x"16CA6E5A",
    x"16CA1F56",
    x"16C9D071",
    x"16C981AB",
    x"16C93304",
    x"16C8E47B",
    x"16C89611",
    x"16C847C6",
    x"16C7F999",
    x"16C7AB8B",
    x"16C75D9B",
    x"16C70FCA",
    x"16C6C217",
    x"16C67482",
    x"16C6270C",
    x"16C5D9B4",
    x"16C58C7A",
    x"16C53F5E",
    x"16C4F260",
    x"16C4A581",
    x"16C458BF",
    x"16C40C1B",
    x"16C3BF95",
    x"16C3732E",
    x"16C326E3",
    x"16C2DAB7",
    x"16C28EA9",
    x"16C242B8",
    x"16C1F6E4",
    x"16C1AB2F",
    x"16C15F97",
    x"16C1141C",
    x"16C0C8BF",
    x"16C07D7F",
    x"16C0325D",
    x"16BFE758",
    x"16BF9C70",
    x"16BF51A6",
    x"16BF06F8",
    x"16BEBC68",
    x"16BE71F5",
    x"16BE279F",
    x"16BDDD66",
    x"16BD934A",
    x"16BD494B",
    x"16BCFF69",
    x"16BCB5A3",
    x"16BC6BFB",
    x"16BC226F",
    x"16BBD900",
    x"16BB8FAE",
    x"16BB4678",
    x"16BAFD5F",
    x"16BAB462",
    x"16BA6B82",
    x"16BA22BE",
    x"16B9DA16",
    x"16B9918B",
    x"16B9491D",
    x"16B900CA",
    x"16B8B894",
    x"16B8707A",
    x"16B8287C",
    x"16B7E09A",
    x"16B798D5",
    x"16B7512B",
    x"16B7099D",
    x"16B6C22B",
    x"16B67AD6",
    x"16B6339B",
    x"16B5EC7D",
    x"16B5A57B",
    x"16B55E94",
    x"16B517C9",
    x"16B4D119",
    x"16B48A85",
    x"16B4440D",
    x"16B3FDB0",
    x"16B3B76F",
    x"16B37149",
    x"16B32B3E",
    x"16B2E54F",
    x"16B29F7B",
    x"16B259C3",
    x"16B21425",
    x"16B1CEA3",
    x"16B1893C",
    x"16B143F0",
    x"16B0FEBF",
    x"16B0B9A9",
    x"16B074AD",
    x"16B02FCD",
    x"16AFEB08",
    x"16AFA65E",
    x"16AF61CE",
    x"16AF1D59",
    x"16AED8FF",
    x"16AE94C0",
    x"16AE509B",
    x"16AE0C91",
    x"16ADC8A1",
    x"16AD84CC",
    x"16AD4111",
    x"16ACFD71",
    x"16ACB9EB",
    x"16AC7680",
    x"16AC332F",
    x"16ABEFF8",
    x"16ABACDB",
    x"16AB69D9",
    x"16AB26F1",
    x"16AAE422",
    x"16AAA16E",
    x"16AA5ED4",
    x"16AA1C54",
    x"16A9D9EE",
    x"16A997A2",
    x"16A95570",
    x"16A91357",
    x"16A8D159",
    x"16A88F74",
    x"16A84DA8",
    x"16A80BF7",
    x"16A7CA5F",
    x"16A788E1",
    x"16A7477C",
    x"16A70631",
    x"16A6C4FF",
    x"16A683E7",
    x"16A642E8",
    x"16A60203",
    x"16A5C137",
    x"16A58084",
    x"16A53FEA",
    x"16A4FF6A",
    x"16A4BF03",
    x"16A47EB5",
    x"16A43E80",
    x"16A3FE64",
    x"16A3BE61",
    x"16A37E77",
    x"16A33EA6",
    x"16A2FEEE",
    x"16A2BF4F",
    x"16A27FC9",
    x"16A2405B",
    x"16A20106",
    x"16A1C1CA",
    x"16A182A7",
    x"16A1439C",
    x"16A104AA",
    x"16A0C5D1",
    x"16A08710",
    x"16A04867",
    x"16A009D7",
    x"169FCB5F",
    x"169F8D00",
    x"169F4EB9",
    x"169F108B",
    x"169ED274",
    x"169E9476",
    x"169E5690",
    x"169E18C2",
    x"169DDB0D",
    x"169D9D6F",
    x"169D5FEA",
    x"169D227C",
    x"169CE527",
    x"169CA7E9",
    x"169C6AC4",
    x"169C2DB6",
    x"169BF0C0",
    x"169BB3E2",
    x"169B771B",
    x"169B3A6D",
    x"169AFDD6",
    x"169AC156",
    x"169A84EF",
    x"169A489F",
    x"169A0C66",
    x"1699D045",
    x"1699943B",
    x"16995849",
    x"16991C6E",
    x"1698E0AB",
    x"1698A4FF",
    x"1698696A",
    x"16982DEC",
    x"1697F286",
    x"1697B737",
    x"16977BFF",
    x"169740DE",
    x"169705D4",
    x"1696CAE1",
    x"16969006",
    x"16965541",
    x"16961A93",
    x"1695DFFC",
    x"1695A57C",
    x"16956B13",
    x"169530C0",
    x"1694F685",
    x"1694BC60",
    x"16948252",
    x"1694485A",
    x"16940E79",
    x"1693D4AF",
    x"16939AFB",
    x"1693615E",
    x"169327D7",
    x"1692EE66",
    x"1692B50D",
    x"16927BC9",
    x"1692429C",
    x"16920985",
    x"1691D084",
    x"1691979A",
    x"16915EC6",
    x"16912608",
    x"1690ED60",
    x"1690B4CE",
    x"16907C53",
    x"169043ED",
    x"16900B9E",
    x"168FD364",
    x"168F9B41",
    x"168F6333",
    x"168F2B3B",
    x"168EF359",
    x"168EBB8D",
    x"168E83D7",
    x"168E4C36",
    x"168E14AB",
    x"168DDD36",
    x"168DA5D6",
    x"168D6E8C",
    x"168D3758",
    x"168D0039",
    x"168CC930",
    x"168C923C",
    x"168C5B5D",
    x"168C2494",
    x"168BEDE1",
    x"168BB743",
    x"168B80BA",
    x"168B4A46",
    x"168B13E8",
    x"168ADD9E",
    x"168AA76A",
    x"168A714C",
    x"168A3B42",
    x"168A054D",
    x"1689CF6E",
    x"168999A3",
    x"168963EE",
    x"16892E4D",
    x"1688F8C2",
    x"1688C34B",
    x"16888DE9",
    x"1688589C",
    x"16882364",
    x"1687EE40",
    x"1687B932",
    x"16878438",
    x"16874F52",
    x"16871A82",
    x"1686E5C6",
    x"1686B11E",
    x"16867C8B",
    x"1686480D",
    x"168613A3",
    x"1685DF4D",
    x"1685AB0C",
    x"168576E0",
    x"168542C8",
    x"16850EC4",
    x"1684DAD4",
    x"1684A6F9",
    x"16847332",
    x"16843F7F",
    x"16840BE0",
    x"1683D855",
    x"1683A4DF",
    x"1683717D",
    x"16833E2E",
    x"16830AF4",
    x"1682D7CE",
    x"1682A4BB",
    x"168271BD",
    x"16823ED2",
    x"16820BFC",
    x"1681D939",
    x"1681A68A",
    x"168173EF",
    x"16814168",
    x"16810EF4",
    x"1680DC94",
    x"1680AA48",
    x"1680780F",
    x"168045EA",
    x"168013D8",
    x"167FC3B4",
    x"167F5FE0",
    x"167EFC32",
    x"167E98AA",
    x"167E354A",
    x"167DD211",
    x"167D6EFE",
    x"167D0C12",
    x"167CA94D",
    x"167C46AE",
    x"167BE435",
    x"167B81E4",
    x"167B1FB8",
    x"167ABDB3",
    x"167A5BD4",
    x"1679FA1B",
    x"16799888",
    x"1679371C",
    x"1678D5D5",
    x"167874B5",
    x"167813BA",
    x"1677B2E5",
    x"16775236",
    x"1676F1AD",
    x"16769149",
    x"1676310B",
    x"1675D0F3",
    x"16757100",
    x"16751133",
    x"1674B18B",
    x"16745208",
    x"1673F2AB",
    x"16739372",
    x"1673345F",
    x"1672D572",
    x"167276A9",
    x"16721805",
    x"1671B986",
    x"16715B2C",
    x"1670FCF7",
    x"16709EE6",
    x"167040FA",
    x"166FE333",
    x"166F8591",
    x"166F2813",
    x"166ECABA",
    x"166E6D85",
    x"166E1074",
    x"166DB388",
    x"166D56C0",
    x"166CFA1C",
    x"166C9D9C",
    x"166C4141",
    x"166BE509",
    x"166B88F6",
    x"166B2D06",
    x"166AD13B",
    x"166A7593",
    x"166A1A0F",
    x"1669BEAF",
    x"16696372",
    x"16690859",
    x"1668AD63",
    x"16685291",
    x"1667F7E3",
    x"16679D58",
    x"166742F0",
    x"1666E8AB",
    x"16668E8A",
    x"1666348C",
    x"1665DAB1",
    x"166580F9",
    x"16652764",
    x"1664CDF2",
    x"166474A3",
    x"16641B77",
    x"1663C26E",
    x"16636987",
    x"166310C3",
    x"1662B822",
    x"16625FA3",
    x"16620747",
    x"1661AF0E",
    x"166156F7",
    x"1660FF02",
    x"1660A72F",
    x"16604F7F",
    x"165FF7F1",
    x"165FA085",
    x"165F493C",
    x"165EF214",
    x"165E9B0F",
    x"165E442B",
    x"165DED69",
    x"165D96CA",
    x"165D404C",
    x"165CE9EF",
    x"165C93B5",
    x"165C3D9C",
    x"165BE7A5",
    x"165B91CF",
    x"165B3C1B",
    x"165AE688",
    x"165A9117",
    x"165A3BC7",
    x"1659E698",
    x"1659918A",
    x"16593C9E",
    x"1658E7D3",
    x"16589329",
    x"16583EA0",
    x"1657EA38",
    x"165795F1",
    x"165741CB",
    x"1656EDC6",
    x"165699E1",
    x"1656461D",
    x"1655F27A",
    x"16559EF8",
    x"16554B96",
    x"1654F855",
    x"1654A534",
    x"16545234",
    x"1653FF54",
    x"1653AC94",
    x"165359F5",
    x"16530776",
    x"1652B517",
    x"165262D9",
    x"165210BA",
    x"1651BEBB",
    x"16516CDD",
    x"16511B1E",
    x"1650C980",
    x"16507801",
    x"165026A2",
    x"164FD563",
    x"164F8443",
    x"164F3343",
    x"164EE263",
    x"164E91A3",
    x"164E4101",
    x"164DF080",
    x"164DA01D",
    x"164D4FDB",
    x"164CFFB7",
    x"164CAFB3",
    x"164C5FCE",
    x"164C1008",
    x"164BC061",
    x"164B70DA",
    x"164B2171",
    x"164AD228",
    x"164A82FD",
    x"164A33F1",
    x"1649E504",
    x"16499636",
    x"16494787",
    x"1648F8F6",
    x"1648AA84",
    x"16485C31",
    x"16480DFC",
    x"1647BFE6",
    x"164771EE",
    x"16472415",
    x"1646D65A",
    x"164688BE",
    x"16463B3F",
    x"1645EDDF",
    x"1645A09E",
    x"1645537A",
    x"16450674",
    x"1644B98D",
    x"16446CC3",
    x"16442018",
    x"1643D38A",
    x"1643871B",
    x"16433AC9",
    x"1642EE95",
    x"1642A27E",
    x"16425686",
    x"16420AAB",
    x"1641BEED",
    x"1641734D",
    x"164127CB",
    x"1640DC66",
    x"1640911F",
    x"164045F5",
    x"163FFAE8",
    x"163FAFF9",
    x"163F6527",
    x"163F1A72",
    x"163ECFDA",
    x"163E855F",
    x"163E3B02",
    x"163DF0C1",
    x"163DA69E",
    x"163D5C97",
    x"163D12AD",
    x"163CC8E1",
    x"163C7F31",
    x"163C359D",
    x"163BEC27",
    x"163BA2CD",
    x"163B598F",
    x"163B106F",
    x"163AC76B",
    x"163A7E83",
    x"163A35B8",
    x"1639ED09",
    x"1639A477",
    x"16395C00",
    x"163913A7",
    x"1638CB69",
    x"16388348",
    x"16383B42",
    x"1637F359",
    x"1637AB8C",
    x"163763DB",
    x"16371C46",
    x"1636D4CD",
    x"16368D70",
    x"1636462F",
    x"1635FF09",
    x"1635B7FF",
    x"16357111",
    x"16352A3F",
    x"1634E388",
    x"16349CED",
    x"1634566E",
    x"1634100A",
    x"1633C9C1",
    x"16338394",
    x"16333D82",
    x"1632F78C",
    x"1632B1B1",
    x"16326BF1",
    x"1632264D",
    x"1631E0C3",
    x"16319B55",
    x"16315602",
    x"163110CA",
    x"1630CBAD",
    x"163086AB",
    x"163041C4",
    x"162FFCF7",
    x"162FB846",
    x"162F73AF",
    x"162F2F34",
    x"162EEAD3",
    x"162EA68C",
    x"162E6260",
    x"162E1E4F",
    x"162DDA59",
    x"162D967D",
    x"162D52BB",
    x"162D0F14",
    x"162CCB87",
    x"162C8815",
    x"162C44BD",
    x"162C017F",
    x"162BBE5C",
    x"162B7B53",
    x"162B3863",
    x"162AF58E",
    x"162AB2D4",
    x"162A7033",
    x"162A2DAC",
    x"1629EB3F",
    x"1629A8EC",
    x"162966B3",
    x"16292494",
    x"1628E28E",
    x"1628A0A3",
    x"16285ED1",
    x"16281D19",
    x"1627DB7A",
    x"162799F5",
    x"1627588A",
    x"16271738",
    x"1626D600",
    x"162694E1",
    x"162653DB",
    x"162612EF",
    x"1625D21D",
    x"16259163",
    x"162550C3",
    x"1625103C",
    x"1624CFCE",
    x"16248F7A",
    x"16244F3E",
    x"16240F1C",
    x"1623CF12",
    x"16238F22",
    x"16234F4B",
    x"16230F8C",
    x"1622CFE6",
    x"1622905A",
    x"162250E6",
    x"1622118A",
    x"1621D248",
    x"1621931E",
    x"1621540D",
    x"16211514",
    x"1620D635",
    x"1620976D",
    x"162058BE",
    x"16201A28",
    x"161FDBAA",
    x"161F9D44",
    x"161F5EF7",
    x"161F20C2",
    x"161EE2A5",
    x"161EA4A1",
    x"161E66B5",
    x"161E28E1",
    x"161DEB25",
    x"161DAD81",
    x"161D6FF5",
    x"161D3281",
    x"161CF526",
    x"161CB7E2",
    x"161C7AB6",
    x"161C3DA2",
    x"161C00A6",
    x"161BC3C1",
    x"161B86F5",
    x"161B4A40",
    x"161B0DA3",
    x"161AD11D",
    x"161A94AF",
    x"161A5859",
    x"161A1C1A",
    x"1619DFF3",
    x"1619A3E3",
    x"161967EB",
    x"16192C0A",
    x"1618F041",
    x"1618B48F",
    x"161878F4",
    x"16183D70",
    x"16180204",
    x"1617C6AE",
    x"16178B70",
    x"1617504A",
    x"1617153A",
    x"1616DA41",
    x"16169F5F",
    x"16166494",
    x"161629E1",
    x"1615EF44",
    x"1615B4BE",
    x"16157A4E",
    x"16153FF6",
    x"161505B4",
    x"1614CB8A",
    x"16149175",
    x"16145778",
    x"16141D91",
    x"1613E3C1",
    x"1613AA07",
    x"16137064",
    x"161336D7",
    x"1612FD61",
    x"1612C401",
    x"16128AB8",
    x"16125185",
    x"16121868",
    x"1611DF62",
    x"1611A672",
    x"16116D98",
    x"161134D4",
    x"1610FC27",
    x"1610C38F",
    x"16108B0E",
    x"161052A3",
    x"16101A4D",
    x"160FE20E",
    x"160FA9E5",
    x"160F71D1",
    x"160F39D4",
    x"160F01EC",
    x"160ECA1A",
    x"160E925E",
    x"160E5AB8",
    x"160E2327",
    x"160DEBAC",
    x"160DB447",
    x"160D7CF7",
    x"160D45BD",
    x"160D0E99",
    x"160CD78A",
    x"160CA091",
    x"160C69AD",
    x"160C32DE",
    x"160BFC25",
    x"160BC581",
    x"160B8EF3",
    x"160B5879",
    x"160B2215",
    x"160AEBC7",
    x"160AB58D",
    x"160A7F69",
    x"160A495A",
    x"160A1360",
    x"1609DD7A",
    x"1609A7AA",
    x"160971EF",
    x"16093C49",
    x"160906B8",
    x"1608D13C",
    x"16089BD5",
    x"16086682",
    x"16083145",
    x"1607FC1C",
    x"1607C708",
    x"16079208",
    x"16075D1E",
    x"16072848",
    x"1606F386",
    x"1606BED9",
    x"16068A41",
    x"160655BD",
    x"1606214E",
    x"1605ECF3",
    x"1605B8AD",
    x"1605847B",
    x"1605505E",
    x"16051C54",
    x"1604E85F",
    x"1604B47F",
    x"160480B2",
    x"16044CFA",
    x"16041956",
    x"1603E5C6",
    x"1603B24B",
    x"16037EE3",
    x"16034B90",
    x"16031850",
    x"1602E525",
    x"1602B20D",
    x"16027F09",
    x"16024C1A",
    x"1602193E",
    x"1601E676",
    x"1601B3C2",
    x"16018122",
    x"16014E95",
    x"16011C1C",
    x"1600E9B7",
    x"1600B766",
    x"16008528",
    x"160052FE",
    x"160020E7",
    x"15FFDDC8",
    x"15FF79E9",
    x"15FF1630",
    x"15FEB29F",
    x"15FE4F35",
    x"15FDEBF1",
    x"15FD88D4",
    x"15FD25DE",
    x"15FCC30F",
    x"15FC6066",
    x"15FBFDE4",
    x"15FB9B88",
    x"15FB3952",
    x"15FAD743",
    x"15FA755A",
    x"15FA1397",
    x"15F9B1FA",
    x"15F95084",
    x"15F8EF34",
    x"15F88E09",
    x"15F82D05",
    x"15F7CC26",
    x"15F76B6D",
    x"15F70ADA",
    x"15F6AA6D",
    x"15F64A25",
    x"15F5EA03",
    x"15F58A06",
    x"15F52A2F",
    x"15F4CA7D",
    x"15F46AF1",
    x"15F40B89",
    x"15F3AC48",
    x"15F34D2B",
    x"15F2EE33",
    x"15F28F61",
    x"15F230B3",
    x"15F1D22B",
    x"15F173C7",
    x"15F11588",
    x"15F0B76E",
    x"15F05979",
    x"15EFFBA8",
    x"15EF9DFC",
    x"15EF4075",
    x"15EEE312",
    x"15EE85D3",
    x"15EE28B9",
    x"15EDCBC4",
    x"15ED6EF2",
    x"15ED1245",
    x"15ECB5BC",
    x"15EC5957",
    x"15EBFD16",
    x"15EBA0F9",
    x"15EB4500",
    x"15EAE92B",
    x"15EA8D7A",
    x"15EA31ED",
    x"15E9D683",
    x"15E97B3D",
    x"15E9201B",
    x"15E8C51C",
    x"15E86A41",
    x"15E80F89",
    x"15E7B4F5",
    x"15E75A83",
    x"15E70036",
    x"15E6A60B",
    x"15E64C04",
    x"15E5F220",
    x"15E5985F",
    x"15E53EC1",
    x"15E4E546",
    x"15E48BEE",
    x"15E432B8",
    x"15E3D9A6",
    x"15E380B6",
    x"15E327E9",
    x"15E2CF3F",
    x"15E276B8",
    x"15E21E52",
    x"15E1C610",
    x"15E16DF0",
    x"15E115F2",
    x"15E0BE17",
    x"15E0665D",
    x"15E00EC7",
    x"15DFB752",
    x"15DF5FFF",
    x"15DF08CF",
    x"15DEB1C0",
    x"15DE5AD4",
    x"15DE0409",
    x"15DDAD61",
    x"15DD56DA",
    x"15DD0075",
    x"15DCAA32",
    x"15DC5410",
    x"15DBFE10",
    x"15DBA831",
    x"15DB5274",
    x"15DAFCD9",
    x"15DAA75F",
    x"15DA5206",
    x"15D9FCCF",
    x"15D9A7B9",
    x"15D952C4",
    x"15D8FDF0",
    x"15D8A93D",
    x"15D854AC",
    x"15D8003B",
    x"15D7ABEC",
    x"15D757BD",
    x"15D703AF",
    x"15D6AFC2",
    x"15D65BF6",
    x"15D6084A",
    x"15D5B4BF",
    x"15D56155",
    x"15D50E0B",
    x"15D4BAE2",
    x"15D467D9",
    x"15D414F1",
    x"15D3C229",
    x"15D36F81",
    x"15D31CFA",
    x"15D2CA92",
    x"15D2784B",
    x"15D22624",
    x"15D1D41E",
    x"15D18237",
    x"15D13070",
    x"15D0DEC9",
    x"15D08D42",
    x"15D03BDA",
    x"15CFEA93",
    x"15CF996B",
    x"15CF4863",
    x"15CEF77B",
    x"15CEA6B2",
    x"15CE5608",
    x"15CE057E",
    x"15CDB514",
    x"15CD64C9",
    x"15CD149D",
    x"15CCC491",
    x"15CC74A4",
    x"15CC24D6",
    x"15CBD527",
    x"15CB8597",
    x"15CB3627",
    x"15CAE6D5",
    x"15CA97A2",
    x"15CA488E",
    x"15C9F999",
    x"15C9AAC3",
    x"15C95C0C",
    x"15C90D73",
    x"15C8BEFA",
    x"15C8709E",
    x"15C82262",
    x"15C7D443",
    x"15C78644",
    x"15C73862",
    x"15C6EAA0",
    x"15C69CFB",
    x"15C64F75",
    x"15C6020D",
    x"15C5B4C3",
    x"15C56798",
    x"15C51A8A",
    x"15C4CD9B",
    x"15C480CA",
    x"15C43416",
    x"15C3E781",
    x"15C39B0A",
    x"15C34EB0",
    x"15C30274",
    x"15C2B656",
    x"15C26A56",
    x"15C21E73",
    x"15C1D2AE",
    x"15C18706",
    x"15C13B7C",
    x"15C0F010",
    x"15C0A4C1",
    x"15C0598F",
    x"15C00E7B",
    x"15BFC384",
    x"15BF78AA",
    x"15BF2DED",
    x"15BEE34E",
    x"15BE98CC",
    x"15BE4E67",
    x"15BE041F",
    x"15BDB9F3",
    x"15BD6FE5",
    x"15BD25F4",
    x"15BCDC20",
    x"15BC9268",
    x"15BC48CD",
    x"15BBFF4F",
    x"15BBB5EE",
    x"15BB6CA9",
    x"15BB2381",
    x"15BADA75",
    x"15BA9186",
    x"15BA48B4",
    x"15B9FFFD",
    x"15B9B764",
    x"15B96EE6",
    x"15B92685",
    x"15B8DE40",
    x"15B89617",
    x"15B84E0B",
    x"15B8061A",
    x"15B7BE46",
    x"15B7768E",
    x"15B72EF1",
    x"15B6E771",
    x"15B6A00C",
    x"15B658C4",
    x"15B61197",
    x"15B5CA86",
    x"15B58391",
    x"15B53CB7",
    x"15B4F5F9",
    x"15B4AF57",
    x"15B468D0",
    x"15B42265",
    x"15B3DC16",
    x"15B395E1",
    x"15B34FC8",
    x"15B309CB",
    x"15B2C3E9",
    x"15B27E22",
    x"15B23876",
    x"15B1F2E6",
    x"15B1AD70",
    x"15B16816",
    x"15B122D7",
    x"15B0DDB3",
    x"15B098AA",
    x"15B053BC",
    x"15B00EE8",
    x"15AFCA30",
    x"15AF8592",
    x"15AF4110",
    x"15AEFCA8",
    x"15AEB85A",
    x"15AE7428",
    x"15AE3010",
    x"15ADEC12",
    x"15ADA82F",
    x"15AD6467",
    x"15AD20B9",
    x"15ACDD25",
    x"15AC99AC",
    x"15AC564D",
    x"15AC1308",
    x"15ABCFDE",
    x"15AB8CCE",
    x"15AB49D8",
    x"15AB06FC",
    x"15AAC43B",
    x"15AA8193",
    x"15AA3F05",
    x"15A9FC92",
    x"15A9BA38",
    x"15A977F8",
    x"15A935D2",
    x"15A8F3C6",
    x"15A8B1D4",
    x"15A86FFB",
    x"15A82E3C",
    x"15A7EC97",
    x"15A7AB0B",
    x"15A76999",
    x"15A72841",
    x"15A6E702",
    x"15A6A5DC",
    x"15A664D0",
    x"15A623DE",
    x"15A5E304",
    x"15A5A244",
    x"15A5619E",
    x"15A52110",
    x"15A4E09C",
    x"15A4A041",
    x"15A45FFF",
    x"15A41FD6",
    x"15A3DFC6",
    x"15A39FCF",
    x"15A35FF1",
    x"15A3202C",
    x"15A2E080",
    x"15A2A0EC",
    x"15A26172",
    x"15A22210",
    x"15A1E2C7",
    x"15A1A397",
    x"15A1647F",
    x"15A12581",
    x"15A0E69A",
    x"15A0A7CC",
    x"15A06917",
    x"15A02A7A",
    x"159FEBF6",
    x"159FAD8A",
    x"159F6F36",
    x"159F30FB",
    x"159EF2D8",
    x"159EB4CD",
    x"159E76DB",
    x"159E3900",
    x"159DFB3E",
    x"159DBD94",
    x"159D8002",
    x"159D4288",
    x"159D0526",
    x"159CC7DC",
    x"159C8AAA",
    x"159C4D90",
    x"159C108D",
    x"159BD3A3",
    x"159B96D0",
    x"159B5A15",
    x"159B1D72",
    x"159AE0E6",
    x"159AA472",
    x"159A6815",
    x"159A2BD1",
    x"1599EFA3",
    x"1599B38D",
    x"1599778F",
    x"15993BA8",
    x"1598FFD8",
    x"1598C420",
    x"1598887F",
    x"15984CF5",
    x"15981183",
    x"1597D628",
    x"15979AE4",
    x"15975FB7",
    x"159724A1",
    x"1596E9A2",
    x"1596AEBA",
    x"159673E9",
    x"15963930",
    x"1595FE8D",
    x"1595C401",
    x"1595898C",
    x"15954F2D",
    x"159514E6",
    x"1594DAB5",
    x"1594A09B",
    x"15946698",
    x"15942CAB",
    x"1593F2D5",
    x"1593B915",
    x"15937F6C",
    x"159345D9",
    x"15930C5D",
    x"1592D2F8",
    x"159299A9",
    x"15926070",
    x"1592274D",
    x"1591EE41",
    x"1591B54B",
    x"15917C6B",
    x"159143A2",
    x"15910AEF",
    x"1590D251",
    x"159099CA",
    x"15906159",
    x"159028FE",
    x"158FF0B9",
    x"158FB88A",
    x"158F8071",
    x"158F486E",
    x"158F1080",
    x"158ED8A9",
    x"158EA0E7",
    x"158E693B",
    x"158E31A5",
    x"158DFA24",
    x"158DC2B9",
    x"158D8B64",
    x"158D5424",
    x"158D1CFA",
    x"158CE5E6",
    x"158CAEE7",
    x"158C77FD",
    x"158C4129",
    x"158C0A6A",
    x"158BD3C1",
    x"158B9D2D",
    x"158B66AE",
    x"158B3045",
    x"158AF9F0",
    x"158AC3B1",
    x"158A8D87",
    x"158A5773",
    x"158A2173",
    x"1589EB89",
    x"1589B5B3",
    x"15897FF3",
    x"15894A47",
    x"158914B1",
    x"1588DF2F",
    x"1588A9C2",
    x"1588746A",
    x"15883F27",
    x"158809F9",
    x"1587D4DF",
    x"15879FDB",
    x"15876AEB",
    x"1587360F",
    x"15870148",
    x"1586CC96",
    x"158697F8",
    x"1586636F",
    x"15862EFB",
    x"1585FA9B",
    x"1585C64F",
    x"15859218",
    x"15855DF5",
    x"158529E6",
    x"1584F5EC",
    x"1584C206",
    x"15848E35",
    x"15845A77",
    x"158426CE",
    x"1583F339",
    x"1583BFB8",
    x"15838C4B",
    x"158358F2",
    x"158325AD",
    x"1582F27D",
    x"1582BF60",
    x"15828C57",
    x"15825962",
    x"15822681",
    x"1581F3B4",
    x"1581C0FB",
    x"15818E55",
    x"15815BC4",
    x"15812946",
    x"1580F6DC",
    x"1580C485",
    x"15809242",
    x"15806013",
    x"15802DF7",
    x"157FF7DD",
    x"157F93F4",
    x"157F3032",
    x"157ECC96",
    x"157E6922",
    x"157E05D4",
    x"157DA2AD",
    x"157D3FAD",
    x"157CDCD4",
    x"157C7A21",
    x"157C1794",
    x"157BB52E",
    x"157B52EF",
    x"157AF0D5",
    x"157A8EE2",
    x"157A2D16",
    x"1579CB6F",
    x"157969EF",
    x"15790894",
    x"1578A760",
    x"15784652",
    x"1577E569",
    x"157784A6",
    x"15772409",
    x"1576C392",
    x"15766341",
    x"15760315",
    x"1575A30E",
    x"1575432D",
    x"1574E372",
    x"157483DC",
    x"1574246B",
    x"1573C51F",
    x"157365F9",
    x"157306F7",
    x"1572A81B",
    x"15724964",
    x"1571EAD2",
    x"15718C65",
    x"15712E1C",
    x"1570CFF9",
    x"157071FA",
    x"1570141F",
    x"156FB66A",
    x"156F58D9",
    x"156EFB6D",
    x"156E9E25",
    x"156E4101",
    x"156DE402",
    x"156D8727",
    x"156D2A70",
    x"156CCDDE",
    x"156C716F",
    x"156C1525",
    x"156BB8FF",
    x"156B5CFC",
    x"156B011E",
    x"156AA564",
    x"156A49CD",
    x"1569EE5A",
    x"1569930B",
    x"156937DF",
    x"1568DCD7",
    x"156881F2",
    x"15682731",
    x"1567CC94",
    x"1567721A",
    x"156717C3",
    x"1566BD8F",
    x"1566637F",
    x"15660991",
    x"1565AFC7",
    x"15655620",
    x"1564FC9C",
    x"1564A33B",
    x"156449FC",
    x"1563F0E1",
    x"156397E8",
    x"15633F12",
    x"1562E65F",
    x"15628DCE",
    x"15623560",
    x"1561DD14",
    x"156184EB",
    x"15612CE4",
    x"1560D500",
    x"15607D3E",
    x"1560259E",
    x"155FCE21",
    x"155F76C5",
    x"155F1F8C",
    x"155EC874",
    x"155E717F",
    x"155E1AAC",
    x"155DC3FA",
    x"155D6D6B",
    x"155D16FD",
    x"155CC0B1",
    x"155C6A86",
    x"155C147D",
    x"155BBE96",
    x"155B68D1",
    x"155B132C",
    x"155ABDAA",
    x"155A6848",
    x"155A1308",
    x"1559BDE9",
    x"155968EC",
    x"1559140F",
    x"1558BF54",
    x"15586ABA",
    x"15581641",
    x"1557C1E8",
    x"15576DB1",
    x"1557199B",
    x"1556C5A5",
    x"155671D0",
    x"15561E1C",
    x"1555CA89",
    x"15557716",
    x"155523C4",
    x"1554D092",
    x"15547D81",
    x"15542A90",
    x"1553D7BF",
    x"1553850F",
    x"1553327F",
    x"1552E010",
    x"15528DC0",
    x"15523B91",
    x"1551E982",
    x"15519793",
    x"155145C3",
    x"1550F414",
    x"1550A285",
    x"15505115",
    x"154FFFC5",
    x"154FAE95",
    x"154F5D85",
    x"154F0C94",
    x"154EBBC3",
    x"154E6B11",
    x"154E1A7F",
    x"154DCA0D",
    x"154D79BA",
    x"154D2986",
    x"154CD971",
    x"154C897C",
    x"154C39A6",
    x"154BE9EF",
    x"154B9A57",
    x"154B4ADE",
    x"154AFB84",
    x"154AAC4A",
    x"154A5D2E",
    x"154A0E31",
    x"1549BF53",
    x"15497093",
    x"154921F3",
    x"1548D371",
    x"1548850D",
    x"154836C9",
    x"1547E8A3",
    x"15479A9B",
    x"15474CB2",
    x"1546FEE7",
    x"1546B13B",
    x"154663AD",
    x"1546163D",
    x"1545C8EB",
    x"15457BB8",
    x"15452EA3",
    x"1544E1AB",
    x"154494D2",
    x"15444817",
    x"1543FB7A",
    x"1543AEFB",
    x"15436299",
    x"15431656",
    x"1542CA30",
    x"15427E28",
    x"1542323D",
    x"1541E670",
    x"15419AC1",
    x"15414F2F",
    x"154103BB",
    x"1540B865",
    x"15406D2B",
    x"1540220F",
    x"153FD711",
    x"153F8C2F",
    x"153F416B",
    x"153EF6C4",
    x"153EAC3A",
    x"153E61CD",
    x"153E177E",
    x"153DCD4B",
    x"153D8335",
    x"153D393D",
    x"153CEF61",
    x"153CA5A2",
    x"153C5BFF",
    x"153C127A",
    x"153BC911",
    x"153B7FC5",
    x"153B3695",
    x"153AED82",
    x"153AA48B",
    x"153A5BB1",
    x"153A12F4",
    x"1539CA53",
    x"153981CE",
    x"15393965",
    x"1538F119",
    x"1538A8E9",
    x"153860D5",
    x"153818DD",
    x"1537D101",
    x"15378942",
    x"1537419E",
    x"1536FA17",
    x"1536B2AB",
    x"15366B5B",
    x"15362427",
    x"1535DD0F",
    x"15359612",
    x"15354F31",
    x"1535086C",
    x"1534C1C3",
    x"15347B35",
    x"153434C3",
    x"1533EE6C",
    x"1533A830",
    x"15336210",
    x"15331C0C",
    x"1532D622",
    x"15329054",
    x"15324AA2",
    x"1532050A",
    x"1531BF8E",
    x"15317A2C",
    x"153134E6",
    x"1530EFBB",
    x"1530AAAB",
    x"153065B6",
    x"153020DB",
    x"152FDC1C",
    x"152F9777",
    x"152F52EE",
    x"152F0E7F",
    x"152ECA2A",
    x"152E85F1",
    x"152E41D2",
    x"152DFDCD",
    x"152DB9E3",
    x"152D7614",
    x"152D325F",
    x"152CEEC5",
    x"152CAB45",
    x"152C67DF",
    x"152C2493",
    x"152BE162",
    x"152B9E4B",
    x"152B5B4F",
    x"152B186C",
    x"152AD5A3",
    x"152A92F5",
    x"152A5061",
    x"152A0DE6",
    x"1529CB86",
    x"1529893F",
    x"15294712",
    x"15290500",
    x"1528C307",
    x"15288127",
    x"15283F62",
    x"1527FDB6",
    x"1527BC23",
    x"15277AAB",
    x"1527394C",
    x"1526F806",
    x"1526B6DA",
    x"152675C7",
    x"152634CE",
    x"1525F3EE",
    x"1525B327",
    x"1525727A",
    x"152531E6",
    x"1524F16B",
    x"1524B109",
    x"152470C1",
    x"15243091",
    x"1523F07B",
    x"1523B07D",
    x"15237099",
    x"152330CD",
    x"1522F11B",
    x"1522B181",
    x"15227200",
    x"15223298",
    x"1521F348",
    x"1521B412",
    x"152174F4",
    x"152135EE",
    x"1520F701",
    x"1520B82D",
    x"15207972",
    x"15203ACE",
    x"151FFC44",
    x"151FBDD1",
    x"151F7F77",
    x"151F4136",
    x"151F030C",
    x"151EC4FB",
    x"151E8702",
    x"151E4922",
    x"151E0B59",
    x"151DCDA9",
    x"151D9011",
    x"151D5290",
    x"151D1528",
    x"151CD7D8",
    x"151C9A9F",
    x"151C5D7F",
    x"151C2076",
    x"151BE386",
    x"151BA6AD",
    x"151B69EB",
    x"151B2D42",
    x"151AF0B0",
    x"151AB436",
    x"151A77D3",
    x"151A3B88",
    x"1519FF55",
    x"1519C339",
    x"15198734",
    x"15194B47",
    x"15190F71",
    x"1518D3B3",
    x"1518980C",
    x"15185C7C",
    x"15182104",
    x"1517E5A2",
    x"1517AA58",
    x"15176F25",
    x"15173409",
    x"1516F905",
    x"1516BE17",
    x"15168340",
    x"15164880",
    x"15160DD7",
    x"1515D346",
    x"151598CA",
    x"15155E66",
    x"15152419",
    x"1514E9E2",
    x"1514AFC2",
    x"151475B9",
    x"15143BC6",
    x"151401EA",
    x"1513C824",
    x"15138E76",
    x"151354DD",
    x"15131B5B",
    x"1512E1F0",
    x"1512A89B",
    x"15126F5C",
    x"15123634",
    x"1511FD22",
    x"1511C426",
    x"15118B40",
    x"15115271",
    x"151119B8",
    x"1510E115",
    x"1510A888",
    x"15107011",
    x"151037B1",
    x"150FFF66",
    x"150FC731",
    x"150F8F12",
    x"150F5709",
    x"150F1F16",
    x"150EE739",
    x"150EAF72",
    x"150E77C0",
    x"150E4024",
    x"150E089E",
    x"150DD12D",
    x"150D99D2",
    x"150D628D",
    x"150D2B5D",
    x"150CF443",
    x"150CBD3E",
    x"150C864F",
    x"150C4F76",
    x"150C18B1",
    x"150BE202",
    x"150BAB69",
    x"150B74E4",
    x"150B3E75",
    x"150B081B",
    x"150AD1D7",
    x"150A9BA8",
    x"150A658D",
    x"150A2F88",
    x"1509F998",
    x"1509C3BD",
    x"15098DF7",
    x"15095846",
    x"150922AA",
    x"1508ED23",
    x"1508B7B1",
    x"15088254",
    x"15084D0B",
    x"150817D7",
    x"1507E2B9",
    x"1507ADAE",
    x"150778B9",
    x"150743D8",
    x"15070F0C",
    x"1506DA54",
    x"1506A5B1",
    x"15067123",
    x"15063CA9",
    x"15060843",
    x"1505D3F2",
    x"15059FB6",
    x"15056B8E",
    x"1505377A",
    x"1505037A",
    x"1504CF8F",
    x"15049BB8",
    x"150467F5",
    x"15043447",
    x"150400AC",
    x"1503CD26",
    x"150399B4",
    x"15036656",
    x"1503330C",
    x"1502FFD6",
    x"1502CCB4",
    x"150299A6",
    x"150266AC",
    x"150233C6",
    x"150200F4",
    x"1501CE35",
    x"15019B8B",
    x"150168F4",
    x"15013671",
    x"15010401",
    x"1500D1A6",
    x"15009F5E",
    x"15006D29",
    x"15003B08",
    x"150008FB",
    x"14FFAE02",
    x"14FF4A36",
    x"14FEE690",
    x"14FE8312",
    x"14FE1FBA",
    x"14FDBC89",
    x"14FD597F",
    x"14FCF69B",
    x"14FC93DE",
    x"14FC3148",
    x"14FBCED7",
    x"14FB6C8E",
    x"14FB0A6B",
    x"14FAA86E",
    x"14FA4697",
    x"14F9E4E7",
    x"14F9835C",
    x"14F921F8",
    x"14F8C0BA",
    x"14F85FA1",
    x"14F7FEAF",
    x"14F79DE2",
    x"14F73D3C",
    x"14F6DCBA",
    x"14F67C5F",
    x"14F61C29",
    x"14F5BC19",
    x"14F55C2E",
    x"14F4FC69",
    x"14F49CC9",
    x"14F43D4F",
    x"14F3DDF9",
    x"14F37EC9",
    x"14F31FBE",
    x"14F2C0D8",
    x"14F26217",
    x"14F2037C",
    x"14F1A505",
    x"14F146B3",
    x"14F0E885",
    x"14F08A7D",
    x"14F02C99",
    x"14EFCEDA",
    x"14EF7140",
    x"14EF13CA",
    x"14EEB678",
    x"14EE594B",
    x"14EDFC42",
    x"14ED9F5E",
    x"14ED429E",
    x"14ECE602",
    x"14EC898A",
    x"14EC2D36",
    x"14EBD107",
    x"14EB74FB",
    x"14EB1913",
    x"14EABD50",
    x"14EA61AF",
    x"14EA0633",
    x"14E9AADB",
    x"14E94FA6",
    x"14E8F494",
    x"14E899A7",
    x"14E83EDC",
    x"14E7E435",
    x"14E789B2",
    x"14E72F52",
    x"14E6D515",
    x"14E67AFB",
    x"14E62105",
    x"14E5C732",
    x"14E56D81",
    x"14E513F4",
    x"14E4BA8A",
    x"14E46142",
    x"14E4081E",
    x"14E3AF1C",
    x"14E3563D",
    x"14E2FD81",
    x"14E2A4E7",
    x"14E24C70",
    x"14E1F41B",
    x"14E19BE9",
    x"14E143D9",
    x"14E0EBEC",
    x"14E09421",
    x"14E03C78",
    x"14DFE4F2",
    x"14DF8D8D",
    x"14DF364B",
    x"14DEDF2B",
    x"14DE882D",
    x"14DE3150",
    x"14DDDA96",
    x"14DD83FE",
    x"14DD2D87",
    x"14DCD732",
    x"14DC80FF",
    x"14DC2AED",
    x"14DBD4FD",
    x"14DB7F2F",
    x"14DB2982",
    x"14DAD3F6",
    x"14DA7E8C",
    x"14DA2944",
    x"14D9D41C",
    x"14D97F16",
    x"14D92A31",
    x"14D8D56D",
    x"14D880CA",
    x"14D82C48",
    x"14D7D7E7",
    x"14D783A8",
    x"14D72F89",
    x"14D6DB8A",
    x"14D687AD",
    x"14D633F0",
    x"14D5E054",
    x"14D58CD9",
    x"14D5397E",
    x"14D4E644",
    x"14D4932A",
    x"14D44031",
    x"14D3ED58",
    x"14D39AA0",
    x"14D34807",
    x"14D2F58F",
    x"14D2A338",
    x"14D25100",
    x"14D1FEE8",
    x"14D1ACF1",
    x"14D15B19",
    x"14D10962",
    x"14D0B7CA",
    x"14D06652",
    x"14D014FA",
    x"14CFC3C2",
    x"14CF72A9",
    x"14CF21B0",
    x"14CED0D7",
    x"14CE801D",
    x"14CE2F82",
    x"14CDDF08",
    x"14CD8EAC",
    x"14CD3E70",
    x"14CCEE53",
    x"14CC9E56",
    x"14CC4E78",
    x"14CBFEB9",
    x"14CBAF19",
    x"14CB5F98",
    x"14CB1036",
    x"14CAC0F3",
    x"14CA71CF",
    x"14CA22CA",
    x"14C9D3E4",
    x"14C9851D",
    x"14C93674",
    x"14C8E7EA",
    x"14C8997F",
    x"14C84B32",
    x"14C7FD04",
    x"14C7AEF4",
    x"14C76103",
    x"14C71331",
    x"14C6C57C",
    x"14C677E6",
    x"14C62A6F",
    x"14C5DD15",
    x"14C58FDA",
    x"14C542BD",
    x"14C4F5BE",
    x"14C4A8DD",
    x"14C45C1A",
    x"14C40F75",
    x"14C3C2EE",
    x"14C37685",
    x"14C32A39",
    x"14C2DE0C",
    x"14C291FC",
    x"14C24609",
    x"14C1FA35",
    x"14C1AE7E",
    x"14C162E5",
    x"14C11769",
    x"14C0CC0A",
    x"14C080C9",
    x"14C035A6",
    x"14BFEA9F",
    x"14BF9FB6",
    x"14BF54EB",
    x"14BF0A3C",
    x"14BEBFAB",
    x"14BE7536",
    x"14BE2ADF",
    x"14BDE0A5",
    x"14BD9687",
    x"14BD4C87",
    x"14BD02A4",
    x"14BCB8DD",
    x"14BC6F33",
    x"14BC25A6",
    x"14BBDC36",
    x"14BB92E2",
    x"14BB49AB",
    x"14BB0091",
    x"14BAB793",
    x"14BA6EB1",
    x"14BA25EC",
    x"14B9DD43",
    x"14B994B7",
    x"14B94C47",
    x"14B903F4",
    x"14B8BBBC",
    x"14B873A1",
    x"14B82BA2",
    x"14B7E3BF",
    x"14B79BF8",
    x"14B7544D",
    x"14B70CBE",
    x"14B6C54B",
    x"14B67DF4",
    x"14B636B9",
    x"14B5EF99",
    x"14B5A895",
    x"14B561AD",
    x"14B51AE1",
    x"14B4D430",
    x"14B48D9B",
    x"14B44722",
    x"14B400C4",
    x"14B3BA81",
    x"14B3745A",
    x"14B32E4E",
    x"14B2E85E",
    x"14B2A289",
    x"14B25CCF",
    x"14B21730",
    x"14B1D1AD",
    x"14B18C44",
    x"14B146F7",
    x"14B101C5",
    x"14B0BCAE",
    x"14B077B1",
    x"14B032D0",
    x"14AFEE0A",
    x"14AFA95E",
    x"14AF64CD",
    x"14AF2057",
    x"14AEDBFC",
    x"14AE97BB",
    x"14AE5396",
    x"14AE0F8A",
    x"14ADCB99",
    x"14AD87C3",
    x"14AD4407",
    x"14AD0066",
    x"14ACBCDF",
    x"14AC7972",
    x"14AC3620",
    x"14ABF2E8",
    x"14ABAFCA",
    x"14AB6CC7",
    x"14AB29DD",
    x"14AAE70E",
    x"14AAA459",
    x"14AA61BE",
    x"14AA1F3C",
    x"14A9DCD5",
    x"14A99A88",
    x"14A95854",
    x"14A9163B",
    x"14A8D43B",
    x"14A89255",
    x"14A85089",
    x"14A80ED6",
    x"14A7CD3D",
    x"14A78BBE",
    x"14A74A58",
    x"14A7090C",
    x"14A6C7D9",
    x"14A686BF",
    x"14A645C0",
    x"14A604D9",
    x"14A5C40C",
    x"14A58358",
    x"14A542BD",
    x"14A5023C",
    x"14A4C1D3",
    x"14A48184",
    x"14A4414E",
    x"14A40131",
    x"14A3C12D",
    x"14A38142",
    x"14A34170",
    x"14A301B7",
    x"14A2C217",
    x"14A2828F",
    x"14A24321",
    x"14A203CB",
    x"14A1C48E",
    x"14A18569",
    x"14A1465E",
    x"14A1076A",
    x"14A0C890",
    x"14A089CE",
    x"14A04B24",
    x"14A00C93",
    x"149FCE1A",
    x"149F8FBA",
    x"149F5172",
    x"149F1342",
    x"149ED52B",
    x"149E972C",
    x"149E5945",
    x"149E1B76",
    x"149DDDBF",
    x"149DA021",
    x"149D629A",
    x"149D252C",
    x"149CE7D5",
    x"149CAA97",
    x"149C6D70",
    x"149C3061",
    x"149BF36A",
    x"149BB68B",
    x"149B79C4",
    x"149B3D14",
    x"149B007C",
    x"149AC3FB",
    x"149A8793",
    x"149A4B41",
    x"149A0F08",
    x"1499D2E6",
    x"149996DB",
    x"14995AE8",
    x"14991F0C",
    x"1498E348",
    x"1498A79A",
    x"14986C05",
    x"14983086",
    x"1497F51F",
    x"1497B9CF",
    x"14977E96",
    x"14974374",
    x"14970869",
    x"1496CD75",
    x"14969298",
    x"149657D3",
    x"14961D24",
    x"1495E28C",
    x"1495A80B",
    x"14956DA0",
    x"1495334D",
    x"1494F910",
    x"1494BEEA",
    x"149484DB",
    x"14944AE3",
    x"14941101",
    x"1493D735",
    x"14939D81",
    x"149363E2",
    x"14932A5B",
    x"1492F0E9",
    x"1492B78E",
    x"14927E4A",
    x"1492451C",
    x"14920C04",
    x"1491D302",
    x"14919A17",
    x"14916142",
    x"14912883",
    x"1490EFDA",
    x"1490B748",
    x"14907ECB",
    x"14904664",
    x"14900E14",
    x"148FD5D9",
    x"148F9DB5",
    x"148F65A6",
    x"148F2DAD",
    x"148EF5CB",
    x"148EBDFD",
    x"148E8646",
    x"148E4EA5",
    x"148E1719",
    x"148DDFA2",
    x"148DA842",
    x"148D70F7",
    x"148D39C2",
    x"148D02A2",
    x"148CCB98",
    x"148C94A3",
    x"148C5DC3",
    x"148C26FA",
    x"148BF045",
    x"148BB9A6",
    x"148B831C",
    x"148B4CA7",
    x"148B1648",
    x"148ADFFE",
    x"148AA9C9",
    x"148A73A9",
    x"148A3D9F",
    x"148A07A9",
    x"1489D1C9",
    x"14899BFD",
    x"14896647",
    x"148930A5",
    x"1488FB19",
    x"1488C5A1",
    x"1488903E",
    x"14885AF0",
    x"148825B7",
    x"1487F093",
    x"1487BB83",
    x"14878688",
    x"148751A2",
    x"14871CD1",
    x"1486E814",
    x"1486B36B",
    x"14867ED8",
    x"14864A58",
    x"148615ED",
    x"1485E197",
    x"1485AD55",
    x"14857928",
    x"1485450F",
    x"1485110A",
    x"1484DD19",
    x"1484A93D",
    x"14847575",
    x"148441C1",
    x"14840E22",
    x"1483DA96",
    x"1483A71F",
    x"148373BC",
    x"1483406C",
    x"14830D31",
    x"1482DA0A",
    x"1482A6F7",
    x"148273F8",
    x"1482410C",
    x"14820E35",
    x"1481DB71",
    x"1481A8C1",
    x"14817625",
    x"1481439D",
    x"14811128",
    x"1480DEC8",
    x"1480AC7A",
    x"14807A41",
    x"1480481B",
    x"14801609",
    x"147FC813",
    x"147F643D",
    x"147F008D",
    x"147E9D04",
    x"147E39A2",
    x"147DD667",
    x"147D7353",
    x"147D1065",
    x"147CAD9E",
    x"147C4AFD",
    x"147BE883",
    x"147B8630",
    x"147B2403",
    x"147AC1FC",
    x"147A601B",
    x"1479FE61",
    x"14799CCC",
    x"14793B5E",
    x"1478DA16",
    x"147878F4",
    x"147817F7",
    x"1477B721",
    x"14775670",
    x"1476F5E5",
    x"14769580",
    x"14763540",
    x"1475D526",
    x"14757532",
    x"14751563",
    x"1474B5B9",
    x"14745635",
    x"1473F6D6",
    x"1473979C",
    x"14733887",
    x"1472D998",
    x"14727ACD",
    x"14721C28",
    x"1471BDA7",
    x"14715F4C",
    x"14710115",
    x"1470A303",
    x"14704516",
    x"146FE74D",
    x"146F89A9",
    x"146F2C29",
    x"146ECECE",
    x"146E7198",
    x"146E1486",
    x"146DB798",
    x"146D5ACE",
    x"146CFE29",
    x"146CA1A7",
    x"146C454A",
    x"146BE911",
    x"146B8CFC",
    x"146B310B",
    x"146AD53E",
    x"146A7995",
    x"146A1E0F",
    x"1469C2AD",
    x"1469676F",
    x"14690C54",
    x"1468B15D",
    x"1468568A",
    x"1467FBDA",
    x"1467A14D",
    x"146746E4",
    x"1466EC9D",
    x"1466927B",
    x"1466387B",
    x"1465DE9F",
    x"146584E5",
    x"14652B4F",
    x"1464D1DB",
    x"1464788B",
    x"14641F5D",
    x"1463C652",
    x"14636D6A",
    x"146314A5",
    x"1462BC02",
    x"14626382",
    x"14620B24",
    x"1461B2E9",
    x"14615AD0",
    x"146102DA",
    x"1460AB06",
    x"14605354",
    x"145FFBC5",
    x"145FA458",
    x"145F4D0D",
    x"145EF5E4",
    x"145E9EDC",
    x"145E47F7",
    x"145DF134",
    x"145D9A93",
    x"145D4413",
    x"145CEDB6",
    x"145C977A",
    x"145C415F",
    x"145BEB67",
    x"145B958F",
    x"145B3FDA",
    x"145AEA46",
    x"145A94D3",
    x"145A3F81",
    x"1459EA51",
    x"14599542",
    x"14594055",
    x"1458EB88",
    x"145896DC",
    x"14584252",
    x"1457EDE9",
    x"145799A0",
    x"14574579",
    x"1456F172",
    x"14569D8C",
    x"145649C7",
    x"1455F622",
    x"1455A29E",
    x"14554F3B",
    x"1454FBF9",
    x"1454A8D6",
    x"145455D5",
    x"145402F3",
    x"1453B032",
    x"14535D92",
    x"14530B11",
    x"1452B8B1",
    x"14526671",
    x"14521451",
    x"1451C251",
    x"14517071",
    x"14511EB1",
    x"1450CD11",
    x"14507B91",
    x"14502A31",
    x"144FD8F0",
    x"144F87CF",
    x"144F36CE",
    x"144EE5EC",
    x"144E952A",
    x"144E4488",
    x"144DF405",
    x"144DA3A1",
    x"144D535D",
    x"144D0338",
    x"144CB332",
    x"144C634C",
    x"144C1385",
    x"144BC3DD",
    x"144B7454",
    x"144B24EA",
    x"144AD59F",
    x"144A8673",
    x"144A3766",
    x"1449E877",
    x"144999A8",
    x"14494AF7",
    x"1448FC66",
    x"1448ADF2",
    x"14485F9E",
    x"14481168",
    x"1447C350",
    x"14477557",
    x"1447277C",
    x"1446D9C0",
    x"14468C22",
    x"14463EA3",
    x"1445F141",
    x"1445A3FE",
    x"144556D9",
    x"144509D2",
    x"1444BCE9",
    x"1444701F",
    x"14442372",
    x"1443D6E3",
    x"14438A72",
    x"14433E1F",
    x"1442F1E9",
    x"1442A5D2",
    x"144259D8",
    x"14420DFC",
    x"1441C23D",
    x"1441769C",
    x"14412B18",
    x"1440DFB2",
    x"14409469",
    x"1440493E",
    x"143FFE30",
    x"143FB33F",
    x"143F686C",
    x"143F1DB6",
    x"143ED31D",
    x"143E88A1",
    x"143E3E42",
    x"143DF400",
    x"143DA9DB",
    x"143D5FD4",
    x"143D15E9",
    x"143CCC1A",
    x"143C8269",
    x"143C38D5",
    x"143BEF5D",
    x"143BA602",
    x"143B5CC3",
    x"143B13A1",
    x"143ACA9C",
    x"143A81B3",
    x"143A38E6",
    x"1439F036",
    x"1439A7A3",
    x"14395F2B",
    x"143916D0",
    x"1438CE91",
    x"1438866F",
    x"14383E68",
    x"1437F67E",
    x"1437AEB0",
    x"143766FE",
    x"14371F67",
    x"1436D7ED",
    x"1436908F",
    x"1436494C",
    x"14360225",
    x"1435BB1A",
    x"1435742B",
    x"14352D58",
    x"1434E6A0",
    x"1434A003",
    x"14345983",
    x"1434131E",
    x"1433CCD4",
    x"143386A5",
    x"14334093",
    x"1432FA9B",
    x"1432B4BF",
    x"14326EFE",
    x"14322958",
    x"1431E3CD",
    x"14319E5E",
    x"1431590A",
    x"143113D0",
    x"1430CEB2",
    x"143089AF",
    x"143044C7",
    x"142FFFF9",
    x"142FBB47",
    x"142F76AF",
    x"142F3232",
    x"142EEDD0",
    x"142EA988",
    x"142E655B",
    x"142E2149",
    x"142DDD51",
    x"142D9974",
    x"142D55B1",
    x"142D1209",
    x"142CCE7B",
    x"142C8B08",
    x"142C47AF",
    x"142C0470",
    x"142BC14B",
    x"142B7E41",
    x"142B3B50",
    x"142AF87A",
    x"142AB5BE",
    x"142A731C",
    x"142A3094",
    x"1429EE26",
    x"1429ABD2",
    x"14296998",
    x"14292778",
    x"1428E571",
    x"1428A385",
    x"142861B2",
    x"14281FF8",
    x"1427DE59",
    x"14279CD2",
    x"14275B66",
    x"14271A13",
    x"1426D8DA",
    x"142697BA",
    x"142656B3",
    x"142615C6",
    x"1425D4F2",
    x"14259438",
    x"14255396",
    x"1425130E",
    x"1424D29F",
    x"1424924A",
    x"1424520D",
    x"142411EA",
    x"1423D1DF",
    x"142391EE",
    x"14235215",
    x"14231255",
    x"1422D2AF",
    x"14229321",
    x"142253AC",
    x"1422144F",
    x"1421D50C",
    x"142195E1",
    x"142156CF",
    x"142117D5",
    x"1420D8F4",
    x"14209A2C",
    x"14205B7C",
    x"14201CE4",
    x"141FDE65",
    x"141F9FFE",
    x"141F61B0",
    x"141F237A",
    x"141EE55C",
    x"141EA757",
    x"141E696A",
    x"141E2B94",
    x"141DEDD8",
    x"141DB033",
    x"141D72A6",
    x"141D3531",
    x"141CF7D4",
    x"141CBA8F",
    x"141C7D63",
    x"141C404D",
    x"141C0350",
    x"141BC66B",
    x"141B899D",
    x"141B4CE7",
    x"141B1049",
    x"141AD3C3",
    x"141A9754",
    x"141A5AFC",
    x"141A1EBD",
    x"1419E294",
    x"1419A684",
    x"14196A8A",
    x"14192EA8",
    x"1418F2DE",
    x"1418B72B",
    x"14187B8F",
    x"1418400A",
    x"1418049D",
    x"1417C946",
    x"14178E07",
    x"141752DF",
    x"141717CF",
    x"1416DCD5",
    x"1416A1F2",
    x"14166726",
    x"14162C71",
    x"1415F1D4",
    x"1415B74D",
    x"14157CDC",
    x"14154283",
    x"14150840",
    x"1414CE15",
    x"141493FF",
    x"14145A01",
    x"14142019",
    x"1413E648",
    x"1413AC8D",
    x"141372E9",
    x"1413395B",
    x"1412FFE4",
    x"1412C683",
    x"14128D39",
    x"14125405",
    x"14121AE7",
    x"1411E1E0",
    x"1411A8EF",
    x"14117014",
    x"1411374F",
    x"1410FEA1",
    x"1410C608",
    x"14108D86",
    x"1410551A",
    x"14101CC4",
    x"140FE483",
    x"140FAC59",
    x"140F7445",
    x"140F3C46",
    x"140F045E",
    x"140ECC8B",
    x"140E94CE",
    x"140E5D27",
    x"140E2595",
    x"140DEE19",
    x"140DB6B3",
    x"140D7F62",
    x"140D4827",
    x"140D1102",
    x"140CD9F2",
    x"140CA2F8",
    x"140C6C13",
    x"140C3543",
    x"140BFE89",
    x"140BC7E4",
    x"140B9155",
    x"140B5ADB",
    x"140B2476",
    x"140AEE26",
    x"140AB7EC",
    x"140A81C7",
    x"140A4BB7",
    x"140A15BC",
    x"1409DFD6",
    x"1409AA05",
    x"14097449",
    x"14093EA2",
    x"14090910",
    x"1408D393",
    x"14089E2B",
    x"140868D7",
    x"14083399",
    x"1407FE6F",
    x"1407C95A",
    x"1407945A",
    x"14075F6E",
    x"14072A97",
    x"1406F5D5",
    x"1406C127",
    x"14068C8E",
    x"14065809",
    x"14062399",
    x"1405EF3D",
    x"1405BAF6",
    x"140586C3",
    x"140552A5",
    x"14051E9B",
    x"1404EAA5",
    x"1404B6C3",
    x"140482F6",
    x"14044F3D",
    x"14041B98",
    x"1403E807",
    x"1403B48B",
    x"14038122",
    x"14034DCE",
    x"14031A8E",
    x"1402E761",
    x"1402B449",
    x"14028144",
    x"14024E54",
    x"14021B77",
    x"1401E8AE",
    x"1401B5F9",
    x"14018358",
    x"140150CB",
    x"14011E51",
    x"1400EBEB",
    x"1400B999",
    x"1400875A",
    x"1400552F",
    x"14002317",
    x"13FFE227",
    x"13FF7E46",
    x"13FF1A8C",
    x"13FEB6F9",
    x"13FE538D",
    x"13FDF048",
    x"13FD8D2A",
    x"13FD2A32",
    x"13FCC761",
    x"13FC64B6",
    x"13FC0232",
    x"13FB9FD4",
    x"13FB3D9D",
    x"13FADB8C",
    x"13FA79A1",
    x"13FA17DD",
    x"13F9B63F",
    x"13F954C7",
    x"13F8F375",
    x"13F89248",
    x"13F83142",
    x"13F7D062",
    x"13F76FA7",
    x"13F70F13",
    x"13F6AEA4",
    x"13F64E5A",
    x"13F5EE36",
    x"13F58E38",
    x"13F52E5F",
    x"13F4CEAC",
    x"13F46F1E",
    x"13F40FB5",
    x"13F3B072",
    x"13F35153",
    x"13F2F25A",
    x"13F29386",
    x"13F234D7",
    x"13F1D64D",
    x"13F177E7",
    x"13F119A7",
    x"13F0BB8B",
    x"13F05D94",
    x"13EFFFC2",
    x"13EFA214",
    x"13EF448B",
    x"13EEE727",
    x"13EE89E7",
    x"13EE2CCB",
    x"13EDCFD4",
    x"13ED7301",
    x"13ED1652",
    x"13ECB9C7",
    x"13EC5D61",
    x"13EC011E",
    x"13EBA500",
    x"13EB4905",
    x"13EAED2F",
    x"13EA917C",
    x"13EA35ED",
    x"13E9DA82",
    x"13E97F3A",
    x"13E92417",
    x"13E8C916",
    x"13E86E39",
    x"13E81380",
    x"13E7B8EA",
    x"13E75E78",
    x"13E70428",
    x"13E6A9FC",
    x"13E64FF4",
    x"13E5F60E",
    x"13E59C4B",
    x"13E542AC",
    x"13E4E92F",
    x"13E48FD6",
    x"13E4369F",
    x"13E3DD8B",
    x"13E3849A",
    x"13E32BCB",
    x"13E2D31F",
    x"13E27A96",
    x"13E22230",
    x"13E1C9EC",
    x"13E171CA",
    x"13E119CB",
    x"13E0C1EE",
    x"13E06A33",
    x"13E0129B",
    x"13DFBB25",
    x"13DF63D1",
    x"13DF0C9F",
    x"13DEB58F",
    x"13DE5EA1",
    x"13DE07D5",
    x"13DDB12B",
    x"13DD5AA2",
    x"13DD043C",
    x"13DCADF7",
    x"13DC57D4",
    x"13DC01D2",
    x"13DBABF2",
    x"13DB5634",
    x"13DB0097",
    x"13DAAB1B",
    x"13DA55C1",
    x"13DA0088",
    x"13D9AB71",
    x"13D9567B",
    x"13D901A5",
    x"13D8ACF1",
    x"13D8585E",
    x"13D803EC",
    x"13D7AF9B",
    x"13D75B6B",
    x"13D7075C",
    x"13D6B36D",
    x"13D65F9F",
    x"13D60BF2",
    x"13D5B866",
    x"13D564FA",
    x"13D511AF",
    x"13D4BE85",
    x"13D46B7A",
    x"13D41891",
    x"13D3C5C7",
    x"13D3731E",
    x"13D32095",
    x"13D2CE2D",
    x"13D27BE4",
    x"13D229BC",
    x"13D1D7B3",
    x"13D185CB",
    x"13D13403",
    x"13D0E25B",
    x"13D090D2",
    x"13D03F69",
    x"13CFEE21",
    x"13CF9CF7",
    x"13CF4BEE",
    x"13CEFB04",
    x"13CEAA3A",
    x"13CE598F",
    x"13CE0904",
    x"13CDB898",
    x"13CD684C",
    x"13CD181E",
    x"13CCC811",
    x"13CC7822",
    x"13CC2853",
    x"13CBD8A3",
    x"13CB8912",
    x"13CB39A0",
    x"13CAEA4D",
    x"13CA9B18",
    x"13CA4C03",
    x"13C9FD0D",
    x"13C9AE36",
    x"13C95F7D",
    x"13C910E3",
    x"13C8C268",
    x"13C8740B",
    x"13C825CD",
    x"13C7D7AE",
    x"13C789AD",
    x"13C73BCA",
    x"13C6EE06",
    x"13C6A060",
    x"13C652D9",
    x"13C6056F",
    x"13C5B824",
    x"13C56AF7",
    x"13C51DE9",
    x"13C4D0F8",
    x"13C48425",
    x"13C43771",
    x"13C3EADA",
    x"13C39E61",
    x"13C35206",
    x"13C305C9",
    x"13C2B9AA",
    x"13C26DA8",
    x"13C221C4",
    x"13C1D5FE",
    x"13C18A55",
    x"13C13ECA",
    x"13C0F35C",
    x"13C0A80B",
    x"13C05CD9",
    x"13C011C3",
    x"13BFC6CB",
    x"13BF7BF0",
    x"13BF3132",
    x"13BEE691",
    x"13BE9C0E",
    x"13BE51A7",
    x"13BE075E",
    x"13BDBD31",
    x"13BD7322",
    x"13BD2930",
    x"13BCDF5A",
    x"13BC95A1",
    x"13BC4C05",
    x"13BC0286",
    x"13BBB923",
    x"13BB6FDD",
    x"13BB26B4",
    x"13BADDA7",
    x"13BA94B6",
    x"13BA4BE2",
    x"13BA032B",
    x"13B9BA90",
    x"13B97211",
    x"13B929AF",
    x"13B8E169",
    x"13B8993F",
    x"13B85131",
    x"13B8093F",
    x"13B7C16A",
    x"13B779B0",
    x"13B73213",
    x"13B6EA91",
    x"13B6A32B",
    x"13B65BE2",
    x"13B614B4",
    x"13B5CDA1",
    x"13B586AB",
    x"13B53FD0",
    x"13B4F911",
    x"13B4B26E",
    x"13B46BE6",
    x"13B42579",
    x"13B3DF28",
    x"13B398F3",
    x"13B352D9",
    x"13B30CDA",
    x"13B2C6F7",
    x"13B2812F",
    x"13B23B82",
    x"13B1F5F0",
    x"13B1B07A",
    x"13B16B1E",
    x"13B125DE",
    x"13B0E0B9",
    x"13B09BAE",
    x"13B056BF",
    x"13B011EB",
    x"13AFCD31",
    x"13AF8892",
    x"13AF440E",
    x"13AEFFA5",
    x"13AEBB57",
    x"13AE7723",
    x"13AE330A",
    x"13ADEF0B",
    x"13ADAB27",
    x"13AD675D",
    x"13AD23AE",
    x"13ACE019",
    x"13AC9C9F",
    x"13AC593F",
    x"13AC15F9",
    x"13ABD2CE",
    x"13AB8FBC",
    x"13AB4CC5",
    x"13AB09E8",
    x"13AAC726",
    x"13AA847D",
    x"13AA41EE",
    x"13A9FF79",
    x"13A9BD1F",
    x"13A97ADE",
    x"13A938B7",
    x"13A8F6A9",
    x"13A8B4B6",
    x"13A872DC",
    x"13A8311C",
    x"13A7EF76",
    x"13A7ADE9",
    x"13A76C76",
    x"13A72B1C",
    x"13A6E9DC",
    x"13A6A8B6",
    x"13A667A8",
    x"13A626B5",
    x"13A5E5DA",
    x"13A5A519",
    x"13A56471",
    x"13A523E2",
    x"13A4E36D",
    x"13A4A311",
    x"13A462CE",
    x"13A422A4",
    x"13A3E293",
    x"13A3A29B",
    x"13A362BB",
    x"13A322F5",
    x"13A2E348",
    x"13A2A3B4",
    x"13A26438",
    x"13A224D6",
    x"13A1E58B",
    x"13A1A65A",
    x"13A16742",
    x"13A12841",
    x"13A0E95A",
    x"13A0AA8B",
    x"13A06BD5",
    x"13A02D37",
    x"139FEEB1",
    x"139FB044",
    x"139F71F0",
    x"139F33B3",
    x"139EF58F",
    x"139EB784",
    x"139E7990",
    x"139E3BB5",
    x"139DFDF1",
    x"139DC046",
    x"139D82B3",
    x"139D4538",
    x"139D07D5",
    x"139CCA8A",
    x"139C8D57",
    x"139C503B",
    x"139C1338",
    x"139BD64C",
    x"139B9979",
    x"139B5CBD",
    x"139B2018",
    x"139AE38B",
    x"139AA716",
    x"139A6AB9",
    x"139A2E73",
    x"1399F245",
    x"1399B62E",
    x"13997A2E",
    x"13993E46",
    x"13990276",
    x"1398C6BC",
    x"13988B1A",
    x"13984F90",
    x"1398141C",
    x"1397D8C0",
    x"13979D7B",
    x"1397624D",
    x"13972736",
    x"1396EC36",
    x"1396B14D",
    x"1396767C",
    x"13963BC1",
    x"1396011D",
    x"1395C690",
    x"13958C1A",
    x"139551BB",
    x"13951772",
    x"1394DD40",
    x"1394A325",
    x"13946921",
    x"13942F33",
    x"1393F55C",
    x"1393BB9B",
    x"139381F1",
    x"1393485E",
    x"13930EE1",
    x"1392D57A",
    x"13929C2A",
    x"139262F0",
    x"139229CD",
    x"1391F0BF",
    x"1391B7C9",
    x"13917EE8",
    x"1391461D",
    x"13910D69",
    x"1390D4CB",
    x"13909C43",
    x"139063D1",
    x"13902B75",
    x"138FF32F",
    x"138FBAFF",
    x"138F82E5",
    x"138F4AE1",
    x"138F12F2",
    x"138EDB1A",
    x"138EA357",
    x"138E6BAA",
    x"138E3413",
    x"138DFC91",
    x"138DC526",
    x"138D8DCF",
    x"138D568F",
    x"138D1F64",
    x"138CE84E",
    x"138CB14E",
    x"138C7A64",
    x"138C438F",
    x"138C0CCF",
    x"138BD625",
    x"138B9F90",
    x"138B6910",
    x"138B32A6",
    x"138AFC50",
    x"138AC610",
    x"138A8FE6",
    x"138A59D0",
    x"138A23CF",
    x"1389EDE4",
    x"1389B80E",
    x"1389824C",
    x"13894CA0",
    x"13891708",
    x"1388E186",
    x"1388AC18",
    x"138876BF",
    x"1388417B",
    x"13880C4C",
    x"1387D732",
    x"1387A22C",
    x"13876D3B",
    x"1387385F",
    x"13870397",
    x"1386CEE4",
    x"13869A45",
    x"138665BB",
    x"13863146",
    x"1385FCE5",
    x"1385C898",
    x"13859460",
    x"1385603C",
    x"13852C2D",
    x"1384F832",
    x"1384C44B",
    x"13849078",
    x"13845CBA",
    x"13842910",
    x"1383F57A",
    x"1383C1F8",
    x"13838E8A",
    x"13835B31",
    x"138327EB",
    x"1382F4BA",
    x"1382C19C",
    x"13828E92",
    x"13825B9D",
    x"138228BB",
    x"1381F5ED",
    x"1381C333",
    x"1381908C",
    x"13815DFA",
    x"13812B7B",
    x"1380F910",
    x"1380C6B8",
    x"13809474",
    x"13806244",
    x"13803028",
    x"137FFC3D",
    x"137F9852",
    x"137F348E",
    x"137ED0F1",
    x"137E6D7B",
    x"137E0A2C",
    x"137DA703",
    x"137D4401",
    x"137CE126",
    x"137C7E71",
    x"137C1BE3",
    x"137BB97B",
    x"137B573A",
    x"137AF51F",
    x"137A932B",
    x"137A315C",
    x"1379CFB4",
    x"13796E32",
    x"13790CD6",
    x"1378ABA0",
    x"13784A90",
    x"1377E9A6",
    x"137788E1",
    x"13772843",
    x"1376C7CA",
    x"13766777",
    x"13760749",
    x"1375A741",
    x"1375475E",
    x"1374E7A1",
    x"13748809",
    x"13742897",
    x"1373C94A",
    x"13736A21",
    x"13730B1F",
    x"1372AC41",
    x"13724D88",
    x"1371EEF4",
    x"13719085",
    x"1371323B",
    x"1370D416",
    x"13707616",
    x"1370183A",
    x"136FBA83",
    x"136F5CF0",
    x"136EFF82",
    x"136EA238",
    x"136E4513",
    x"136DE812",
    x"136D8B36",
    x"136D2E7E",
    x"136CD1EA",
    x"136C757A",
    x"136C192E",
    x"136BBD06",
    x"136B6102",
    x"136B0522",
    x"136AA966",
    x"136A4DCE",
    x"1369F259",
    x"13699708",
    x"13693BDB",
    x"1368E0D2",
    x"136885EC",
    x"13682B29",
    x"1367D08A",
    x"1367760E",
    x"13671BB6",
    x"1366C180",
    x"1366676E",
    x"13660D80",
    x"1365B3B4",
    x"13655A0B",
    x"13650085",
    x"1364A723",
    x"13644DE3",
    x"1363F4C6",
    x"13639BCC",
    x"136342F4",
    x"1362EA3F",
    x"136291AD",
    x"1362393D",
    x"1361E0F0",
    x"136188C6",
    x"136130BD",
    x"1360D8D8",
    x"13608114",
    x"13602973",
    x"135FD1F4",
    x"135F7A97",
    x"135F235C",
    x"135ECC43",
    x"135E754C",
    x"135E1E77",
    x"135DC7C4",
    x"135D7133",
    x"135D1AC4",
    x"135CC476",
    x"135C6E4B",
    x"135C1840",
    x"135BC258",
    x"135B6C90",
    x"135B16EB",
    x"135AC166",
    x"135A6C04",
    x"135A16C2",
    x"1359C1A2",
    x"13596CA3",
    x"135917C5",
    x"1358C308",
    x"13586E6D",
    x"135819F2",
    x"1357C598",
    x"13577160",
    x"13571D48",
    x"1356C951",
    x"1356757A",
    x"135621C5",
    x"1355CE30",
    x"13557ABC",
    x"13552768",
    x"1354D435",
    x"13548122",
    x"13542E30",
    x"1353DB5E",
    x"135388AD",
    x"1353361B",
    x"1352E3AA",
    x"13529159",
    x"13523F29",
    x"1351ED18",
    x"13519B28",
    x"13514957",
    x"1350F7A6",
    x"1350A615",
    x"135054A4",
    x"13500353",
    x"134FB222",
    x"134F6110",
    x"134F101E",
    x"134EBF4B",
    x"134E6E99",
    x"134E1E05",
    x"134DCD91",
    x"134D7D3C",
    x"134D2D07",
    x"134CDCF1",
    x"134C8CFB",
    x"134C3D23",
    x"134BED6B",
    x"134B9DD2",
    x"134B4E57",
    x"134AFEFC",
    x"134AAFC0",
    x"134A60A3",
    x"134A11A5",
    x"1349C2C5",
    x"13497405",
    x"13492563",
    x"1348D6DF",
    x"1348887B",
    x"13483A35",
    x"1347EC0D",
    x"13479E04",
    x"1347501A",
    x"1347024E",
    x"1346B4A0",
    x"13466711",
    x"1346199F",
    x"1345CC4C",
    x"13457F18",
    x"13453201",
    x"1344E509",
    x"1344982E",
    x"13444B72",
    x"1343FED3",
    x"1343B253",
    x"134365F0",
    x"134319AB",
    x"1342CD84",
    x"1342817A",
    x"1342358F",
    x"1341E9C1",
    x"13419E10",
    x"1341527D",
    x"13410708",
    x"1340BBB0",
    x"13407075",
    x"13402558",
    x"133FDA58",
    x"133F8F75",
    x"133F44B0",
    x"133EFA07",
    x"133EAF7C",
    x"133E650E",
    x"133E1ABD",
    x"133DD089",
    x"133D8672",
    x"133D3C78",
    x"133CF29B",
    x"133CA8DB",
    x"133C5F37",
    x"133C15B0",
    x"133BCC46",
    x"133B82F9",
    x"133B39C8",
    x"133AF0B4",
    x"133AA7BC",
    x"133A5EE1",
    x"133A1622",
    x"1339CD7F",
    x"133984F9",
    x"13393C8F",
    x"1338F442",
    x"1338AC11",
    x"133863FB",
    x"13381C02",
    x"1337D426",
    x"13378C65",
    x"133744C0",
    x"1336FD37",
    x"1336B5CA",
    x"13366E79",
    x"13362744",
    x"1335E02A",
    x"1335992D",
    x"1335524B",
    x"13350B84",
    x"1334C4DA",
    x"13347E4A",
    x"133437D7",
    x"1333F17F",
    x"1333AB42",
    x"13336521",
    x"13331F1B",
    x"1332D931",
    x"13329361",
    x"13324DAE",
    x"13320815",
    x"1331C297",
    x"13317D35",
    x"133137ED",
    x"1330F2C1",
    x"1330ADB0",
    x"133068B9",
    x"133023DE",
    x"132FDF1D",
    x"132F9A78",
    x"132F55ED",
    x"132F117C",
    x"132ECD27",
    x"132E88EC",
    x"132E44CC",
    x"132E00C6",
    x"132DBCDB",
    x"132D790B",
    x"132D3555",
    x"132CF1B9",
    x"132CAE38",
    x"132C6AD1",
    x"132C2784",
    x"132BE452",
    x"132BA13A",
    x"132B5E3C",
    x"132B1B58",
    x"132AD88F",
    x"132A95DF",
    x"132A534A",
    x"132A10CE",
    x"1329CE6D",
    x"13298C25",
    x"132949F7",
    x"132907E3",
    x"1328C5E9",
    x"13288408",
    x"13284242",
    x"13280095",
    x"1327BF01",
    x"13277D87",
    x"13273C27",
    x"1326FAE0",
    x"1326B9B3",
    x"1326789F",
    x"132637A5",
    x"1325F6C4",
    x"1325B5FC",
    x"1325754E",
    x"132534B8",
    x"1324F43C",
    x"1324B3DA",
    x"13247390",
    x"1324335F",
    x"1323F348",
    x"1323B349",
    x"13237364",
    x"13233397",
    x"1322F3E3",
    x"1322B449",
    x"132274C6",
    x"1322355D",
    x"1321F60D",
    x"1321B6D5",
    x"132177B6",
    x"132138AF",
    x"1320F9C2",
    x"1320BAEC",
    x"13207C30",
    x"13203D8B",
    x"131FFF00",
    x"131FC08C",
    x"131F8231",
    x"131F43EE",
    x"131F05C4",
    x"131EC7B2",
    x"131E89B8",
    x"131E4BD6",
    x"131E0E0D",
    x"131DD05B",
    x"131D92C2",
    x"131D5541",
    x"131D17D7",
    x"131CDA86",
    x"131C9D4D",
    x"131C602B",
    x"131C2321",
    x"131BE630",
    x"131BA956",
    x"131B6C93",
    x"131B2FE9",
    x"131AF356",
    x"131AB6DB",
    x"131A7A77",
    x"131A3E2B",
    x"131A01F6",
    x"1319C5D9",
    x"131989D4",
    x"13194DE6",
    x"1319120F",
    x"1318D650",
    x"13189AA8",
    x"13185F17",
    x"1318239D",
    x"1317E83B",
    x"1317ACF0",
    x"131771BC",
    x"1317369F",
    x"1316FB99",
    x"1316C0AA",
    x"131685D3",
    x"13164B12",
    x"13161068",
    x"1315D5D5",
    x"13159B59",
    x"131560F4",
    x"131526A5",
    x"1314EC6D",
    x"1314B24C",
    x"13147842",
    x"13143E4E",
    x"13140471",
    x"1313CAAB",
    x"131390FB",
    x"13135762",
    x"13131DDF",
    x"1312E472",
    x"1312AB1C",
    x"131271DD",
    x"131238B3",
    x"1311FFA0",
    x"1311C6A4",
    x"13118DBD",
    x"131154ED",
    x"13111C33",
    x"1310E38F",
    x"1310AB01",
    x"13107289",
    x"13103A27",
    x"131001DC",
    x"130FC9A6",
    x"130F9186",
    x"130F597C",
    x"130F2188",
    x"130EE9AA",
    x"130EB1E2",
    x"130E7A2F",
    x"130E4292",
    x"130E0B0B",
    x"130DD39A",
    x"130D9C3E",
    x"130D64F8",
    x"130D2DC7",
    x"130CF6AC",
    x"130CBFA6",
    x"130C88B6",
    x"130C51DB",
    x"130C1B16",
    x"130BE466",
    x"130BADCC",
    x"130B7746",
    x"130B40D6",
    x"130B0A7C",
    x"130AD436",
    x"130A9E06",
    x"130A67EB",
    x"130A31E5",
    x"1309FBF4",
    x"1309C618",
    x"13099051",
    x"13095A9F",
    x"13092502",
    x"1308EF7A",
    x"1308BA07",
    x"130884A9",
    x"13084F5F",
    x"13081A2B",
    x"1307E50B",
    x"1307B000",
    x"13077B09",
    x"13074628",
    x"1307115B",
    x"1306DCA2",
    x"1306A7FE",
    x"1306736F",
    x"13063EF4",
    x"13060A8E",
    x"1305D63C",
    x"1305A1FE",
    x"13056DD5",
    x"130539C1",
    x"130505C0",
    x"1304D1D4",
    x"13049DFC",
    x"13046A39",
    x"13043689",
    x"130402EE",
    x"1303CF67",
    x"13039BF4",
    x"13036895",
    x"1303354A",
    x"13030213",
    x"1302CEF1",
    x"13029BE2",
    x"130268E7",
    x"13023600",
    x"1302032D",
    x"1301D06D",
    x"13019DC2",
    x"13016B2A",
    x"130138A6",
    x"13010636",
    x"1300D3D9",
    x"1300A190",
    x"13006F5B",
    x"13003D39",
    x"13000B2B",
    x"12FFB261",
    x"12FF4E93",
    x"12FEEAEC",
    x"12FE876B",
    x"12FE2412",
    x"12FDC0DF",
    x"12FD5DD3",
    x"12FCFAEE",
    x"12FC982F",
    x"12FC3597",
    x"12FBD325",
    x"12FB70DA",
    x"12FB0EB5",
    x"12FAACB6",
    x"12FA4ADE",
    x"12F9E92C",
    x"12F987A0",
    x"12F9263A",
    x"12F8C4FA",
    x"12F863E0",
    x"12F802EC",
    x"12F7A21E",
    x"12F74175",
    x"12F6E0F2",
    x"12F68095",
    x"12F6205E",
    x"12F5C04C",
    x"12F56060",
    x"12F50099",
    x"12F4A0F7",
    x"12F4417B",
    x"12F3E224",
    x"12F382F2",
    x"12F323E6",
    x"12F2C4FE",
    x"12F2663C",
    x"12F2079E",
    x"12F1A926",
    x"12F14AD2",
    x"12F0ECA3",
    x"12F08E99",
    x"12F030B4",
    x"12EFD2F3",
    x"12EF7557",
    x"12EF17E0",
    x"12EEBA8C",
    x"12EE5D5E",
    x"12EE0053",
    x"12EDA36E",
    x"12ED46AC",
    x"12ECEA0E",
    x"12EC8D95",
    x"12EC3140",
    x"12EBD50E",
    x"12EB7901",
    x"12EB1D18",
    x"12EAC152",
    x"12EA65B1",
    x"12EA0A33",
    x"12E9AED9",
    x"12E953A2",
    x"12E8F88F",
    x"12E89DA0",
    x"12E842D4",
    x"12E7E82C",
    x"12E78DA7",
    x"12E73345",
    x"12E6D907",
    x"12E67EEC",
    x"12E624F4",
    x"12E5CB1F",
    x"12E5716D",
    x"12E517DE",
    x"12E4BE72",
    x"12E46529",
    x"12E40C03",
    x"12E3B300",
    x"12E35A1F",
    x"12E30162",
    x"12E2A8C6",
    x"12E2504E",
    x"12E1F7F8",
    x"12E19FC4",
    x"12E147B3",
    x"12E0EFC4",
    x"12E097F7",
    x"12E0404D",
    x"12DFE8C5",
    x"12DF915F",
    x"12DF3A1C",
    x"12DEE2FA",
    x"12DE8BFA",
    x"12DE351C",
    x"12DDDE61",
    x"12DD87C7",
    x"12DD314F",
    x"12DCDAF8",
    x"12DC84C3",
    x"12DC2EB0",
    x"12DBD8BF",
    x"12DB82EF",
    x"12DB2D41",
    x"12DAD7B4",
    x"12DA8248",
    x"12DA2CFE",
    x"12D9D7D5",
    x"12D982CD",
    x"12D92DE7",
    x"12D8D921",
    x"12D8847D",
    x"12D82FFA",
    x"12D7DB98",
    x"12D78756",
    x"12D73336",
    x"12D6DF36",
    x"12D68B57",
    x"12D63799",
    x"12D5E3FC",
    x"12D5907F",
    x"12D53D23",
    x"12D4E9E7",
    x"12D496CC",
    x"12D443D2",
    x"12D3F0F7",
    x"12D39E3D",
    x"12D34BA4",
    x"12D2F92A",
    x"12D2A6D1",
    x"12D25498",
    x"12D2027F",
    x"12D1B086",
    x"12D15EAD",
    x"12D10CF4",
    x"12D0BB5B",
    x"12D069E2",
    x"12D01888",
    x"12CFC74E",
    x"12CF7634",
    x"12CF253A",
    x"12CED45F",
    x"12CE83A4",
    x"12CE3308",
    x"12CDE28C",
    x"12CD922F",
    x"12CD41F2",
    x"12CCF1D4",
    x"12CCA1D5",
    x"12CC51F5",
    x"12CC0235",
    x"12CBB294",
    x"12CB6312",
    x"12CB13AE",
    x"12CAC46A",
    x"12CA7545",
    x"12CA263E",
    x"12C9D757",
    x"12C9888E",
    x"12C939E4",
    x"12C8EB59",
    x"12C89CEC",
    x"12C84E9E",
    x"12C8006F",
    x"12C7B25E",
    x"12C7646C",
    x"12C71698",
    x"12C6C8E2",
    x"12C67B4B",
    x"12C62DD2",
    x"12C5E077",
    x"12C5933A",
    x"12C5461C",
    x"12C4F91B",
    x"12C4AC39",
    x"12C45F75",
    x"12C412CF",
    x"12C3C646",
    x"12C379DC",
    x"12C32D8F",
    x"12C2E160",
    x"12C2954F",
    x"12C2495B",
    x"12C1FD86",
    x"12C1B1CD",
    x"12C16633",
    x"12C11AB5",
    x"12C0CF56",
    x"12C08413",
    x"12C038EF",
    x"12BFEDE7",
    x"12BFA2FD",
    x"12BF5830",
    x"12BF0D80",
    x"12BEC2ED",
    x"12BE7877",
    x"12BE2E1F",
    x"12BDE3E3",
    x"12BD99C5",
    x"12BD4FC3",
    x"12BD05DF",
    x"12BCBC17",
    x"12BC726C",
    x"12BC28DD",
    x"12BBDF6C",
    x"12BB9617",
    x"12BB4CDE",
    x"12BB03C3",
    x"12BABAC3",
    x"12BA71E1",
    x"12BA291A",
    x"12B9E071",
    x"12B997E3",
    x"12B94F72",
    x"12B9071D",
    x"12B8BEE4",
    x"12B876C8",
    x"12B82EC7",
    x"12B7E6E3",
    x"12B79F1B",
    x"12B7576F",
    x"12B70FDF",
    x"12B6C86B",
    x"12B68112",
    x"12B639D6",
    x"12B5F2B5",
    x"12B5ABB0",
    x"12B564C7",
    x"12B51DF9",
    x"12B4D747",
    x"12B490B1",
    x"12B44A36",
    x"12B403D7",
    x"12B3BD93",
    x"12B3776B",
    x"12B3315E",
    x"12B2EB6C",
    x"12B2A596",
    x"12B25FDB",
    x"12B21A3B",
    x"12B1D4B7",
    x"12B18F4D",
    x"12B149FF",
    x"12B104CB",
    x"12B0BFB3",
    x"12B07AB5",
    x"12B035D3",
    x"12AFF10B",
    x"12AFAC5F",
    x"12AF67CD",
    x"12AF2355",
    x"12AEDEF9",
    x"12AE9AB7",
    x"12AE5690",
    x"12AE1284",
    x"12ADCE92",
    x"12AD8ABA",
    x"12AD46FD",
    x"12AD035B",
    x"12ACBFD3",
    x"12AC7C65",
    x"12AC3911",
    x"12ABF5D8",
    x"12ABB2B9",
    x"12AB6FB5",
    x"12AB2CCA",
    x"12AAE9FA",
    x"12AAA743",
    x"12AA64A7",
    x"12AA2225",
    x"12A9DFBC",
    x"12A99D6E",
    x"12A95B39",
    x"12A9191F",
    x"12A8D71E",
    x"12A89536",
    x"12A85369",
    x"12A811B5",
    x"12A7D01B",
    x"12A78E9B",
    x"12A74D34",
    x"12A70BE6",
    x"12A6CAB2",
    x"12A68998",
    x"12A64897",
    x"12A607AF",
    x"12A5C6E1",
    x"12A5862C",
    x"12A54590",
    x"12A5050E",
    x"12A4C4A4",
    x"12A48454",
    x"12A4441D",
    x"12A403FF",
    x"12A3C3FA",
    x"12A3840E",
    x"12A3443A",
    x"12A30480",
    x"12A2C4DF",
    x"12A28556",
    x"12A245E7",
    x"12A20690",
    x"12A1C752",
    x"12A1882C",
    x"12A1491F",
    x"12A10A2B",
    x"12A0CB4F",
    x"12A08C8C",
    x"12A04DE1",
    x"12A00F4F",
    x"129FD0D5",
    x"129F9274",
    x"129F542B",
    x"129F15FA",
    x"129ED7E2",
    x"129E99E2",
    x"129E5BFA",
    x"129E1E2A",
    x"129DE072",
    x"129DA2D2",
    x"129D654B",
    x"129D27DB",
    x"129CEA84",
    x"129CAD44",
    x"129C701C",
    x"129C330C",
    x"129BF614",
    x"129BB934",
    x"129B7C6C",
    x"129B3FBB",
    x"129B0322",
    x"129AC6A0",
    x"129A8A37",
    x"129A4DE4",
    x"129A11AA",
    x"1299D587",
    x"1299997B",
    x"12995D87",
    x"129921AA",
    x"1298E5E4",
    x"1298AA36",
    x"12986E9F",
    x"12983320",
    x"1297F7B7",
    x"1297BC66",
    x"1297812C",
    x"12974609",
    x"12970AFE",
    x"1296D009",
    x"1296952B",
    x"12965A64",
    x"12961FB4",
    x"1295E51B",
    x"1295AA99",
    x"1295702E",
    x"129535DA",
    x"1294FB9C",
    x"1294C175",
    x"12948765",
    x"12944D6B",
    x"12941388",
    x"1293D9BC",
    x"1293A006",
    x"12936667",
    x"12932CDE",
    x"1292F36C",
    x"1292BA10",
    x"129280CB",
    x"1292479B",
    x"12920E83",
    x"1291D580",
    x"12919C94",
    x"129163BE",
    x"12912AFE",
    x"1290F254",
    x"1290B9C1",
    x"12908143",
    x"129048DC",
    x"1290108A",
    x"128FD84F",
    x"128FA029",
    x"128F681A",
    x"128F3020",
    x"128EF83C",
    x"128EC06E",
    x"128E88B6",
    x"128E5113",
    x"128E1986",
    x"128DE20F",
    x"128DAAAE",
    x"128D7362",
    x"128D3C2B",
    x"128D050B",
    x"128CCE00",
    x"128C970A",
    x"128C602A",
    x"128C295F",
    x"128BF2A9",
    x"128BBC09",
    x"128B857E",
    x"128B4F09",
    x"128B18A9",
    x"128AE25D",
    x"128AAC28",
    x"128A7607",
    x"128A3FFB",
    x"128A0A05",
    x"1289D424",
    x"12899E57",
    x"128968A0",
    x"128932FD",
    x"1288FD70",
    x"1288C7F7",
    x"12889294",
    x"12885D45",
    x"1288280B",
    x"1287F2E6",
    x"1287BDD5",
    x"128788D9",
    x"128753F2",
    x"12871F20",
    x"1286EA62",
    x"1286B5B9",
    x"12868124",
    x"12864CA4",
    x"12861838",
    x"1285E3E1",
    x"1285AF9E",
    x"12857B70",
    x"12854756",
    x"12851350",
    x"1284DF5E",
    x"1284AB81",
    x"128477B8",
    x"12844404",
    x"12841063",
    x"1283DCD7",
    x"1283A95F",
    x"128375FB",
    x"128342AB",
    x"12830F6F",
    x"1282DC47",
    x"1282A932",
    x"12827632",
    x"12824346",
    x"1282106E",
    x"1281DDA9",
    x"1281AAF9",
    x"1281785C",
    x"128145D3",
    x"1281135D",
    x"1280E0FB",
    x"1280AEAD",
    x"12807C73",
    x"12804A4C",
    x"12801839",
    x"127FCC72",
    x"127F689A",
    x"127F04E9",
    x"127EA15E",
    x"127E3DFA",
    x"127DDABE",
    x"127D77A8",
    x"127D14B8",
    x"127CB1EF",
    x"127C4F4D",
    x"127BECD1",
    x"127B8A7C",
    x"127B284D",
    x"127AC645",
    x"127A6462",
    x"127A02A6",
    x"1279A110",
    x"12793FA0",
    x"1278DE56",
    x"12787D33",
    x"12781C35",
    x"1277BB5D",
    x"12775AAA",
    x"1276FA1E",
    x"127699B7",
    x"12763976",
    x"1275D95A",
    x"12757964",
    x"12751993",
    x"1274B9E8",
    x"12745A62",
    x"1273FB01",
    x"12739BC6",
    x"12733CAF",
    x"1272DDBE",
    x"12727EF2",
    x"1272204B",
    x"1271C1C9",
    x"1271636C",
    x"12710533",
    x"1270A720",
    x"12704931",
    x"126FEB66",
    x"126F8DC1",
    x"126F3040",
    x"126ED2E3",
    x"126E75AB",
    x"126E1897",
    x"126DBBA8",
    x"126D5EDC",
    x"126D0235",
    x"126CA5B3",
    x"126C4954",
    x"126BED19",
    x"126B9103",
    x"126B3510",
    x"126AD941",
    x"126A7D96",
    x"126A220F",
    x"1269C6AC",
    x"12696B6C",
    x"12691050",
    x"1268B557",
    x"12685A82",
    x"1267FFD0",
    x"1267A542",
    x"12674AD7",
    x"1266F090",
    x"1266966B",
    x"12663C6A",
    x"1265E28C",
    x"126588D1",
    x"12652F39",
    x"1264D5C4",
    x"12647C72",
    x"12642343",
    x"1263CA37",
    x"1263714D",
    x"12631886",
    x"1262BFE2",
    x"12626760",
    x"12620F01",
    x"1261B6C4",
    x"12615EAA",
    x"126106B2",
    x"1260AEDD",
    x"1260572A",
    x"125FFF99",
    x"125FA82A",
    x"125F50DD",
    x"125EF9B3",
    x"125EA2AA",
    x"125E4BC4",
    x"125DF4FF",
    x"125D9E5C",
    x"125D47DB",
    x"125CF17C",
    x"125C9B3F",
    x"125C4523",
    x"125BEF29",
    x"125B9950",
    x"125B4399",
    x"125AEE03",
    x"125A988F",
    x"125A433C",
    x"1259EE0A",
    x"125998FA",
    x"1259440B",
    x"1258EF3D",
    x"12589A90",
    x"12584604",
    x"1257F199",
    x"12579D4F",
    x"12574926",
    x"1256F51E",
    x"1256A137",
    x"12564D70",
    x"1255F9CA",
    x"1255A645",
    x"125552E0",
    x"1254FF9C",
    x"1254AC79",
    x"12545976",
    x"12540693",
    x"1253B3D0",
    x"1253612E",
    x"12530EAC",
    x"1252BC4B",
    x"12526A09",
    x"125217E8",
    x"1251C5E7",
    x"12517405",
    x"12512244",
    x"1250D0A3",
    x"12507F21",
    x"12502DBF",
    x"124FDC7D",
    x"124F8B5B",
    x"124F3A58",
    x"124EE975",
    x"124E98B2",
    x"124E480E",
    x"124DF78A",
    x"124DA725",
    x"124D56DF",
    x"124D06B9",
    x"124CB6B2",
    x"124C66CA",
    x"124C1701",
    x"124BC758",
    x"124B77CE",
    x"124B2862",
    x"124AD916",
    x"124A89E9",
    x"124A3ADA",
    x"1249EBEB",
    x"12499D1A",
    x"12494E68",
    x"1248FFD5",
    x"1248B160",
    x"1248630A",
    x"124814D3",
    x"1247C6BA",
    x"124778BF",
    x"12472AE4",
    x"1246DD26",
    x"12468F87",
    x"12464206",
    x"1245F4A3",
    x"1245A75F",
    x"12455A38",
    x"12450D30",
    x"1244C046",
    x"1244737A",
    x"124426CC",
    x"1243DA3C",
    x"12438DC9",
    x"12434175",
    x"1242F53E",
    x"1242A925",
    x"12425D2A",
    x"1242114C",
    x"1241C58C",
    x"124179EA",
    x"12412E65",
    x"1240E2FE",
    x"124097B4",
    x"12404C87",
    x"12400178",
    x"123FB686",
    x"123F6BB1",
    x"123F20FA",
    x"123ED660",
    x"123E8BE2",
    x"123E4182",
    x"123DF73F",
    x"123DAD19",
    x"123D6310",
    x"123D1924",
    x"123CCF54",
    x"123C85A2",
    x"123C3C0C",
    x"123BF293",
    x"123BA936",
    x"123B5FF7",
    x"123B16D3",
    x"123ACDCD",
    x"123A84E3",
    x"123A3C15",
    x"1239F364",
    x"1239AACF",
    x"12396256",
    x"123919FA",
    x"1238D1BA",
    x"12388996",
    x"1238418E",
    x"1237F9A3",
    x"1237B1D3",
    x"12376A20",
    x"12372288",
    x"1236DB0D",
    x"123693AD",
    x"12364C6A",
    x"12360542",
    x"1235BE35",
    x"12357745",
    x"12353070",
    x"1234E9B7",
    x"1234A31A",
    x"12345C98",
    x"12341631",
    x"1233CFE6",
    x"123389B7",
    x"123343A3",
    x"1232FDAA",
    x"1232B7CD",
    x"1232720A",
    x"12322C63",
    x"1231E6D8",
    x"1231A167",
    x"12315C12",
    x"123116D7",
    x"1230D1B8",
    x"12308CB3",
    x"123047CA",
    x"123002FB",
    x"122FBE47",
    x"122F79AF",
    x"122F3530",
    x"122EF0CD",
    x"122EAC84",
    x"122E6856",
    x"122E2443",
    x"122DE04A",
    x"122D9C6B",
    x"122D58A8",
    x"122D14FE",
    x"122CD16F",
    x"122C8DFB",
    x"122C4AA0",
    x"122C0760",
    x"122BC43A",
    x"122B812F",
    x"122B3E3E",
    x"122AFB66",
    x"122AB8A9",
    x"122A7606",
    x"122A337D",
    x"1229F10E",
    x"1229AEB9",
    x"12296C7D",
    x"12292A5C",
    x"1228E854",
    x"1228A666",
    x"12286492",
    x"122822D8",
    x"1227E137",
    x"12279FB0",
    x"12275E42",
    x"12271CEE",
    x"1226DBB4",
    x"12269A92",
    x"1226598B",
    x"1226189C",
    x"1225D7C8",
    x"1225970C",
    x"12255669",
    x"122515E0",
    x"1224D570",
    x"1224951A",
    x"122454DC",
    x"122414B7",
    x"1223D4AC",
    x"122394B9",
    x"122354DF",
    x"1223151F",
    x"1222D577",
    x"122295E8",
    x"12225672",
    x"12221714",
    x"1221D7D0",
    x"122198A4",
    x"12215991",
    x"12211A96",
    x"1220DBB4",
    x"12209CEA",
    x"12205E39",
    x"12201FA1",
    x"121FE120",
    x"121FA2B9",
    x"121F6469",
    x"121F2632",
    x"121EE813",
    x"121EAA0D",
    x"121E6C1F",
    x"121E2E48",
    x"121DF08A",
    x"121DB2E4",
    x"121D7557",
    x"121D37E1",
    x"121CFA83",
    x"121CBD3D",
    x"121C800F",
    x"121C42F9",
    x"121C05FB",
    x"121BC914",
    x"121B8C46",
    x"121B4F8F",
    x"121B12F0",
    x"121AD668",
    x"121A99F8",
    x"121A5DA0",
    x"121A215F",
    x"1219E536",
    x"1219A924",
    x"12196D29",
    x"12193146",
    x"1218F57B",
    x"1218B9C7",
    x"12187E2A",
    x"121842A4",
    x"12180736",
    x"1217CBDE",
    x"1217909E",
    x"12175575",
    x"12171A64",
    x"1216DF69",
    x"1216A485",
    x"121669B8",
    x"12162F02",
    x"1215F464",
    x"1215B9DC",
    x"12157F6A",
    x"12154510",
    x"12150ACC",
    x"1214D0A0",
    x"12149689",
    x"12145C8A",
    x"121422A1",
    x"1213E8CF",
    x"1213AF13",
    x"1213756E",
    x"12133BDF",
    x"12130267",
    x"1212C906",
    x"12128FBA",
    x"12125685",
    x"12121D67",
    x"1211E45E",
    x"1211AB6C",
    x"12117290",
    x"121139CB",
    x"1211011B",
    x"1210C882",
    x"12108FFE",
    x"12105791",
    x"12101F3A",
    x"120FE6F9",
    x"120FAECE",
    x"120F76B8",
    x"120F3EB9",
    x"120F06CF",
    x"120ECEFC",
    x"120E973E",
    x"120E5F95",
    x"120E2803",
    x"120DF086",
    x"120DB91F",
    x"120D81CD",
    x"120D4A92",
    x"120D136B",
    x"120CDC5A",
    x"120CA55F",
    x"120C6E79",
    x"120C37A9",
    x"120C00EE",
    x"120BCA48",
    x"120B93B8",
    x"120B5D3D",
    x"120B26D7",
    x"120AF086",
    x"120ABA4B",
    x"120A8425",
    x"120A4E14",
    x"120A1818",
    x"1209E231",
    x"1209AC5F",
    x"120976A2",
    x"120940FA",
    x"12090B67",
    x"1208D5E9",
    x"1208A080",
    x"12086B2C",
    x"120835EC",
    x"120800C2",
    x"1207CBAC",
    x"120796AB",
    x"120761BE",
    x"12072CE6",
    x"1206F823",
    x"1206C374",
    x"12068EDA",
    x"12065A55",
    x"120625E4",
    x"1205F187",
    x"1205BD3F",
    x"1205890B",
    x"120554EC",
    x"120520E1",
    x"1204ECEA",
    x"1204B908",
    x"1204853A",
    x"12045180",
    x"12041DDA",
    x"1203EA48",
    x"1203B6CB",
    x"12038362",
    x"1203500C",
    x"12031CCB",
    x"1202E99E",
    x"1202B685",
    x"1202837F",
    x"1202508E",
    x"12021DB0",
    x"1201EAE7",
    x"1201B831",
    x"1201858F",
    x"12015300",
    x"12012086",
    x"1200EE1F",
    x"1200BBCC",
    x"1200898C",
    x"12005760",
    x"12002548",
    x"11FFE686",
    x"11FF82A4",
    x"11FF1EE8",
    x"11FEBB54",
    x"11FE57E6",
    x"11FDF49F",
    x"11FD917F",
    x"11FD2E85",
    x"11FCCBB2",
    x"11FC6906",
    x"11FC0680",
    x"11FBA421",
    x"11FB41E8",
    x"11FADFD6",
    x"11FA7DE9",
    x"11FA1C23",
    x"11F9BA83",
    x"11F95909",
    x"11F8F7B6",
    x"11F89688",
    x"11F83580",
    x"11F7D49E",
    x"11F773E2",
    x"11F7134B",
    x"11F6B2DB",
    x"11F65290",
    x"11F5F26A",
    x"11F5926A",
    x"11F53290",
    x"11F4D2DB",
    x"11F4734B",
    x"11F413E1",
    x"11F3B49C",
    x"11F3557C",
    x"11F2F681",
    x"11F297AB",
    x"11F238FA",
    x"11F1DA6E",
    x"11F17C08",
    x"11F11DC6",
    x"11F0BFA8",
    x"11F061B0",
    x"11F003DC",
    x"11EFA62D",
    x"11EF48A2",
    x"11EEEB3C",
    x"11EE8DFA",
    x"11EE30DD",
    x"11EDD3E4",
    x"11ED7710",
    x"11ED1A5F",
    x"11ECBDD3",
    x"11EC616B",
    x"11EC0527",
    x"11EBA907",
    x"11EB4D0B",
    x"11EAF133",
    x"11EA957E",
    x"11EA39EE",
    x"11E9DE81",
    x"11E98338",
    x"11E92812",
    x"11E8CD11",
    x"11E87232",
    x"11E81777",
    x"11E7BCE0",
    x"11E7626C",
    x"11E7081B",
    x"11E6ADED",
    x"11E653E3",
    x"11E5F9FC",
    x"11E5A038",
    x"11E54697",
    x"11E4ED19",
    x"11E493BD",
    x"11E43A85",
    x"11E3E170",
    x"11E3887D",
    x"11E32FAD",
    x"11E2D700",
    x"11E27E75",
    x"11E2260D",
    x"11E1CDC7",
    x"11E175A4",
    x"11E11DA3",
    x"11E0C5C5",
    x"11E06E09",
    x"11E0166F",
    x"11DFBEF7",
    x"11DF67A2",
    x"11DF106E",
    x"11DEB95D",
    x"11DE626D",
    x"11DE0BA0",
    x"11DDB4F4",
    x"11DD5E6B",
    x"11DD0803",
    x"11DCB1BC",
    x"11DC5B98",
    x"11DC0595",
    x"11DBAFB3",
    x"11DB59F3",
    x"11DB0455",
    x"11DAAED8",
    x"11DA597C",
    x"11DA0442",
    x"11D9AF29",
    x"11D95A31",
    x"11D9055B",
    x"11D8B0A5",
    x"11D85C11",
    x"11D8079D",
    x"11D7B34B",
    x"11D75F19",
    x"11D70B08",
    x"11D6B718",
    x"11D66349",
    x"11D60F9B",
    x"11D5BC0D",
    x"11D568A0",
    x"11D51553",
    x"11D4C227",
    x"11D46F1C",
    x"11D41C30",
    x"11D3C966",
    x"11D376BB",
    x"11D32431",
    x"11D2D1C7",
    x"11D27F7D",
    x"11D22D53",
    x"11D1DB49",
    x"11D18960",
    x"11D13796",
    x"11D0E5EC",
    x"11D09462",
    x"11D042F8",
    x"11CFF1AE",
    x"11CFA084",
    x"11CF4F79",
    x"11CEFE8D",
    x"11CEADC2",
    x"11CE5D16",
    x"11CE0C89",
    x"11CDBC1C",
    x"11CD6BCE",
    x"11CD1BA0",
    x"11CCCB91",
    x"11CC7BA1",
    x"11CC2BD0",
    x"11CBDC1E",
    x"11CB8C8C",
    x"11CB3D19",
    x"11CAEDC4",
    x"11CA9E8F",
    x"11CA4F78",
    x"11CA0081",
    x"11C9B1A8",
    x"11C962EE",
    x"11C91453",
    x"11C8C5D6",
    x"11C87778",
    x"11C82939",
    x"11C7DB18",
    x"11C78D15",
    x"11C73F32",
    x"11C6F16C",
    x"11C6A3C5",
    x"11C6563C",
    x"11C608D2",
    x"11C5BB85",
    x"11C56E57",
    x"11C52147",
    x"11C4D455",
    x"11C48781",
    x"11C43ACB",
    x"11C3EE33",
    x"11C3A1B9",
    x"11C3555D",
    x"11C3091E",
    x"11C2BCFE",
    x"11C270FB",
    x"11C22515",
    x"11C1D94E",
    x"11C18DA4",
    x"11C14217",
    x"11C0F6A8",
    x"11C0AB56",
    x"11C06022",
    x"11C0150B",
    x"11BFCA12",
    x"11BF7F35",
    x"11BF3476",
    x"11BEE9D4",
    x"11BE9F50",
    x"11BE54E8",
    x"11BE0A9D",
    x"11BDC070",
    x"11BD765F",
    x"11BD2C6B",
    x"11BCE294",
    x"11BC98DA",
    x"11BC4F3D",
    x"11BC05BC",
    x"11BBBC58",
    x"11BB7311",
    x"11BB29E6",
    x"11BAE0D8",
    x"11BA97E7",
    x"11BA4F11",
    x"11BA0659",
    x"11B9BDBD",
    x"11B9753D",
    x"11B92CD9",
    x"11B8E491",
    x"11B89C66",
    x"11B85457",
    x"11B80C64",
    x"11B7C48E",
    x"11B77CD3",
    x"11B73534",
    x"11B6EDB1",
    x"11B6A64A",
    x"11B65EFF",
    x"11B617D0",
    x"11B5D0BD",
    x"11B589C5",
    x"11B542E9",
    x"11B4FC29",
    x"11B4B584",
    x"11B46EFB",
    x"11B4288D",
    x"11B3E23B",
    x"11B39C05",
    x"11B355E9",
    x"11B30FE9",
    x"11B2CA05",
    x"11B2843C",
    x"11B23E8E",
    x"11B1F8FB",
    x"11B1B383",
    x"11B16E26",
    x"11B128E5",
    x"11B0E3BE",
    x"11B09EB3",
    x"11B059C3",
    x"11B014ED",
    x"11AFD032",
    x"11AF8B92",
    x"11AF470D",
    x"11AF02A3",
    x"11AEBE53",
    x"11AE7A1E",
    x"11AE3604",
    x"11ADF204",
    x"11ADAE1F",
    x"11AD6A54",
    x"11AD26A3",
    x"11ACE30E",
    x"11AC9F92",
    x"11AC5C31",
    x"11AC18EA",
    x"11ABD5BD",
    x"11AB92AB",
    x"11AB4FB3",
    x"11AB0CD5",
    x"11AACA11",
    x"11AA8767",
    x"11AA44D7",
    x"11AA0261",
    x"11A9C005",
    x"11A97DC3",
    x"11A93B9B",
    x"11A8F98C",
    x"11A8B798",
    x"11A875BD",
    x"11A833FC",
    x"11A7F254",
    x"11A7B0C7",
    x"11A76F52",
    x"11A72DF8",
    x"11A6ECB6",
    x"11A6AB8F",
    x"11A66A80",
    x"11A6298B",
    x"11A5E8B0",
    x"11A5A7EE",
    x"11A56745",
    x"11A526B5",
    x"11A4E63E",
    x"11A4A5E1",
    x"11A4659D",
    x"11A42572",
    x"11A3E55F",
    x"11A3A566",
    x"11A36586",
    x"11A325BF",
    x"11A2E611",
    x"11A2A67B",
    x"11A266FF",
    x"11A2279B",
    x"11A1E850",
    x"11A1A91D",
    x"11A16A04",
    x"11A12B02",
    x"11A0EC1A",
    x"11A0AD4A",
    x"11A06E93",
    x"11A02FF4",
    x"119FF16D",
    x"119FB2FF",
    x"119F74A9",
    x"119F366C",
    x"119EF847",
    x"119EBA3A",
    x"119E7C45",
    x"119E3E69",
    x"119E00A4",
    x"119DC2F8",
    x"119D8564",
    x"119D47E8",
    x"119D0A84",
    x"119CCD38",
    x"119C9004",
    x"119C52E7",
    x"119C15E3",
    x"119BD8F6",
    x"119B9C21",
    x"119B5F64",
    x"119B22BF",
    x"119AE631",
    x"119AA9BB",
    x"119A6D5C",
    x"119A3115",
    x"1199F4E6",
    x"1199B8CE",
    x"11997CCE",
    x"119940E5",
    x"11990513",
    x"1198C959",
    x"11988DB6",
    x"1198522A",
    x"119816B5",
    x"1197DB58",
    x"1197A012",
    x"119764E3",
    x"119729CB",
    x"1196EECA",
    x"1196B3E1",
    x"1196790E",
    x"11963E52",
    x"119603AD",
    x"1195C91F",
    x"11958EA8",
    x"11955448",
    x"119519FE",
    x"1194DFCB",
    x"1194A5AF",
    x"11946BAA",
    x"119431BB",
    x"1193F7E3",
    x"1193BE22",
    x"11938477",
    x"11934AE2",
    x"11931164",
    x"1192D7FC",
    x"11929EAB",
    x"11926570",
    x"11922C4C",
    x"1191F33E",
    x"1191BA46",
    x"11918164",
    x"11914899",
    x"11910FE4",
    x"1190D744",
    x"11909EBB",
    x"11906648",
    x"11902DEB",
    x"118FF5A5",
    x"118FBD74",
    x"118F8559",
    x"118F4D53",
    x"118F1564",
    x"118EDD8B",
    x"118EA5C7",
    x"118E6E19",
    x"118E3681",
    x"118DFEFF",
    x"118DC792",
    x"118D903B",
    x"118D58F9",
    x"118D21CD",
    x"118CEAB7",
    x"118CB3B6",
    x"118C7CCA",
    x"118C45F4",
    x"118C0F34",
    x"118BD888",
    x"118BA1F2",
    x"118B6B72",
    x"118B3506",
    x"118AFEB0",
    x"118AC86F",
    x"118A9244",
    x"118A5C2D",
    x"118A262C",
    x"1189F03F",
    x"1189BA68",
    x"118984A6",
    x"11894EF8",
    x"11891960",
    x"1188E3DD",
    x"1188AE6E",
    x"11887914",
    x"118843CF",
    x"11880E9F",
    x"1187D984",
    x"1187A47D",
    x"11876F8B",
    x"11873AAE",
    x"118705E6",
    x"1186D132",
    x"11869C92",
    x"11866807",
    x"11863391",
    x"1185FF2F",
    x"1185CAE1",
    x"118596A8",
    x"11856284",
    x"11852E73",
    x"1184FA77",
    x"1184C690",
    x"118492BC",
    x"11845EFD",
    x"11842B52",
    x"1183F7BB",
    x"1183C439",
    x"118390CA",
    x"11835D6F",
    x"11832A29",
    x"1182F6F6",
    x"1182C3D8",
    x"118290CD",
    x"11825DD7",
    x"11822AF4",
    x"1181F825",
    x"1181C56A",
    x"118192C3",
    x"11816030",
    x"11812DB0",
    x"1180FB44",
    x"1180C8EC",
    x"118096A7",
    x"11806476",
    x"11803258",
    x"1180004F",
    x"117F9CB0",
    x"117F38EB",
    x"117ED54C",
    x"117E71D4",
    x"117E0E83",
    x"117DAB59",
    x"117D4855",
    x"117CE578",
    x"117C82C2",
    x"117C2032",
    x"117BBDC9",
    x"117B5B86",
    x"117AF969",
    x"117A9773",
    x"117A35A3",
    x"1179D3F9",
    x"11797275",
    x"11791117",
    x"1178AFE0",
    x"11784ECE",
    x"1177EDE2",
    x"11778D1C",
    x"11772C7C",
    x"1176CC01",
    x"11766BAC",
    x"11760B7D",
    x"1175AB73",
    x"11754B8F",
    x"1174EBD0",
    x"11748C37",
    x"11742CC3",
    x"1173CD74",
    x"11736E4A",
    x"11730F46",
    x"1172B066",
    x"117251AC",
    x"1171F317",
    x"117194A6",
    x"1171365A",
    x"1170D834",
    x"11707A31",
    x"11701C54",
    x"116FBE9B",
    x"116F6107",
    x"116F0398",
    x"116EA64C",
    x"116E4926",
    x"116DEC23",
    x"116D8F45",
    x"116D328B",
    x"116CD5F6",
    x"116C7984",
    x"116C1D37",
    x"116BC10D",
    x"116B6508",
    x"116B0926",
    x"116AAD69",
    x"116A51CF",
    x"1169F659",
    x"11699B06",
    x"11693FD8",
    x"1168E4CC",
    x"116889E5",
    x"11682F21",
    x"1167D480",
    x"11677A03",
    x"11671FA9",
    x"1166C572",
    x"11666B5E",
    x"1166116E",
    x"1165B7A1",
    x"11655DF6",
    x"1165046F",
    x"1164AB0B",
    x"116451CA",
    x"1163F8AB",
    x"11639FAF",
    x"116346D6",
    x"1162EE20",
    x"1162958C",
    x"11623D1B",
    x"1161E4CC",
    x"11618CA0",
    x"11613497",
    x"1160DCAF",
    x"116084EA",
    x"11602D47",
    x"115FD5C7",
    x"115F7E68",
    x"115F272C",
    x"115ED012",
    x"115E7919",
    x"115E2243",
    x"115DCB8F",
    x"115D74FC",
    x"115D1E8B",
    x"115CC83C",
    x"115C720F",
    x"115C1C03",
    x"115BC619",
    x"115B7050",
    x"115B1AA9",
    x"115AC523",
    x"115A6FBF",
    x"115A1A7C",
    x"1159C55A",
    x"1159705A",
    x"11591B7B",
    x"1158C6BC",
    x"1158721F",
    x"11581DA3",
    x"1157C948",
    x"1157750E",
    x"115720F5",
    x"1156CCFC",
    x"11567925",
    x"1156256E",
    x"1155D1D7",
    x"11557E62",
    x"11552B0D",
    x"1154D7D8",
    x"115484C4",
    x"115431D0",
    x"1153DEFD",
    x"11538C4A",
    x"115339B7",
    x"1152E745",
    x"115294F3",
    x"115242C1",
    x"1151F0AE",
    x"11519EBC",
    x"11514CEA",
    x"1150FB38",
    x"1150A9A6",
    x"11505834",
    x"115006E1",
    x"114FB5AE",
    x"114F649B",
    x"114F13A8",
    x"114EC2D4",
    x"114E7220",
    x"114E218B",
    x"114DD115",
    x"114D80BF",
    x"114D3089",
    x"114CE071",
    x"114C9079",
    x"114C40A1",
    x"114BF0E7",
    x"114BA14C",
    x"114B51D1",
    x"114B0274",
    x"114AB337",
    x"114A6418",
    x"114A1519",
    x"1149C638",
    x"11497776",
    x"114928D3",
    x"1148DA4E",
    x"11488BE8",
    x"11483DA1",
    x"1147EF78",
    x"1147A16E",
    x"11475382",
    x"114705B4",
    x"1146B805",
    x"11466A74",
    x"11461D02",
    x"1145CFAE",
    x"11458278",
    x"11453560",
    x"1144E866",
    x"11449B8A",
    x"11444ECD",
    x"1144022D",
    x"1143B5AB",
    x"11436947",
    x"11431D01",
    x"1142D0D8",
    x"114284CD",
    x"114238E0",
    x"1141ED11",
    x"1141A15F",
    x"114155CB",
    x"11410A54",
    x"1140BEFB",
    x"114073BF",
    x"114028A0",
    x"113FDD9F",
    x"113F92BB",
    x"113F47F4",
    x"113EFD4B",
    x"113EB2BF",
    x"113E684F",
    x"113E1DFD",
    x"113DD3C8",
    x"113D89B0",
    x"113D3FB4",
    x"113CF5D6",
    x"113CAC14",
    x"113C626F",
    x"113C18E7",
    x"113BCF7C",
    x"113B862D",
    x"113B3CFB",
    x"113AF3E5",
    x"113AAAEC",
    x"113A6210",
    x"113A1950",
    x"1139D0AC",
    x"11398825",
    x"11393FBA",
    x"1138F76B",
    x"1138AF38",
    x"11386722",
    x"11381F28",
    x"1137D74A",
    x"11378F88",
    x"113747E2",
    x"11370057",
    x"1136B8E9",
    x"11367197",
    x"11362A61",
    x"1135E346",
    x"11359C47",
    x"11355564",
    x"11350E9C",
    x"1134C7F0",
    x"11348160",
    x"11343AEB",
    x"1133F492",
    x"1133AE54",
    x"11336832",
    x"1133222B",
    x"1132DC3F",
    x"1132966F",
    x"113250BA",
    x"11320B20",
    x"1131C5A1",
    x"1131803D",
    x"11313AF5",
    x"1130F5C7",
    x"1130B0B5",
    x"11306BBD",
    x"113026E0",
    x"112FE21F",
    x"112F9D78",
    x"112F58EC",
    x"112F147A",
    x"112ED024",
    x"112E8BE8",
    x"112E47C6",
    x"112E03C0",
    x"112DBFD3",
    x"112D7C02",
    x"112D384A",
    x"112CF4AE",
    x"112CB12B",
    x"112C6DC3",
    x"112C2A76",
    x"112BE742",
    x"112BA429",
    x"112B612A",
    x"112B1E45",
    x"112ADB7A",
    x"112A98C9",
    x"112A5633",
    x"112A13B6",
    x"1129D153",
    x"11298F0B",
    x"11294CDC",
    x"11290AC6",
    x"1128C8CB",
    x"112886EA",
    x"11284522",
    x"11280374",
    x"1127C1DF",
    x"11278064",
    x"11273F03",
    x"1126FDBB",
    x"1126BC8C",
    x"11267B78",
    x"11263A7C",
    x"1125F99A",
    x"1125B8D1",
    x"11257821",
    x"1125378B",
    x"1124F70E",
    x"1124B6AA",
    x"1124765F",
    x"1124362E",
    x"1123F615",
    x"1123B615",
    x"1123762F",
    x"11233661",
    x"1122F6AC",
    x"1122B710",
    x"1122778D",
    x"11223823",
    x"1121F8D1",
    x"1121B998",
    x"11217A78",
    x"11213B71",
    x"1120FC82",
    x"1120BDAB",
    x"11207EEE",
    x"11204048",
    x"112001BB",
    x"111FC347",
    x"111F84EB",
    x"111F46A7",
    x"111F087C",
    x"111ECA68",
    x"111E8C6E",
    x"111E4E8B",
    x"111E10C0",
    x"111DD30E",
    x"111D9573",
    x"111D57F1",
    x"111D1A87",
    x"111CDD34",
    x"111C9FFA",
    x"111C62D7",
    x"111C25CC",
    x"111BE8DA",
    x"111BABFF",
    x"111B6F3B",
    x"111B3290",
    x"111AF5FC",
    x"111AB97F",
    x"111A7D1B",
    x"111A40CE",
    x"111A0498",
    x"1119C87A",
    x"11198C73",
    x"11195084",
    x"111914AD",
    x"1118D8EC",
    x"11189D43",
    x"111861B1",
    x"11182637",
    x"1117EAD3",
    x"1117AF87",
    x"11177452",
    x"11173934",
    x"1116FE2E",
    x"1116C33E",
    x"11168865",
    x"11164DA3",
    x"111612F8",
    x"1115D864",
    x"11159DE7",
    x"11156381",
    x"11152932",
    x"1114EEF9",
    x"1114B4D7",
    x"11147ACC",
    x"111440D7",
    x"111406F9",
    x"1113CD31",
    x"11139381",
    x"111359E6",
    x"11132062",
    x"1112E6F5",
    x"1112AD9E",
    x"1112745D",
    x"11123B33",
    x"1112021F",
    x"1111C921",
    x"1111903A",
    x"11115769",
    x"11111EAE",
    x"1110E609",
    x"1110AD7A",
    x"11107501",
    x"11103C9E",
    x"11100452",
    x"110FCC1B",
    x"110F93FA",
    x"110F5BEF",
    x"110F23FA",
    x"110EEC1B",
    x"110EB452",
    x"110E7C9E",
    x"110E4501",
    x"110E0D78",
    x"110DD606",
    x"110D9EA9",
    x"110D6762",
    x"110D3030",
    x"110CF914",
    x"110CC20E",
    x"110C8B1D",
    x"110C5441",
    x"110C1D7B",
    x"110BE6CA",
    x"110BB02F",
    x"110B79A8",
    x"110B4338",
    x"110B0CDC",
    x"110AD696",
    x"110AA064",
    x"110A6A48",
    x"110A3441",
    x"1109FE4F",
    x"1109C873",
    x"110992AB",
    x"11095CF8",
    x"1109275A",
    x"1108F1D1",
    x"1108BC5D",
    x"110886FE",
    x"110851B4",
    x"11081C7E",
    x"1107E75D",
    x"1107B251",
    x"11077D5A",
    x"11074877",
    x"110713AA",
    x"1106DEF0",
    x"1106AA4B",
    x"110675BB",
    x"1106413F",
    x"11060CD8",
    x"1105D885",
    x"1105A447",
    x"1105701D",
    x"11053C07",
    x"11050806",
    x"1104D419",
    x"1104A040",
    x"11046C7C",
    x"110438CC",
    x"1104052F",
    x"1103D1A7",
    x"11039E34",
    x"11036AD4",
    x"11033788",
    x"11030450",
    x"1102D12D",
    x"11029E1D",
    x"11026B21",
    x"11023839",
    x"11020565",
    x"1101D2A5",
    x"11019FF9",
    x"11016D60",
    x"11013ADB",
    x"1101086A",
    x"1100D60D",
    x"1100A3C3",
    x"1100718D",
    x"11003F6A",
    x"11000D5B",
    x"10FFB6C0",
    x"10FF52F0",
    x"10FEEF47",
    x"10FE8BC5",
    x"10FE2869",
    x"10FDC535",
    x"10FD6227",
    x"10FCFF40",
    x"10FC9C80",
    x"10FC39E6",
    x"10FBD773",
    x"10FB7526",
    x"10FB12FF",
    x"10FAB0FF",
    x"10FA4F25",
    x"10F9ED71",
    x"10F98BE3",
    x"10F92A7C",
    x"10F8C93A",
    x"10F8681F",
    x"10F80729",
    x"10F7A659",
    x"10F745AF",
    x"10F6E52A",
    x"10F684CC",
    x"10F62493",
    x"10F5C47F",
    x"10F56491",
    x"10F504C9",
    x"10F4A525",
    x"10F445A8",
    x"10F3E64F",
    x"10F3871C",
    x"10F3280D",
    x"10F2C924",
    x"10F26A60",
    x"10F20BC1",
    x"10F1AD47",
    x"10F14EF2",
    x"10F0F0C1",
    x"10F092B6",
    x"10F034CF",
    x"10EFD70C",
    x"10EF796F",
    x"10EF1BF5",
    x"10EEBEA1",
    x"10EE6171",
    x"10EE0465",
    x"10EDA77D",
    x"10ED4ABA",
    x"10ECEE1B",
    x"10EC91A0",
    x"10EC3549",
    x"10EBD916",
    x"10EB7D07",
    x"10EB211C",
    x"10EAC555",
    x"10EA69B2",
    x"10EA0E33",
    x"10E9B2D7",
    x"10E9579F",
    x"10E8FC8B",
    x"10E8A19A",
    x"10E846CC",
    x"10E7EC22",
    x"10E7919C",
    x"10E73739",
    x"10E6DCF9",
    x"10E682DC",
    x"10E628E2",
    x"10E5CF0C",
    x"10E57559",
    x"10E51BC8",
    x"10E4C25B",
    x"10E46910",
    x"10E40FE9",
    x"10E3B6E4",
    x"10E35E02",
    x"10E30543",
    x"10E2ACA6",
    x"10E2542C",
    x"10E1FBD4",
    x"10E1A39F",
    x"10E14B8C",
    x"10E0F39C",
    x"10E09BCE",
    x"10E04422",
    x"10DFEC99",
    x"10DF9531",
    x"10DF3DEC",
    x"10DEE6C9",
    x"10DE8FC8",
    x"10DE38E9",
    x"10DDE22B",
    x"10DD8B90",
    x"10DD3516",
    x"10DCDEBE",
    x"10DC8888",
    x"10DC3274",
    x"10DBDC81",
    x"10DB86AF",
    x"10DB3100",
    x"10DADB71",
    x"10DA8604",
    x"10DA30B8",
    x"10D9DB8E",
    x"10D98685",
    x"10D9319D",
    x"10D8DCD6",
    x"10D88830",
    x"10D833AC",
    x"10D7DF48",
    x"10D78B05",
    x"10D736E3",
    x"10D6E2E2",
    x"10D68F02",
    x"10D63B43",
    x"10D5E7A4",
    x"10D59426",
    x"10D540C8",
    x"10D4ED8B",
    x"10D49A6E",
    x"10D44772",
    x"10D3F497",
    x"10D3A1DB",
    x"10D34F40",
    x"10D2FCC5",
    x"10D2AA6B",
    x"10D25830",
    x"10D20616",
    x"10D1B41B",
    x"10D16241",
    x"10D11087",
    x"10D0BEEC",
    x"10D06D71",
    x"10D01C16",
    x"10CFCADB",
    x"10CF79C0",
    x"10CF28C4",
    x"10CED7E8",
    x"10CE872C",
    x"10CE368F",
    x"10CDE611",
    x"10CD95B3",
    x"10CD4574",
    x"10CCF554",
    x"10CCA554",
    x"10CC5573",
    x"10CC05B2",
    x"10CBB60F",
    x"10CB668B",
    x"10CB1727",
    x"10CAC7E1",
    x"10CA78BB",
    x"10CA29B3",
    x"10C9DACA",
    x"10C98C00",
    x"10C93D55",
    x"10C8EEC8",
    x"10C8A05A",
    x"10C8520B",
    x"10C803DA",
    x"10C7B5C8",
    x"10C767D4",
    x"10C719FE",
    x"10C6CC48",
    x"10C67EAF",
    x"10C63135",
    x"10C5E3D8",
    x"10C5969B",
    x"10C5497B",
    x"10C4FC79",
    x"10C4AF95",
    x"10C462D0",
    x"10C41628",
    x"10C3C99F",
    x"10C37D33",
    x"10C330E5",
    x"10C2E4B5",
    x"10C298A2",
    x"10C24CAD",
    x"10C200D6",
    x"10C1B51D",
    x"10C16981",
    x"10C11E02",
    x"10C0D2A1",
    x"10C0875E",
    x"10C03C37",
    x"10BFF12F",
    x"10BFA643",
    x"10BF5B75",
    x"10BF10C4",
    x"10BEC630",
    x"10BE7BB9",
    x"10BE315F",
    x"10BDE722",
    x"10BD9D02",
    x"10BD52FF",
    x"10BD0919",
    x"10BCBF50",
    x"10BC75A4",
    x"10BC2C14",
    x"10BBE2A1",
    x"10BB994B",
    x"10BB5012",
    x"10BB06F5",
    x"10BABDF4",
    x"10BA7510",
    x"10BA2C49",
    x"10B9E39E",
    x"10B99B0F",
    x"10B9529D",
    x"10B90A46",
    x"10B8C20C",
    x"10B879EF",
    x"10B831ED",
    x"10B7EA08",
    x"10B7A23E",
    x"10B75A91",
    x"10B71300",
    x"10B6CB8A",
    x"10B68431",
    x"10B63CF3",
    x"10B5F5D1",
    x"10B5AECB",
    x"10B567E0",
    x"10B52112",
    x"10B4DA5F",
    x"10B493C7",
    x"10B44D4B",
    x"10B406EB",
    x"10B3C0A6",
    x"10B37A7C",
    x"10B3346E",
    x"10B2EE7B",
    x"10B2A8A4",
    x"10B262E7",
    x"10B21D46",
    x"10B1D7C0",
    x"10B19256",
    x"10B14D06",
    x"10B107D2",
    x"10B0C2B8",
    x"10B07DB9",
    x"10B038D6",
    x"10AFF40D",
    x"10AFAF5F",
    x"10AF6ACC",
    x"10AF2654",
    x"10AEE1F6",
    x"10AE9DB3",
    x"10AE598B",
    x"10AE157D",
    x"10ADD18A",
    x"10AD8DB1",
    x"10AD49F3",
    x"10AD0650",
    x"10ACC2C6",
    x"10AC7F57",
    x"10AC3C03",
    x"10ABF8C9",
    x"10ABB5A8",
    x"10AB72A3",
    x"10AB2FB7",
    x"10AAECE5",
    x"10AAAA2E",
    x"10AA6790",
    x"10AA250D",
    x"10A9E2A3",
    x"10A9A054",
    x"10A95E1E",
    x"10A91C02",
    x"10A8DA00",
    x"10A89818",
    x"10A85649",
    x"10A81495",
    x"10A7D2F9",
    x"10A79178",
    x"10A75010",
    x"10A70EC1",
    x"10A6CD8C",
    x"10A68C71",
    x"10A64B6E",
    x"10A60A86",
    x"10A5C9B6",
    x"10A58900",
    x"10A54863",
    x"10A507DF",
    x"10A4C775",
    x"10A48724",
    x"10A446EB",
    x"10A406CC",
    x"10A3C6C6",
    x"10A386D9",
    x"10A34705",
    x"10A30749",
    x"10A2C7A7",
    x"10A2881D",
    x"10A248AD",
    x"10A20955",
    x"10A1CA15",
    x"10A18AEF",
    x"10A14BE1",
    x"10A10CEB",
    x"10A0CE0F",
    x"10A08F4A",
    x"10A0509F",
    x"10A0120B",
    x"109FD391",
    x"109F952E",
    x"109F56E4",
    x"109F18B2",
    x"109EDA99",
    x"109E9C97",
    x"109E5EAE",
    x"109E20DD",
    x"109DE325",
    x"109DA584",
    x"109D67FB",
    x"109D2A8B",
    x"109CED32",
    x"109CAFF1",
    x"109C72C9",
    x"109C35B8",
    x"109BF8BF",
    x"109BBBDD",
    x"109B7F14",
    x"109B4262",
    x"109B05C8",
    x"109AC946",
    x"109A8CDB",
    x"109A5088",
    x"109A144C",
    x"1099D828",
    x"10999C1B",
    x"10996026",
    x"10992448",
    x"1098E881",
    x"1098ACD2",
    x"1098713A",
    x"109835BA",
    x"1097FA50",
    x"1097BEFE",
    x"109783C3",
    x"1097489F",
    x"10970D92",
    x"1096D29D",
    x"109697BE",
    x"10965CF6",
    x"10962245",
    x"1095E7AB",
    x"1095AD28",
    x"109572BC",
    x"10953866",
    x"1094FE28",
    x"1094C400",
    x"109489EF",
    x"10944FF4",
    x"10941610",
    x"1093DC43",
    x"1093A28C",
    x"109368EC",
    x"10932F62",
    x"1092F5EF",
    x"1092BC92",
    x"1092834C",
    x"10924A1B",
    x"10921102",
    x"1091D7FE",
    x"10919F11",
    x"1091663A",
    x"10912D79",
    x"1090F4CE",
    x"1090BC3A",
    x"109083BB",
    x"10904B53",
    x"10901300",
    x"108FDAC4",
    x"108FA29D",
    x"108F6A8D",
    x"108F3292",
    x"108EFAAD",
    x"108EC2DE",
    x"108E8B25",
    x"108E5382",
    x"108E1BF4",
    x"108DE47C",
    x"108DAD19",
    x"108D75CD",
    x"108D3E95",
    x"108D0774",
    x"108CD067",
    x"108C9971",
    x"108C6290",
    x"108C2BC4",
    x"108BF50D",
    x"108BBE6C",
    x"108B87E1",
    x"108B516A",
    x"108B1B09",
    x"108AE4BD",
    x"108AAE86",
    x"108A7865",
    x"108A4258",
    x"108A0C61",
    x"1089D67F",
    x"1089A0B1",
    x"10896AF9",
    x"10893556",
    x"1088FFC7",
    x"1088CA4E",
    x"108894E9",
    x"10885F99",
    x"10882A5F",
    x"1087F538",
    x"1087C027",
    x"10878B2A",
    x"10875642",
    x"1087216F",
    x"1086ECB0",
    x"1086B806",
    x"10868370",
    x"10864EEF",
    x"10861A83",
    x"1085E62B",
    x"1085B1E7",
    x"10857DB8",
    x"1085499D",
    x"10851596",
    x"1084E1A4",
    x"1084ADC6",
    x"108479FC",
    x"10844646",
    x"108412A5",
    x"1083DF18",
    x"1083AB9F",
    x"1083783A",
    x"108344E9",
    x"108311AC",
    x"1082DE83",
    x"1082AB6E",
    x"1082786D",
    x"10824580",
    x"108212A7",
    x"1081DFE1",
    x"1081AD30",
    x"10817A92",
    x"10814808",
    x"10811592",
    x"1080E32F",
    x"1080B0E0",
    x"10807EA5",
    x"10804C7D",
    x"10801A69",
    x"107FD0D1",
    x"107F6CF7",
    x"107F0944",
    x"107EA5B8",
    x"107E4253",
    x"107DDF14",
    x"107D7BFC",
    x"107D190B",
    x"107CB641",
    x"107C539D",
    x"107BF11F",
    x"107B8EC9",
    x"107B2C98",
    x"107ACA8E",
    x"107A68AA",
    x"107A06EC",
    x"1079A554",
    x"107943E3",
    x"1078E297",
    x"10788172",
    x"10782072",
    x"1077BF98",
    x"10775EE4",
    x"1076FE56",
    x"10769DEE",
    x"10763DAB",
    x"1075DD8D",
    x"10757D96",
    x"10751DC3",
    x"1074BE16",
    x"10745E8F",
    x"1073FF2C",
    x"10739FEF",
    x"107340D7",
    x"1072E1E5",
    x"10728317",
    x"1072246E",
    x"1071C5EA",
    x"1071678C",
    x"10710952",
    x"1070AB3C",
    x"10704D4C",
    x"106FEF80",
    x"106F91D9",
    x"106F3456",
    x"106ED6F8",
    x"106E79BE",
    x"106E1CA9",
    x"106DBFB8",
    x"106D62EB",
    x"106D0642",
    x"106CA9BE",
    x"106C4D5E",
    x"106BF121",
    x"106B9509",
    x"106B3915",
    x"106ADD45",
    x"106A8198",
    x"106A260F",
    x"1069CAAA",
    x"10696F69",
    x"1069144B",
    x"1068B951",
    x"10685E7B",
    x"106803C7",
    x"1067A938",
    x"10674ECB",
    x"1066F482",
    x"10669A5C",
    x"10664059",
    x"1065E67A",
    x"10658CBD",
    x"10653324",
    x"1064D9AD",
    x"1064805A",
    x"10642729",
    x"1063CE1B",
    x"10637530",
    x"10631C68",
    x"1062C3C2",
    x"10626B3F",
    x"106212DE",
    x"1061BAA0",
    x"10616284",
    x"10610A8B",
    x"1060B2B4",
    x"10605AFF",
    x"1060036D",
    x"105FABFD",
    x"105F54AE",
    x"105EFD82",
    x"105EA678",
    x"105E4F90",
    x"105DF8CA",
    x"105DA226",
    x"105D4BA3",
    x"105CF543",
    x"105C9F04",
    x"105C48E7",
    x"105BF2EB",
    x"105B9D11",
    x"105B4758",
    x"105AF1C1",
    x"105A9C4B",
    x"105A46F7",
    x"1059F1C4",
    x"10599CB2",
    x"105947C1",
    x"1058F2F2",
    x"10589E44",
    x"105849B6",
    x"1057F54A",
    x"1057A0FF",
    x"10574CD4",
    x"1056F8CB",
    x"1056A4E2",
    x"1056511A",
    x"1055FD72",
    x"1055A9EC",
    x"10555686",
    x"10550340",
    x"1054B01B",
    x"10545D16",
    x"10540A32",
    x"1053B76F",
    x"105364CB",
    x"10531248",
    x"1052BFE5",
    x"10526DA2",
    x"10521B7F",
    x"1051C97C",
    x"1051779A",
    x"105125D7",
    x"1050D434",
    x"105082B1",
    x"1050314E",
    x"104FE00B",
    x"104F8EE7",
    x"104F3DE3",
    x"104EECFE",
    x"104E9C3A",
    x"104E4B94",
    x"104DFB0F",
    x"104DAAA8",
    x"104D5A61",
    x"104D0A3A",
    x"104CBA31",
    x"104C6A48",
    x"104C1A7E",
    x"104BCAD3",
    x"104B7B48",
    x"104B2BDB",
    x"104ADC8D",
    x"104A8D5F",
    x"104A3E4F",
    x"1049EF5E",
    x"1049A08C",
    x"104951D9",
    x"10490344",
    x"1048B4CE",
    x"10486677",
    x"1048183E",
    x"1047CA24",
    x"10477C28",
    x"10472E4B",
    x"1046E08C",
    x"104692EB",
    x"10464569",
    x"1045F805",
    x"1045AABF",
    x"10455D98",
    x"1045108E",
    x"1044C3A3",
    x"104476D5",
    x"10442A26",
    x"1043DD94",
    x"10439121",
    x"104344CB",
    x"1042F893",
    x"1042AC79",
    x"1042607C",
    x"1042149D",
    x"1041C8DC",
    x"10417D38",
    x"104131B2",
    x"1040E64A",
    x"10409AFE",
    x"10404FD1",
    x"104004C0",
    x"103FB9CD",
    x"103F6EF7",
    x"103F243E",
    x"103ED9A3",
    x"103E8F24",
    x"103E44C3",
    x"103DFA7E",
    x"103DB057",
    x"103D664D",
    x"103D1C5F",
    x"103CD28E",
    x"103C88DB",
    x"103C3F43",
    x"103BF5C9",
    x"103BAC6B",
    x"103B632A",
    x"103B1A06",
    x"103AD0FE",
    x"103A8813",
    x"103A3F44",
    x"1039F691",
    x"1039ADFB",
    x"10396581",
    x"10391D24",
    x"1038D4E2",
    x"10388CBD",
    x"103844B4",
    x"1037FCC8",
    x"1037B4F7",
    x"10376D42",
    x"103725AA",
    x"1036DE2D",
    x"103696CC",
    x"10364F87",
    x"1036085E",
    x"1035C150",
    x"10357A5F",
    x"10353389",
    x"1034ECCF",
    x"1034A630",
    x"10345FAD",
    x"10341945",
    x"1033D2F9",
    x"10338CC8",
    x"103346B3",
    x"103300B9",
    x"1032BADA",
    x"10327517",
    x"10322F6F",
    x"1031E9E2",
    x"1031A470",
    x"10315F19",
    x"103119DE",
    x"1030D4BD",
    x"10308FB8",
    x"10304ACD",
    x"103005FD",
    x"102FC148",
    x"102F7CAE",
    x"102F382F",
    x"102EF3CA",
    x"102EAF80",
    x"102E6B51",
    x"102E273D",
    x"102DE342",
    x"102D9F63",
    x"102D5B9E",
    x"102D17F3",
    x"102CD463",
    x"102C90ED",
    x"102C4D92",
    x"102C0A51",
    x"102BC72A",
    x"102B841D",
    x"102B412B",
    x"102AFE52",
    x"102ABB94",
    x"102A78F0",
    x"102A3665",
    x"1029F3F5",
    x"1029B19F",
    x"10296F62",
    x"10292D40",
    x"1028EB37",
    x"1028A948",
    x"10286773",
    x"102825B7",
    x"1027E415",
    x"1027A28D",
    x"1027611E",
    x"10271FC9",
    x"1026DE8D",
    x"10269D6B",
    x"10265C62",
    x"10261B73",
    x"1025DA9D",
    x"102599E0",
    x"1025593D",
    x"102518B3",
    x"1024D841",
    x"102497EA",
    x"102457AB",
    x"10241785",
    x"1023D778",
    x"10239785",
    x"102357AA",
    x"102317E8",
    x"1022D83F",
    x"102298AF",
    x"10225938",
    x"102219DA",
    x"1021DA94",
    x"10219B67",
    x"10215C52",
    x"10211D57",
    x"1020DE73",
    x"10209FA9",
    x"102060F7",
    x"1020225D",
    x"101FE3DC",
    x"101FA573",
    x"101F6723",
    x"101F28EA",
    x"101EEACB",
    x"101EACC3",
    x"101E6ED4",
    x"101E30FC",
    x"101DF33D",
    x"101DB596",
    x"101D7807",
    x"101D3A91",
    x"101CFD32",
    x"101CBFEB",
    x"101C82BC",
    x"101C45A5",
    x"101C08A5",
    x"101BCBBE",
    x"101B8EEE",
    x"101B5236",
    x"101B1596",
    x"101AD90D",
    x"101A9C9C",
    x"101A6043",
    x"101A2401",
    x"1019E7D7",
    x"1019ABC4",
    x"10196FC9",
    x"101933E5",
    x"1018F818",
    x"1018BC63",
    x"101880C5",
    x"1018453E",
    x"101809CF",
    x"1017CE77",
    x"10179335",
    x"1017580B",
    x"10171CF9",
    x"1016E1FD",
    x"1016A718",
    x"10166C4A",
    x"10163193",
    x"1015F6F4",
    x"1015BC6B",
    x"101581F8",
    x"1015479D",
    x"10150D58",
    x"1014D32B",
    x"10149913",
    x"10145F13",
    x"10142529",
    x"1013EB56",
    x"1013B199",
    x"101377F3",
    x"10133E64",
    x"101304EA",
    x"1012CB88",
    x"1012923B",
    x"10125905",
    x"10121FE6",
    x"1011E6DC",
    x"1011ADE9",
    x"1011750D",
    x"10113C46",
    x"10110395",
    x"1010CAFB",
    x"10109277",
    x"10105A09",
    x"101021B1",
    x"100FE96E",
    x"100FB142",
    x"100F792C",
    x"100F412B",
    x"100F0941",
    x"100ED16C",
    x"100E99AD",
    x"100E6204",
    x"100E2A71",
    x"100DF2F3",
    x"100DBB8B",
    x"100D8438",
    x"100D4CFC",
    x"100D15D4",
    x"100CDEC3",
    x"100CA7C6",
    x"100C70DF",
    x"100C3A0E",
    x"100C0352",
    x"100BCCAB",
    x"100B961A",
    x"100B5F9E",
    x"100B2937",
    x"100AF2E6",
    x"100ABCAA",
    x"100A8683",
    x"100A5071",
    x"100A1A74",
    x"1009E48C",
    x"1009AEB9",
    x"100978FB",
    x"10094353",
    x"10090DBF",
    x"1008D840",
    x"1008A2D6",
    x"10086D81",
    x"10083840",
    x"10080315",
    x"1007CDFE",
    x"100798FC",
    x"1007640E",
    x"10072F36",
    x"1006FA71",
    x"1006C5C2",
    x"10069127",
    x"10065CA1",
    x"1006282F",
    x"1005F3D1",
    x"1005BF88",
    x"10058B53",
    x"10055733",
    x"10052327",
    x"1004EF30",
    x"1004BB4C",
    x"1004877D",
    x"100453C3",
    x"1004201C",
    x"1003EC8A",
    x"1003B90B",
    x"100385A1",
    x"1003524B",
    x"10031F09",
    x"1002EBDB",
    x"1002B8C0",
    x"100285BA",
    x"100252C8",
    x"10021FE9",
    x"1001ED1F",
    x"1001BA68",
    x"100187C5",
    x"10015536",
    x"100122BB",
    x"1000F053",
    x"1000BDFF",
    x"10008BBF",
    x"10005992",
    x"10002779",
    x"0FFFEAE6",
    x"0FFF8702",
    x"0FFF2344",
    x"0FFEBFAE",
    x"0FFE5C3F",
    x"0FFDF8F6",
    x"0FFD95D4",
    x"0FFD32D9",
    x"0FFCD004",
    x"0FFC6D56",
    x"0FFC0ACF",
    x"0FFBA86E",
    x"0FFB4633",
    x"0FFAE41F",
    x"0FFA8231",
    x"0FFA2069",
    x"0FF9BEC8",
    x"0FF95D4C",
    x"0FF8FBF7",
    x"0FF89AC7",
    x"0FF839BE",
    x"0FF7D8DA",
    x"0FF7781C",
    x"0FF71784",
    x"0FF6B712",
    x"0FF656C5",
    x"0FF5F69E",
    x"0FF5969D",
    x"0FF536C1",
    x"0FF4D70A",
    x"0FF47778",
    x"0FF4180C",
    x"0FF3B8C6",
    x"0FF359A4",
    x"0FF2FAA8",
    x"0FF29BD0",
    x"0FF23D1E",
    x"0FF1DE90",
    x"0FF18028",
    x"0FF121E4",
    x"0FF0C3C5",
    x"0FF065CB",
    x"0FF007F6",
    x"0FEFAA45",
    x"0FEF4CB9",
    x"0FEEEF51",
    x"0FEE920E",
    x"0FEE34EF",
    x"0FEDD7F5",
    x"0FED7B1E",
    x"0FED1E6C",
    x"0FECC1DF",
    x"0FEC6575",
    x"0FEC092F",
    x"0FEBAD0E",
    x"0FEB5110",
    x"0FEAF536",
    x"0FEA9980",
    x"0FEA3DEE",
    x"0FE9E280",
    x"0FE98735",
    x"0FE92C0E",
    x"0FE8D10B",
    x"0FE8762B",
    x"0FE81B6F",
    x"0FE7C0D6",
    x"0FE76660",
    x"0FE70C0E",
    x"0FE6B1DF",
    x"0FE657D3",
    x"0FE5FDEA",
    x"0FE5A424",
    x"0FE54A82",
    x"0FE4F102",
    x"0FE497A5",
    x"0FE43E6C",
    x"0FE3E555",
    x"0FE38C60",
    x"0FE3338F",
    x"0FE2DAE0",
    x"0FE28254",
    x"0FE229EA",
    x"0FE1D1A3",
    x"0FE1797E",
    x"0FE1217C",
    x"0FE0C99C",
    x"0FE071DF",
    x"0FE01A43",
    x"0FDFC2CA",
    x"0FDF6B73",
    x"0FDF143E",
    x"0FDEBD2B",
    x"0FDE663A",
    x"0FDE0F6B",
    x"0FDDB8BE",
    x"0FDD6233",
    x"0FDD0BCA",
    x"0FDCB582",
    x"0FDC5F5C",
    x"0FDC0957",
    x"0FDBB374",
    x"0FDB5DB3",
    x"0FDB0813",
    x"0FDAB295",
    x"0FDA5D38",
    x"0FDA07FC",
    x"0FD9B2E1",
    x"0FD95DE8",
    x"0FD90910",
    x"0FD8B459",
    x"0FD85FC3",
    x"0FD80B4E",
    x"0FD7B6FA",
    x"0FD762C7",
    x"0FD70EB5",
    x"0FD6BAC4",
    x"0FD666F3",
    x"0FD61343",
    x"0FD5BFB4",
    x"0FD56C45",
    x"0FD518F7",
    x"0FD4C5CA",
    x"0FD472BD",
    x"0FD41FD0",
    x"0FD3CD04",
    x"0FD37A58",
    x"0FD327CC",
    x"0FD2D561",
    x"0FD28316",
    x"0FD230EB",
    x"0FD1DEE0",
    x"0FD18CF4",
    x"0FD13B29",
    x"0FD0E97E",
    x"0FD097F3",
    x"0FD04687",
    x"0FCFF53C",
    x"0FCFA410",
    x"0FCF5304",
    x"0FCF0217",
    x"0FCEB14A",
    x"0FCE609C",
    x"0FCE100E",
    x"0FCDBFA0",
    x"0FCD6F51",
    x"0FCD1F21",
    x"0FCCCF10",
    x"0FCC7F1F",
    x"0FCC2F4D",
    x"0FCBDF9A",
    x"0FCB9006",
    x"0FCB4092",
    x"0FCAF13C",
    x"0FCAA205",
    x"0FCA52ED",
    x"0FCA03F4",
    x"0FC9B51A",
    x"0FC9665F",
    x"0FC917C2",
    x"0FC8C944",
    x"0FC87AE5",
    x"0FC82CA4",
    x"0FC7DE82",
    x"0FC7907E",
    x"0FC74299",
    x"0FC6F4D2",
    x"0FC6A72A",
    x"0FC659A0",
    x"0FC60C34",
    x"0FC5BEE6",
    x"0FC571B7",
    x"0FC524A5",
    x"0FC4D7B2",
    x"0FC48ADD",
    x"0FC43E26",
    x"0FC3F18C",
    x"0FC3A511",
    x"0FC358B3",
    x"0FC30C74",
    x"0FC2C052",
    x"0FC2744D",
    x"0FC22867",
    x"0FC1DC9E",
    x"0FC190F2",
    x"0FC14564",
    x"0FC0F9F4",
    x"0FC0AEA1",
    x"0FC0636C",
    x"0FC01853",
    x"0FBFCD59",
    x"0FBF827B",
    x"0FBF37BB",
    x"0FBEED17",
    x"0FBEA291",
    x"0FBE5828",
    x"0FBE0DDD",
    x"0FBDC3AE",
    x"0FBD799C",
    x"0FBD2FA7",
    x"0FBCE5CE",
    x"0FBC9C13",
    x"0FBC5274",
    x"0FBC08F3",
    x"0FBBBF8D",
    x"0FBB7645",
    x"0FBB2D19",
    x"0FBAE40A",
    x"0FBA9B17",
    x"0FBA5241",
    x"0FBA0987",
    x"0FB9C0E9",
    x"0FB97868",
    x"0FB93003",
    x"0FB8E7BA",
    x"0FB89F8E",
    x"0FB8577E",
    x"0FB80F8A",
    x"0FB7C7B2",
    x"0FB77FF6",
    x"0FB73856",
    x"0FB6F0D2",
    x"0FB6A969",
    x"0FB6621D",
    x"0FB61AED",
    x"0FB5D3D8",
    x"0FB58CDF",
    x"0FB54602",
    x"0FB4FF40",
    x"0FB4B89B",
    x"0FB47210",
    x"0FB42BA1",
    x"0FB3E54E",
    x"0FB39F16",
    x"0FB358FA",
    x"0FB312F9",
    x"0FB2CD13",
    x"0FB28749",
    x"0FB24199",
    x"0FB1FC05",
    x"0FB1B68C",
    x"0FB1712F",
    x"0FB12BEC",
    x"0FB0E6C4",
    x"0FB0A1B8",
    x"0FB05CC6",
    x"0FB017EF",
    x"0FAFD333",
    x"0FAF8E92",
    x"0FAF4A0C",
    x"0FAF05A0",
    x"0FAEC14F",
    x"0FAE7D19",
    x"0FAE38FE",
    x"0FADF4FD",
    x"0FADB116",
    x"0FAD6D4A",
    x"0FAD2999",
    x"0FACE602",
    x"0FACA285",
    x"0FAC5F23",
    x"0FAC1BDB",
    x"0FABD8AD",
    x"0FAB959A",
    x"0FAB52A0",
    x"0FAB0FC1",
    x"0FAACCFC",
    x"0FAA8A51",
    x"0FAA47C0",
    x"0FAA0549",
    x"0FA9C2EC",
    x"0FA980A8",
    x"0FA93E7F",
    x"0FA8FC70",
    x"0FA8BA7A",
    x"0FA8789E",
    x"0FA836DC",
    x"0FA7F533",
    x"0FA7B3A4",
    x"0FA7722F",
    x"0FA730D3",
    x"0FA6EF91",
    x"0FA6AE68",
    x"0FA66D58",
    x"0FA62C62",
    x"0FA5EB86",
    x"0FA5AAC2",
    x"0FA56A18",
    x"0FA52987",
    x"0FA4E910",
    x"0FA4A8B1",
    x"0FA4686C",
    x"0FA42840",
    x"0FA3E82C",
    x"0FA3A832",
    x"0FA36851",
    x"0FA32889",
    x"0FA2E8D9",
    x"0FA2A943",
    x"0FA269C5",
    x"0FA22A60",
    x"0FA1EB14",
    x"0FA1ABE1",
    x"0FA16CC6",
    x"0FA12DC4",
    x"0FA0EEDA",
    x"0FA0B009",
    x"0FA07150",
    x"0FA032B0",
    x"0F9FF429",
    x"0F9FB5BA",
    x"0F9F7763",
    x"0F9F3924",
    x"0F9EFAFE",
    x"0F9EBCF0",
    x"0F9E7EFB",
    x"0F9E411D",
    x"0F9E0358",
    x"0F9DC5AA",
    x"0F9D8815",
    x"0F9D4A98",
    x"0F9D0D33",
    x"0F9CCFE6",
    x"0F9C92B0",
    x"0F9C5593",
    x"0F9C188E",
    x"0F9BDBA0",
    x"0F9B9ECA",
    x"0F9B620C",
    x"0F9B2565",
    x"0F9AE8D7",
    x"0F9AAC60",
    x"0F9A7000",
    x"0F9A33B8",
    x"0F99F788",
    x"0F99BB6F",
    x"0F997F6D",
    x"0F994383",
    x"0F9907B0",
    x"0F98CBF5",
    x"0F989051",
    x"0F9854C4",
    x"0F98194F",
    x"0F97DDF0",
    x"0F97A2A9",
    x"0F976779",
    x"0F972C61",
    x"0F96F15F",
    x"0F96B674",
    x"0F967BA0",
    x"0F9640E3",
    x"0F96063D",
    x"0F95CBAE",
    x"0F959136",
    x"0F9556D5",
    x"0F951C8A",
    x"0F94E257",
    x"0F94A83A",
    x"0F946E33",
    x"0F943444",
    x"0F93FA6A",
    x"0F93C0A8",
    x"0F9386FC",
    x"0F934D66",
    x"0F9313E7",
    x"0F92DA7F",
    x"0F92A12D",
    x"0F9267F1",
    x"0F922ECB",
    x"0F91F5BC",
    x"0F91BCC3",
    x"0F9183E1",
    x"0F914B14",
    x"0F91125E",
    x"0F90D9BE",
    x"0F90A134",
    x"0F9068C0",
    x"0F903062",
    x"0F8FF81A",
    x"0F8FBFE8",
    x"0F8F87CC",
    x"0F8F4FC6",
    x"0F8F17D6",
    x"0F8EDFFC",
    x"0F8EA837",
    x"0F8E7088",
    x"0F8E38EF",
    x"0F8E016C",
    x"0F8DC9FE",
    x"0F8D92A6",
    x"0F8D5B63",
    x"0F8D2436",
    x"0F8CED1F",
    x"0F8CB61D",
    x"0F8C7F31",
    x"0F8C485A",
    x"0F8C1198",
    x"0F8BDAEC",
    x"0F8BA455",
    x"0F8B6DD4",
    x"0F8B3767",
    x"0F8B0110",
    x"0F8ACACF",
    x"0F8A94A2",
    x"0F8A5E8A",
    x"0F8A2888",
    x"0F89F29B",
    x"0F89BCC3",
    x"0F8986FF",
    x"0F895151",
    x"0F891BB8",
    x"0F88E633",
    x"0F88B0C4",
    x"0F887B69",
    x"0F884623",
    x"0F8810F2",
    x"0F87DBD6",
    x"0F87A6CF",
    x"0F8771DC",
    x"0F873CFE",
    x"0F870834",
    x"0F86D37F",
    x"0F869EDF",
    x"0F866A53",
    x"0F8635DC",
    x"0F860179",
    x"0F85CD2B",
    x"0F8598F1",
    x"0F8564CB",
    x"0F8530BA",
    x"0F84FCBD",
    x"0F84C8D5",
    x"0F849500",
    x"0F846140",
    x"0F842D94",
    x"0F83F9FD",
    x"0F83C679",
    x"0F83930A",
    x"0F835FAE",
    x"0F832C67",
    x"0F82F933",
    x"0F82C614",
    x"0F829309",
    x"0F826011",
    x"0F822D2E",
    x"0F81FA5E",
    x"0F81C7A2",
    x"0F8194FA",
    x"0F816266",
    x"0F812FE5",
    x"0F80FD78",
    x"0F80CB1F",
    x"0F8098D9",
    x"0F8066A8",
    x"0F803489",
    x"0F80027E",
    x"0F7FA10F",
    x"0F7F3D47",
    x"0F7ED9A7",
    x"0F7E762D",
    x"0F7E12DA",
    x"0F7DAFAE",
    x"0F7D4CA9",
    x"0F7CE9CA",
    x"0F7C8712",
    x"0F7C2481",
    x"0F7BC216",
    x"0F7B5FD1",
    x"0F7AFDB3",
    x"0F7A9BBB",
    x"0F7A39E9",
    x"0F79D83E",
    x"0F7976B8",
    x"0F791559",
    x"0F78B420",
    x"0F78530C",
    x"0F77F21F",
    x"0F779157",
    x"0F7730B5",
    x"0F76D039",
    x"0F766FE2",
    x"0F760FB2",
    x"0F75AFA6",
    x"0F754FC0",
    x"0F74F000",
    x"0F749065",
    x"0F7430EF",
    x"0F73D19F",
    x"0F737273",
    x"0F73136D",
    x"0F72B48C",
    x"0F7255D0",
    x"0F71F739",
    x"0F7198C7",
    x"0F713A7A",
    x"0F70DC51",
    x"0F707E4D",
    x"0F70206E",
    x"0F6FC2B4",
    x"0F6F651E",
    x"0F6F07AD",
    x"0F6EAA60",
    x"0F6E4D38",
    x"0F6DF034",
    x"0F6D9354",
    x"0F6D3699",
    x"0F6CDA02",
    x"0F6C7D8F",
    x"0F6C2140",
    x"0F6BC515",
    x"0F6B690E",
    x"0F6B0D2A",
    x"0F6AB16B",
    x"0F6A55D0",
    x"0F69FA58",
    x"0F699F04",
    x"0F6943D4",
    x"0F68E8C7",
    x"0F688DDE",
    x"0F683318",
    x"0F67D876",
    x"0F677DF7",
    x"0F67239C",
    x"0F66C963",
    x"0F666F4E",
    x"0F66155C",
    x"0F65BB8E",
    x"0F6561E2",
    x"0F650859",
    x"0F64AEF3",
    x"0F6455B0",
    x"0F63FC90",
    x"0F63A393",
    x"0F634AB9",
    x"0F62F201",
    x"0F62996B",
    x"0F6240F9",
    x"0F61E8A9",
    x"0F61907B",
    x"0F613870",
    x"0F60E087",
    x"0F6088C0",
    x"0F60311C",
    x"0F5FD99A",
    x"0F5F823A",
    x"0F5F2AFC",
    x"0F5ED3E0",
    x"0F5E7CE7",
    x"0F5E260F",
    x"0F5DCF59",
    x"0F5D78C5",
    x"0F5D2253",
    x"0F5CCC02",
    x"0F5C75D3",
    x"0F5C1FC6",
    x"0F5BC9DA",
    x"0F5B7410",
    x"0F5B1E68",
    x"0F5AC8E0",
    x"0F5A737B",
    x"0F5A1E36",
    x"0F59C913",
    x"0F597411",
    x"0F591F30",
    x"0F58CA71",
    x"0F5875D2",
    x"0F582155",
    x"0F57CCF8",
    x"0F5778BD",
    x"0F5724A2",
    x"0F56D0A8",
    x"0F567CCF",
    x"0F562916",
    x"0F55D57F",
    x"0F558208",
    x"0F552EB1",
    x"0F54DB7B",
    x"0F548866",
    x"0F543571",
    x"0F53E29C",
    x"0F538FE7",
    x"0F533D53",
    x"0F52EAE0",
    x"0F52988C",
    x"0F524658",
    x"0F51F445",
    x"0F51A251",
    x"0F51507E",
    x"0F50FECB",
    x"0F50AD37",
    x"0F505BC3",
    x"0F500A6F",
    x"0F4FB93B",
    x"0F4F6827",
    x"0F4F1732",
    x"0F4EC65C",
    x"0F4E75A7",
    x"0F4E2510",
    x"0F4DD49A",
    x"0F4D8442",
    x"0F4D340A",
    x"0F4CE3F2",
    x"0F4C93F8",
    x"0F4C441E",
    x"0F4BF463",
    x"0F4BA4C7",
    x"0F4B554A",
    x"0F4B05EC",
    x"0F4AB6AE",
    x"0F4A678E",
    x"0F4A188D",
    x"0F49C9AB",
    x"0F497AE7",
    x"0F492C43",
    x"0F48DDBD",
    x"0F488F55",
    x"0F48410D",
    x"0F47F2E2",
    x"0F47A4D7",
    x"0F4756EA",
    x"0F47091B",
    x"0F46BB6B",
    x"0F466DD8",
    x"0F462065",
    x"0F45D30F",
    x"0F4585D8",
    x"0F4538BF",
    x"0F44EBC3",
    x"0F449EE6",
    x"0F445227",
    x"0F440586",
    x"0F43B903",
    x"0F436C9E",
    x"0F432056",
    x"0F42D42C",
    x"0F428820",
    x"0F423C32",
    x"0F41F061",
    x"0F41A4AE",
    x"0F415919",
    x"0F410DA1",
    x"0F40C246",
    x"0F407709",
    x"0F402BE9",
    x"0F3FE0E6",
    x"0F3F9601",
    x"0F3F4B39",
    x"0F3F008E",
    x"0F3EB601",
    x"0F3E6B90",
    x"0F3E213D",
    x"0F3DD706",
    x"0F3D8CED",
    x"0F3D42F0",
    x"0F3CF910",
    x"0F3CAF4E",
    x"0F3C65A7",
    x"0F3C1C1E",
    x"0F3BD2B1",
    x"0F3B8961",
    x"0F3B402E",
    x"0F3AF717",
    x"0F3AAE1D",
    x"0F3A653F",
    x"0F3A1C7E",
    x"0F39D3D9",
    x"0F398B50",
    x"0F3942E4",
    x"0F38FA94",
    x"0F38B260",
    x"0F386A49",
    x"0F38224D",
    x"0F37DA6E",
    x"0F3792AB",
    x"0F374B03",
    x"0F370378",
    x"0F36BC09",
    x"0F3674B5",
    x"0F362D7D",
    x"0F35E662",
    x"0F359F61",
    x"0F35587D",
    x"0F3511B4",
    x"0F34CB07",
    x"0F348476",
    x"0F343E00",
    x"0F33F7A5",
    x"0F33B166",
    x"0F336B43",
    x"0F33253A",
    x"0F32DF4E",
    x"0F32997C",
    x"0F3253C6",
    x"0F320E2A",
    x"0F31C8AB",
    x"0F318346",
    x"0F313DFC",
    x"0F30F8CD",
    x"0F30B3BA",
    x"0F306EC1",
    x"0F3029E3",
    x"0F2FE520",
    x"0F2FA078",
    x"0F2F5BEB",
    x"0F2F1778",
    x"0F2ED320",
    x"0F2E8EE3",
    x"0F2E4AC1",
    x"0F2E06B9",
    x"0F2DC2CB",
    x"0F2D7EF9",
    x"0F2D3B40",
    x"0F2CF7A2",
    x"0F2CB41F",
    x"0F2C70B6",
    x"0F2C2D67",
    x"0F2BEA32",
    x"0F2BA718",
    x"0F2B6418",
    x"0F2B2132",
    x"0F2ADE66",
    x"0F2A9BB4",
    x"0F2A591C",
    x"0F2A169E",
    x"0F29D43A",
    x"0F2991F0",
    x"0F294FC0",
    x"0F290DAA",
    x"0F28CBAE",
    x"0F2889CB",
    x"0F284802",
    x"0F280653",
    x"0F27C4BD",
    x"0F278341",
    x"0F2741DE",
    x"0F270095",
    x"0F26BF66",
    x"0F267E50",
    x"0F263D53",
    x"0F25FC70",
    x"0F25BBA6",
    x"0F257AF5",
    x"0F253A5E",
    x"0F24F9E0",
    x"0F24B97B",
    x"0F24792F",
    x"0F2438FC",
    x"0F23F8E2",
    x"0F23B8E2",
    x"0F2378FA",
    x"0F23392B",
    x"0F22F975",
    x"0F22B9D8",
    x"0F227A54",
    x"0F223AE9",
    x"0F21FB96",
    x"0F21BC5C",
    x"0F217D3B",
    x"0F213E32",
    x"0F20FF42",
    x"0F20C06B",
    x"0F2081AC",
    x"0F204305",
    x"0F200477",
    x"0F1FC602",
    x"0F1F87A5",
    x"0F1F4960",
    x"0F1F0B33",
    x"0F1ECD1F",
    x"0F1E8F23",
    x"0F1E513F",
    x"0F1E1374",
    x"0F1DD5C0",
    x"0F1D9825",
    x"0F1D5AA1",
    x"0F1D1D36",
    x"0F1CDFE2",
    x"0F1CA2A7",
    x"0F1C6583",
    x"0F1C2878",
    x"0F1BEB84",
    x"0F1BAEA8",
    x"0F1B71E3",
    x"0F1B3537",
    x"0F1AF8A2",
    x"0F1ABC24",
    x"0F1A7FBF",
    x"0F1A4370",
    x"0F1A073A",
    x"0F19CB1B",
    x"0F198F13",
    x"0F195323",
    x"0F19174A",
    x"0F18DB89",
    x"0F189FDF",
    x"0F18644C",
    x"0F1828D0",
    x"0F17ED6C",
    x"0F17B21F",
    x"0F1776E9",
    x"0F173BCA",
    x"0F1700C2",
    x"0F16C5D1",
    x"0F168AF8",
    x"0F165035",
    x"0F161589",
    x"0F15DAF4",
    x"0F15A076",
    x"0F15660F",
    x"0F152BBE",
    x"0F14F184",
    x"0F14B761",
    x"0F147D55",
    x"0F14435F",
    x"0F140980",
    x"0F13CFB8",
    x"0F139606",
    x"0F135C6B",
    x"0F1322E6",
    x"0F12E978",
    x"0F12B020",
    x"0F1276DE",
    x"0F123DB3",
    x"0F12049E",
    x"0F11CB9F",
    x"0F1192B7",
    x"0F1159E4",
    x"0F112128",
    x"0F10E883",
    x"0F10AFF3",
    x"0F107779",
    x"0F103F15",
    x"0F1006C8",
    x"0F0FCE90",
    x"0F0F966E",
    x"0F0F5E63",
    x"0F0F266D",
    x"0F0EEE8D",
    x"0F0EB6C2",
    x"0F0E7F0E",
    x"0F0E476F",
    x"0F0E0FE6",
    x"0F0DD873",
    x"0F0DA115",
    x"0F0D69CD",
    x"0F0D329A",
    x"0F0CFB7D",
    x"0F0CC476",
    x"0F0C8D84",
    x"0F0C56A7",
    x"0F0C1FE0",
    x"0F0BE92E",
    x"0F0BB292",
    x"0F0B7C0B",
    x"0F0B4599",
    x"0F0B0F3C",
    x"0F0AD8F5",
    x"0F0AA2C3",
    x"0F0A6CA6",
    x"0F0A369E",
    x"0F0A00AB",
    x"0F09CACD",
    x"0F099505",
    x"0F095F51",
    x"0F0929B2",
    x"0F08F428",
    x"0F08BEB3",
    x"0F088953",
    x"0F085408",
    x"0F081ED2",
    x"0F07E9B0",
    x"0F07B4A3",
    x"0F077FAB",
    x"0F074AC7",
    x"0F0715F8",
    x"0F06E13E",
    x"0F06AC98",
    x"0F067807",
    x"0F06438B",
    x"0F060F23",
    x"0F05DACF",
    x"0F05A690",
    x"0F057265",
    x"0F053E4E",
    x"0F050A4C",
    x"0F04D65E",
    x"0F04A285",
    x"0F046EBF",
    x"0F043B0E",
    x"0F040771",
    x"0F03D3E8",
    x"0F03A073",
    x"0F036D13",
    x"0F0339C6",
    x"0F03068E",
    x"0F02D369",
    x"0F02A058",
    x"0F026D5C",
    x"0F023A73",
    x"0F02079E",
    x"0F01D4DD",
    x"0F01A230",
    x"0F016F96",
    x"0F013D11",
    x"0F010A9F",
    x"0F00D840",
    x"0F00A5F6",
    x"0F0073BF",
    x"0F00419B",
    x"0F000F8B",
    x"0EFFBB1E",
    x"0EFF574D",
    x"0EFEF3A2",
    x"0EFE901E",
    x"0EFE2CC1",
    x"0EFDC98B",
    x"0EFD667C",
    x"0EFD0393",
    x"0EFCA0D1",
    x"0EFC3E35",
    x"0EFBDBC0",
    x"0EFB7972",
    x"0EFB174A",
    x"0EFAB548",
    x"0EFA536C",
    x"0EF9F1B6",
    x"0EF99027",
    x"0EF92EBE",
    x"0EF8CD7A",
    x"0EF86C5D",
    x"0EF80B66",
    x"0EF7AA94",
    x"0EF749E9",
    x"0EF6E963",
    x"0EF68902",
    x"0EF628C7",
    x"0EF5C8B2",
    x"0EF568C3",
    x"0EF508F8",
    x"0EF4A954",
    x"0EF449D4",
    x"0EF3EA7A",
    x"0EF38B45",
    x"0EF32C35",
    x"0EF2CD4A",
    x"0EF26E85",
    x"0EF20FE4",
    x"0EF1B168",
    x"0EF15311",
    x"0EF0F4DF",
    x"0EF096D2",
    x"0EF038EA",
    x"0EEFDB26",
    x"0EEF7D86",
    x"0EEF200C",
    x"0EEEC2B5",
    x"0EEE6583",
    x"0EEE0876",
    x"0EEDAB8D",
    x"0EED4EC8",
    x"0EECF227",
    x"0EEC95AB",
    x"0EEC3952",
    x"0EEBDD1E",
    x"0EEB810D",
    x"0EEB2521",
    x"0EEAC958",
    x"0EEA6DB4",
    x"0EEA1233",
    x"0EE9B6D5",
    x"0EE95B9C",
    x"0EE90086",
    x"0EE8A593",
    x"0EE84AC4",
    x"0EE7F019",
    x"0EE79591",
    x"0EE73B2C",
    x"0EE6E0EB",
    x"0EE686CC",
    x"0EE62CD1",
    x"0EE5D2F9",
    x"0EE57944",
    x"0EE51FB3",
    x"0EE4C644",
    x"0EE46CF8",
    x"0EE413CF",
    x"0EE3BAC8",
    x"0EE361E5",
    x"0EE30924",
    x"0EE2B085",
    x"0EE2580A",
    x"0EE1FFB1",
    x"0EE1A77A",
    x"0EE14F66",
    x"0EE0F774",
    x"0EE09FA4",
    x"0EE047F7",
    x"0EDFF06C",
    x"0EDF9903",
    x"0EDF41BD",
    x"0EDEEA98",
    x"0EDE9395",
    x"0EDE3CB5",
    x"0EDDE5F6",
    x"0EDD8F59",
    x"0EDD38DE",
    x"0EDCE285",
    x"0EDC8C4D",
    x"0EDC3637",
    x"0EDBE043",
    x"0EDB8A70",
    x"0EDB34BE",
    x"0EDADF2F",
    x"0EDA89C0",
    x"0EDA3473",
    x"0ED9DF47",
    x"0ED98A3C",
    x"0ED93553",
    x"0ED8E08B",
    x"0ED88BE4",
    x"0ED8375D",
    x"0ED7E2F8",
    x"0ED78EB4",
    x"0ED73A91",
    x"0ED6E68E",
    x"0ED692AD",
    x"0ED63EEC",
    x"0ED5EB4B",
    x"0ED597CC",
    x"0ED5446D",
    x"0ED4F12E",
    x"0ED49E10",
    x"0ED44B13",
    x"0ED3F836",
    x"0ED3A579",
    x"0ED352DC",
    x"0ED30060",
    x"0ED2AE04",
    x"0ED25BC8",
    x"0ED209AC",
    x"0ED1B7B1",
    x"0ED165D5",
    x"0ED11419",
    x"0ED0C27D",
    x"0ED07101",
    x"0ED01FA5",
    x"0ECFCE68",
    x"0ECF7D4C",
    x"0ECF2C4F",
    x"0ECEDB71",
    x"0ECE8AB3",
    x"0ECE3A15",
    x"0ECDE996",
    x"0ECD9936",
    x"0ECD48F6",
    x"0ECCF8D5",
    x"0ECCA8D4",
    x"0ECC58F1",
    x"0ECC092E",
    x"0ECBB98A",
    x"0ECB6A05",
    x"0ECB1A9F",
    x"0ECACB58",
    x"0ECA7C30",
    x"0ECA2D27",
    x"0EC9DE3D",
    x"0EC98F72",
    x"0EC940C5",
    x"0EC8F237",
    x"0EC8A3C8",
    x"0EC85577",
    x"0EC80745",
    x"0EC7B931",
    x"0EC76B3C",
    x"0EC71D65",
    x"0EC6CFAD",
    x"0EC68213",
    x"0EC63498",
    x"0EC5E73A",
    x"0EC599FB",
    x"0EC54CDA",
    x"0EC4FFD7",
    x"0EC4B2F2",
    x"0EC4662B",
    x"0EC41982",
    x"0EC3CCF7",
    x"0EC3808A",
    x"0EC3343B",
    x"0EC2E809",
    x"0EC29BF5",
    x"0EC24FFF",
    x"0EC20427",
    x"0EC1B86C",
    x"0EC16CCF",
    x"0EC1214F",
    x"0EC0D5ED",
    x"0EC08AA8",
    x"0EC03F80",
    x"0EBFF476",
    x"0EBFA989",
    x"0EBF5EBA",
    x"0EBF1407",
    x"0EBEC972",
    x"0EBE7EFA",
    x"0EBE349F",
    x"0EBDEA61",
    x"0EBDA040",
    x"0EBD563C",
    x"0EBD0C54",
    x"0EBCC28A",
    x"0EBC78DC",
    x"0EBC2F4C",
    x"0EBBE5D7",
    x"0EBB9C80",
    x"0EBB5345",
    x"0EBB0A27",
    x"0EBAC125",
    x"0EBA7840",
    x"0EBA2F77",
    x"0EB9E6CB",
    x"0EB99E3B",
    x"0EB955C7",
    x"0EB90D70",
    x"0EB8C535",
    x"0EB87D16",
    x"0EB83513",
    x"0EB7ED2C",
    x"0EB7A562",
    x"0EB75DB3",
    x"0EB71620",
    x"0EB6CEAA",
    x"0EB6874F",
    x"0EB64010",
    x"0EB5F8ED",
    x"0EB5B1E6",
    x"0EB56AFA",
    x"0EB5242A",
    x"0EB4DD76",
    x"0EB496DD",
    x"0EB45060",
    x"0EB409FE",
    x"0EB3C3B8",
    x"0EB37D8D",
    x"0EB3377E",
    x"0EB2F18A",
    x"0EB2ABB1",
    x"0EB265F4",
    x"0EB22052",
    x"0EB1DACA",
    x"0EB1955F",
    x"0EB1500E",
    x"0EB10AD8",
    x"0EB0C5BD",
    x"0EB080BE",
    x"0EB03BD9",
    x"0EAFF70F",
    x"0EAFB260",
    x"0EAF6DCB",
    x"0EAF2952",
    x"0EAEE4F3",
    x"0EAEA0AF",
    x"0EAE5C86",
    x"0EAE1877",
    x"0EADD482",
    x"0EAD90A9",
    x"0EAD4CE9",
    x"0EAD0945",
    x"0EACC5BA",
    x"0EAC824A",
    x"0EAC3EF4",
    x"0EABFBB9",
    x"0EABB898",
    x"0EAB7591",
    x"0EAB32A4",
    x"0EAAEFD1",
    x"0EAAAD18",
    x"0EAA6A7A",
    x"0EAA27F5",
    x"0EA9E58B",
    x"0EA9A33A",
    x"0EA96103",
    x"0EA91EE6",
    x"0EA8DCE3",
    x"0EA89AF9",
    x"0EA8592A",
    x"0EA81774",
    x"0EA7D5D7",
    x"0EA79455",
    x"0EA752EC",
    x"0EA7119C",
    x"0EA6D066",
    x"0EA68F49",
    x"0EA64E46",
    x"0EA60D5C",
    x"0EA5CC8B",
    x"0EA58BD4",
    x"0EA54B36",
    x"0EA50AB1",
    x"0EA4CA46",
    x"0EA489F3",
    x"0EA449BA",
    x"0EA4099A",
    x"0EA3C992",
    x"0EA389A4",
    x"0EA349CF",
    x"0EA30A13",
    x"0EA2CA6F",
    x"0EA28AE4",
    x"0EA24B73",
    x"0EA20C19",
    x"0EA1CCD9",
    x"0EA18DB1",
    x"0EA14EA2",
    x"0EA10FAC",
    x"0EA0D0CE",
    x"0EA09209",
    x"0EA0535C",
    x"0EA014C8",
    x"0E9FD64C",
    x"0E9F97E8",
    x"0E9F599D",
    x"0E9F1B6A",
    x"0E9EDD50",
    x"0E9E9F4D",
    x"0E9E6163",
    x"0E9E2391",
    x"0E9DE5D7",
    x"0E9DA836",
    x"0E9D6AAC",
    x"0E9D2D3A",
    x"0E9CEFE1",
    x"0E9CB29F",
    x"0E9C7575",
    x"0E9C3863",
    x"0E9BFB69",
    x"0E9BBE87",
    x"0E9B81BC",
    x"0E9B4509",
    x"0E9B086E",
    x"0E9ACBEB",
    x"0E9A8F7F",
    x"0E9A532B",
    x"0E9A16EE",
    x"0E99DAC9",
    x"0E999EBB",
    x"0E9962C5",
    x"0E9926E6",
    x"0E98EB1E",
    x"0E98AF6E",
    x"0E9873D5",
    x"0E983854",
    x"0E97FCE9",
    x"0E97C196",
    x"0E97865A",
    x"0E974B35",
    x"0E971027",
    x"0E96D530",
    x"0E969A51",
    x"0E965F88",
    x"0E9624D6",
    x"0E95EA3B",
    x"0E95AFB7",
    x"0E95754A",
    x"0E953AF3",
    x"0E9500B4",
    x"0E94C68B",
    x"0E948C79",
    x"0E94527D",
    x"0E941898",
    x"0E93DECA",
    x"0E93A512",
    x"0E936B71",
    x"0E9331E6",
    x"0E92F872",
    x"0E92BF14",
    x"0E9285CC",
    x"0E924C9B",
    x"0E921381",
    x"0E91DA7C",
    x"0E91A18E",
    x"0E9168B6",
    x"0E912FF4",
    x"0E90F748",
    x"0E90BEB3",
    x"0E908633",
    x"0E904DCA",
    x"0E901577",
    x"0E8FDD39",
    x"0E8FA512",
    x"0E8F6D00",
    x"0E8F3505",
    x"0E8EFD1F",
    x"0E8EC54F",
    x"0E8E8D95",
    x"0E8E55F0",
    x"0E8E1E62",
    x"0E8DE6E9",
    x"0E8DAF85",
    x"0E8D7837",
    x"0E8D40FF",
    x"0E8D09DD",
    x"0E8CD2CF",
    x"0E8C9BD8",
    x"0E8C64F6",
    x"0E8C2E29",
    x"0E8BF772",
    x"0E8BC0D0",
    x"0E8B8A43",
    x"0E8B53CC",
    x"0E8B1D6A",
    x"0E8AE71D",
    x"0E8AB0E5",
    x"0E8A7AC2",
    x"0E8A44B5",
    x"0E8A0EBD",
    x"0E89D8DA",
    x"0E89A30B",
    x"0E896D52",
    x"0E8937AE",
    x"0E89021F",
    x"0E88CCA4",
    x"0E88973F",
    x"0E8861EE",
    x"0E882CB2",
    x"0E87F78B",
    x"0E87C279",
    x"0E878D7B",
    x"0E875892",
    x"0E8723BE",
    x"0E86EEFE",
    x"0E86BA53",
    x"0E8685BD",
    x"0E86513B",
    x"0E861CCD",
    x"0E85E874",
    x"0E85B430",
    x"0E857FFF",
    x"0E854BE4",
    x"0E8517DC",
    x"0E84E3E9",
    x"0E84B00A",
    x"0E847C3F",
    x"0E844889",
    x"0E8414E7",
    x"0E83E159",
    x"0E83ADDF",
    x"0E837A79",
    x"0E834727",
    x"0E8313E9",
    x"0E82E0BF",
    x"0E82ADAA",
    x"0E827AA8",
    x"0E8247BA",
    x"0E8214E0",
    x"0E81E21A",
    x"0E81AF67",
    x"0E817CC8",
    x"0E814A3E",
    x"0E8117C6",
    x"0E80E563",
    x"0E80B313",
    x"0E8080D7",
    x"0E804EAF",
    x"0E801C9A",
    x"0E7FD530",
    x"0E7F7155",
    x"0E7F0DA0",
    x"0E7EAA12",
    x"0E7E46AB",
    x"0E7DE36B",
    x"0E7D8051",
    x"0E7D1D5F",
    x"0E7CBA92",
    x"0E7C57ED",
    x"0E7BF56E",
    x"0E7B9315",
    x"0E7B30E3",
    x"0E7ACED7",
    x"0E7A6CF1",
    x"0E7A0B32",
    x"0E79A998",
    x"0E794825",
    x"0E78E6D8",
    x"0E7885B1",
    x"0E7824AF",
    x"0E77C3D4",
    x"0E77631E",
    x"0E77028F",
    x"0E76A224",
    x"0E7641E0",
    x"0E75E1C1",
    x"0E7581C8",
    x"0E7521F4",
    x"0E74C245",
    x"0E7462BC",
    x"0E740358",
    x"0E73A419",
    x"0E734500",
    x"0E72E60B",
    x"0E72873C",
    x"0E722892",
    x"0E71CA0C",
    x"0E716BAC",
    x"0E710D70",
    x"0E70AF59",
    x"0E705167",
    x"0E6FF39A",
    x"0E6F95F1",
    x"0E6F386C",
    x"0E6EDB0D",
    x"0E6E7DD1",
    x"0E6E20BA",
    x"0E6DC3C8",
    x"0E6D66F9",
    x"0E6D0A4F",
    x"0E6CADC9",
    x"0E6C5167",
    x"0E6BF52A",
    x"0E6B9910",
    x"0E6B3D1A",
    x"0E6AE148",
    x"0E6A859A",
    x"0E6A2A10",
    x"0E69CEA9",
    x"0E697366",
    x"0E691847",
    x"0E68BD4B",
    x"0E686273",
    x"0E6807BE",
    x"0E67AD2D",
    x"0E6752BF",
    x"0E66F874",
    x"0E669E4D",
    x"0E664449",
    x"0E65EA68",
    x"0E6590A9",
    x"0E65370E",
    x"0E64DD96",
    x"0E648441",
    x"0E642B0F",
    x"0E63D200",
    x"0E637913",
    x"0E632049",
    x"0E62C7A2",
    x"0E626F1D",
    x"0E6216BB",
    x"0E61BE7B",
    x"0E61665E",
    x"0E610E63",
    x"0E60B68B",
    x"0E605ED5",
    x"0E600741",
    x"0E5FAFCF",
    x"0E5F587F",
    x"0E5F0152",
    x"0E5EAA46",
    x"0E5E535D",
    x"0E5DFC95",
    x"0E5DA5EF",
    x"0E5D4F6C",
    x"0E5CF909",
    x"0E5CA2C9",
    x"0E5C4CAA",
    x"0E5BF6AD",
    x"0E5BA0D1",
    x"0E5B4B17",
    x"0E5AF57F",
    x"0E5AA008",
    x"0E5A4AB2",
    x"0E59F57D",
    x"0E59A06A",
    x"0E594B78",
    x"0E58F6A7",
    x"0E58A1F7",
    x"0E584D68",
    x"0E57F8FB",
    x"0E57A4AE",
    x"0E575082",
    x"0E56FC77",
    x"0E56A88D",
    x"0E5654C3",
    x"0E56011B",
    x"0E55AD92",
    x"0E555A2B",
    x"0E5506E4",
    x"0E54B3BD",
    x"0E5460B8",
    x"0E540DD2",
    x"0E53BB0D",
    x"0E536868",
    x"0E5315E3",
    x"0E52C37F",
    x"0E52713A",
    x"0E521F16",
    x"0E51CD12",
    x"0E517B2E",
    x"0E51296A",
    x"0E50D7C6",
    x"0E508641",
    x"0E5034DD",
    x"0E4FE398",
    x"0E4F9273",
    x"0E4F416D",
    x"0E4EF088",
    x"0E4E9FC2",
    x"0E4E4F1B",
    x"0E4DFE94",
    x"0E4DAE2C",
    x"0E4D5DE4",
    x"0E4D0DBB",
    x"0E4CBDB1",
    x"0E4C6DC6",
    x"0E4C1DFB",
    x"0E4BCE4F",
    x"0E4B7EC2",
    x"0E4B2F54",
    x"0E4AE005",
    x"0E4A90D5",
    x"0E4A41C4",
    x"0E49F2D2",
    x"0E49A3FE",
    x"0E495549",
    x"0E4906B3",
    x"0E48B83C",
    x"0E4869E3",
    x"0E481BA9",
    x"0E47CD8E",
    x"0E477F91",
    x"0E4731B2",
    x"0E46E3F2",
    x"0E469650",
    x"0E4648CC",
    x"0E45FB67",
    x"0E45AE20",
    x"0E4560F7",
    x"0E4513EC",
    x"0E44C700",
    x"0E447A31",
    x"0E442D80",
    x"0E43E0ED",
    x"0E439478",
    x"0E434821",
    x"0E42FBE8",
    x"0E42AFCC",
    x"0E4263CF",
    x"0E4217EE",
    x"0E41CC2C",
    x"0E418087",
    x"0E4134FF",
    x"0E40E995",
    x"0E409E49",
    x"0E40531A",
    x"0E400808",
    x"0E3FBD14",
    x"0E3F723C",
    x"0E3F2782",
    x"0E3EDCE5",
    x"0E3E9266",
    x"0E3E4803",
    x"0E3DFDBD",
    x"0E3DB395",
    x"0E3D6989",
    x"0E3D1F9A",
    x"0E3CD5C8",
    x"0E3C8C13",
    x"0E3C427B",
    x"0E3BF8FF",
    x"0E3BAFA0",
    x"0E3B665E",
    x"0E3B1D38",
    x"0E3AD42F",
    x"0E3A8B43",
    x"0E3A4272",
    x"0E39F9BF",
    x"0E39B127",
    x"0E3968AC",
    x"0E39204E",
    x"0E38D80B",
    x"0E388FE5",
    x"0E3847DB",
    x"0E37FFED",
    x"0E37B81B",
    x"0E377065",
    x"0E3728CB",
    x"0E36E14D",
    x"0E3699EB",
    x"0E3652A5",
    x"0E360B7A",
    x"0E35C46C",
    x"0E357D79",
    x"0E3536A2",
    x"0E34EFE6",
    x"0E34A946",
    x"0E3462C2",
    x"0E341C59",
    x"0E33D60C",
    x"0E338FDA",
    x"0E3349C3",
    x"0E3303C8",
    x"0E32BDE8",
    x"0E327824",
    x"0E32327A",
    x"0E31ECEC",
    x"0E31A779",
    x"0E316221",
    x"0E311CE5",
    x"0E30D7C3",
    x"0E3092BC",
    x"0E304DD0",
    x"0E3008FF",
    x"0E2FC449",
    x"0E2F7FAE",
    x"0E2F3B2D",
    x"0E2EF6C8",
    x"0E2EB27D",
    x"0E2E6E4C",
    x"0E2E2A36",
    x"0E2DE63B",
    x"0E2DA25A",
    x"0E2D5E94",
    x"0E2D1AE9",
    x"0E2CD757",
    x"0E2C93E0",
    x"0E2C5084",
    x"0E2C0D41",
    x"0E2BCA19",
    x"0E2B870C",
    x"0E2B4418",
    x"0E2B013E",
    x"0E2ABE7F",
    x"0E2A7BD9",
    x"0E2A394E",
    x"0E29F6DD",
    x"0E29B485",
    x"0E297248",
    x"0E293024",
    x"0E28EE1A",
    x"0E28AC2A",
    x"0E286A54",
    x"0E282897",
    x"0E27E6F4",
    x"0E27A56A",
    x"0E2763FB",
    x"0E2722A4",
    x"0E26E167",
    x"0E26A044",
    x"0E265F3A",
    x"0E261E4A",
    x"0E25DD73",
    x"0E259CB5",
    x"0E255C10",
    x"0E251B85",
    x"0E24DB13",
    x"0E249ABA",
    x"0E245A7A",
    x"0E241A53",
    x"0E23DA45",
    x"0E239A50",
    x"0E235A75",
    x"0E231AB2",
    x"0E22DB08",
    x"0E229B77",
    x"0E225BFE",
    x"0E221C9F",
    x"0E21DD58",
    x"0E219E2A",
    x"0E215F14",
    x"0E212017",
    x"0E20E133",
    x"0E20A268",
    x"0E2063B4",
    x"0E20251A",
    x"0E1FE697",
    x"0E1FA82D",
    x"0E1F69DC",
    x"0E1F2BA3",
    x"0E1EED82",
    x"0E1EAF79",
    x"0E1E7189",
    x"0E1E33B0",
    x"0E1DF5F0",
    x"0E1DB848",
    x"0E1D7AB8",
    x"0E1D3D40",
    x"0E1CFFE0",
    x"0E1CC298",
    x"0E1C8568",
    x"0E1C4850",
    x"0E1C0B50",
    x"0E1BCE67",
    x"0E1B9197",
    x"0E1B54DE",
    x"0E1B183C",
    x"0E1ADBB3",
    x"0E1A9F41",
    x"0E1A62E6",
    x"0E1A26A3",
    x"0E19EA78",
    x"0E19AE64",
    x"0E197268",
    x"0E193683",
    x"0E18FAB5",
    x"0E18BEFF",
    x"0E188360",
    x"0E1847D8",
    x"0E180C68",
    x"0E17D10F",
    x"0E1795CD",
    x"0E175AA2",
    x"0E171F8E",
    x"0E16E491",
    x"0E16A9AB",
    x"0E166EDC",
    x"0E163424",
    x"0E15F984",
    x"0E15BEFA",
    x"0E158486",
    x"0E154A2A",
    x"0E150FE4",
    x"0E14D5B6",
    x"0E149B9D",
    x"0E14619C",
    x"0E1427B1",
    x"0E13EDDD",
    x"0E13B41F",
    x"0E137A78",
    x"0E1340E8",
    x"0E13076E",
    x"0E12CE0A",
    x"0E1294BD",
    x"0E125B86",
    x"0E122265",
    x"0E11E95B",
    x"0E11B067",
    x"0E117789",
    x"0E113EC1",
    x"0E110610",
    x"0E10CD75",
    x"0E1094EF",
    x"0E105C80",
    x"0E102427",
    x"0E0FEBE4",
    x"0E0FB3B7",
    x"0E0F7BA0",
    x"0E0F439E",
    x"0E0F0BB3",
    x"0E0ED3DD",
    x"0E0E9C1D",
    x"0E0E6473",
    x"0E0E2CDF",
    x"0E0DF560",
    x"0E0DBDF7",
    x"0E0D86A4",
    x"0E0D4F66",
    x"0E0D183E",
    x"0E0CE12B",
    x"0E0CAA2E",
    x"0E0C7346",
    x"0E0C3C74",
    x"0E0C05B7",
    x"0E0BCF0F",
    x"0E0B987D",
    x"0E0B6200",
    x"0E0B2B98",
    x"0E0AF546",
    x"0E0ABF09",
    x"0E0A88E1",
    x"0E0A52CE",
    x"0E0A1CD0",
    x"0E09E6E7",
    x"0E09B113",
    x"0E097B55",
    x"0E0945AB",
    x"0E091016",
    x"0E08DA97",
    x"0E08A52C",
    x"0E086FD6",
    x"0E083A94",
    x"0E080568",
    x"0E07D050",
    x"0E079B4D",
    x"0E07665F",
    x"0E073185",
    x"0E06FCC0",
    x"0E06C810",
    x"0E069374",
    x"0E065EEC",
    x"0E062A79",
    x"0E05F61B",
    x"0E05C1D1",
    x"0E058D9C",
    x"0E05597B",
    x"0E05256E",
    x"0E04F175",
    x"0E04BD91",
    x"0E0489C1",
    x"0E045605",
    x"0E04225E",
    x"0E03EECB",
    x"0E03BB4B",
    x"0E0387E0",
    x"0E035489",
    x"0E032146",
    x"0E02EE17",
    x"0E02BAFC",
    x"0E0287F5",
    x"0E025502",
    x"0E022223",
    x"0E01EF57",
    x"0E01BCA0",
    x"0E0189FC",
    x"0E01576C",
    x"0E0124F0",
    x"0E00F287",
    x"0E00C032",
    x"0E008DF1",
    x"0E005BC3",
    x"0E0029A9",
    x"0DFFEF45",
    x"0DFF8B5F",
    x"0DFF27A0",
    x"0DFEC408",
    x"0DFE6097",
    x"0DFDFD4D",
    x"0DFD9A29",
    x"0DFD372D",
    x"0DFCD456",
    x"0DFC71A7",
    x"0DFC0F1D",
    x"0DFBACBB",
    x"0DFB4A7E",
    x"0DFAE869",
    x"0DFA8679",
    x"0DFA24AF",
    x"0DF9C30C",
    x"0DF9618F",
    x"0DF90038",
    x"0DF89F07",
    x"0DF83DFC",
    x"0DF7DD16",
    x"0DF77C57",
    x"0DF71BBD",
    x"0DF6BB49",
    x"0DF65AFB",
    x"0DF5FAD2",
    x"0DF59ACF",
    x"0DF53AF1",
    x"0DF4DB39",
    x"0DF47BA6",
    x"0DF41C38",
    x"0DF3BCF0",
    x"0DF35DCD",
    x"0DF2FECF",
    x"0DF29FF6",
    x"0DF24142",
    x"0DF1E2B3",
    x"0DF18448",
    x"0DF12603",
    x"0DF0C7E3",
    x"0DF069E7",
    x"0DF00C10",
    x"0DEFAE5E",
    x"0DEF50D0",
    x"0DEEF366",
    x"0DEE9622",
    x"0DEE3901",
    x"0DEDDC05",
    x"0DED7F2D",
    x"0DED227A",
    x"0DECC5EA",
    x"0DEC697F",
    x"0DEC0D38",
    x"0DEBB115",
    x"0DEB5515",
    x"0DEAF93A",
    x"0DEA9D83",
    x"0DEA41EF",
    x"0DE9E67F",
    x"0DE98B33",
    x"0DE9300A",
    x"0DE8D505",
    x"0DE87A24",
    x"0DE81F66",
    x"0DE7C4CB",
    x"0DE76A54",
    x"0DE71000",
    x"0DE6B5D0",
    x"0DE65BC2",
    x"0DE601D8",
    x"0DE5A811",
    x"0DE54E6D",
    x"0DE4F4EC",
    x"0DE49B8D",
    x"0DE44252",
    x"0DE3E93A",
    x"0DE39044",
    x"0DE33771",
    x"0DE2DEC0",
    x"0DE28633",
    x"0DE22DC8",
    x"0DE1D57F",
    x"0DE17D59",
    x"0DE12555",
    x"0DE0CD74",
    x"0DE075B5",
    x"0DE01E18",
    x"0DDFC69D",
    x"0DDF6F44",
    x"0DDF180E",
    x"0DDEC0FA",
    x"0DDE6A07",
    x"0DDE1337",
    x"0DDDBC88",
    x"0DDD65FB",
    x"0DDD0F91",
    x"0DDCB947",
    x"0DDC6320",
    x"0DDC0D1A",
    x"0DDBB736",
    x"0DDB6173",
    x"0DDB0BD1",
    x"0DDAB651",
    x"0DDA60F3",
    x"0DDA0BB6",
    x"0DD9B69A",
    x"0DD9619F",
    x"0DD90CC5",
    x"0DD8B80D",
    x"0DD86376",
    x"0DD80EFF",
    x"0DD7BAAA",
    x"0DD76675",
    x"0DD71262",
    x"0DD6BE6F",
    x"0DD66A9D",
    x"0DD616EC",
    x"0DD5C35B",
    x"0DD56FEB",
    x"0DD51C9C",
    x"0DD4C96D",
    x"0DD4765E",
    x"0DD42370",
    x"0DD3D0A3",
    x"0DD37DF5",
    x"0DD32B68",
    x"0DD2D8FB",
    x"0DD286AF",
    x"0DD23482",
    x"0DD1E276",
    x"0DD19089",
    x"0DD13EBD",
    x"0DD0ED10",
    x"0DD09B83",
    x"0DD04A17",
    x"0DCFF8CA",
    x"0DCFA79C",
    x"0DCF568F",
    x"0DCF05A1",
    x"0DCEB4D2",
    x"0DCE6423",
    x"0DCE1394",
    x"0DCDC324",
    x"0DCD72D3",
    x"0DCD22A2",
    x"0DCCD290",
    x"0DCC829E",
    x"0DCC32CA",
    x"0DCBE316",
    x"0DCB9381",
    x"0DCB440B",
    x"0DCAF4B4",
    x"0DCAA57C",
    x"0DCA5662",
    x"0DCA0768",
    x"0DC9B88D",
    x"0DC969D0",
    x"0DC91B32",
    x"0DC8CCB3",
    x"0DC87E52",
    x"0DC83010",
    x"0DC7E1EC",
    x"0DC793E7",
    x"0DC74601",
    x"0DC6F839",
    x"0DC6AA8F",
    x"0DC65D03",
    x"0DC60F96",
    x"0DC5C247",
    x"0DC57516",
    x"0DC52804",
    x"0DC4DB0F",
    x"0DC48E39",
    x"0DC44180",
    x"0DC3F4E5",
    x"0DC3A869",
    x"0DC35C0A",
    x"0DC30FC9",
    x"0DC2C3A6",
    x"0DC277A0",
    x"0DC22BB8",
    x"0DC1DFEE",
    x"0DC19441",
    x"0DC148B2",
    x"0DC0FD40",
    x"0DC0B1EC",
    x"0DC066B5",
    x"0DC01B9C",
    x"0DBFD0A0",
    x"0DBF85C1",
    x"0DBF3AFF",
    x"0DBEF05B",
    x"0DBEA5D3",
    x"0DBE5B69",
    x"0DBE111C",
    x"0DBDC6EC",
    x"0DBD7CD9",
    x"0DBD32E2",
    x"0DBCE909",
    x"0DBC9F4C",
    x"0DBC55AC",
    x"0DBC0C29",
    x"0DBBC2C3",
    x"0DBB7979",
    x"0DBB304C",
    x"0DBAE73B",
    x"0DBA9E47",
    x"0DBA5570",
    x"0DBA0CB4",
    x"0DB9C416",
    x"0DB97B93",
    x"0DB9332D",
    x"0DB8EAE3",
    x"0DB8A2B6",
    x"0DB85AA4",
    x"0DB812AF",
    x"0DB7CAD5",
    x"0DB78318",
    x"0DB73B77",
    x"0DB6F3F2",
    x"0DB6AC88",
    x"0DB6653B",
    x"0DB61E09",
    x"0DB5D6F4",
    x"0DB58FF9",
    x"0DB5491B",
    x"0DB50258",
    x"0DB4BBB1",
    x"0DB47526",
    x"0DB42EB6",
    x"0DB3E861",
    x"0DB3A228",
    x"0DB35C0A",
    x"0DB31608",
    x"0DB2D021",
    x"0DB28A56",
    x"0DB244A5",
    x"0DB1FF10",
    x"0DB1B996",
    x"0DB17437",
    x"0DB12EF3",
    x"0DB0E9CA",
    x"0DB0A4BC",
    x"0DB05FC9",
    x"0DB01AF2",
    x"0DAFD634",
    x"0DAF9192",
    x"0DAF4D0B",
    x"0DAF089E",
    x"0DAEC44C",
    x"0DAE8015",
    x"0DAE3BF8",
    x"0DADF7F6",
    x"0DADB40E",
    x"0DAD7041",
    x"0DAD2C8E",
    x"0DACE8F6",
    x"0DACA578",
    x"0DAC6215",
    x"0DAC1ECC",
    x"0DABDB9D",
    x"0DAB9888",
    x"0DAB558E",
    x"0DAB12AD",
    x"0DAACFE7",
    x"0DAA8D3B",
    x"0DAA4AA9",
    x"0DAA0831",
    x"0DA9C5D2",
    x"0DA9838E",
    x"0DA94164",
    x"0DA8FF53",
    x"0DA8BD5C",
    x"0DA87B7F",
    x"0DA839BC",
    x"0DA7F812",
    x"0DA7B682",
    x"0DA7750B",
    x"0DA733AE",
    x"0DA6F26B",
    x"0DA6B141",
    x"0DA67030",
    x"0DA62F39",
    x"0DA5EE5B",
    x"0DA5AD97",
    x"0DA56CEC",
    x"0DA52C5A",
    x"0DA4EBE1",
    x"0DA4AB82",
    x"0DA46B3B",
    x"0DA42B0E",
    x"0DA3EAFA",
    x"0DA3AAFE",
    x"0DA36B1C",
    x"0DA32B53",
    x"0DA2EBA2",
    x"0DA2AC0A",
    x"0DA26C8C",
    x"0DA22D26",
    x"0DA1EDD8",
    x"0DA1AEA4",
    x"0DA16F88",
    x"0DA13085",
    x"0DA0F19A",
    x"0DA0B2C8",
    x"0DA0740E",
    x"0DA0356D",
    x"0D9FF6E5",
    x"0D9FB874",
    x"0D9F7A1C",
    x"0D9F3BDD",
    x"0D9EFDB6",
    x"0D9EBFA7",
    x"0D9E81B0",
    x"0D9E43D1",
    x"0D9E060B",
    x"0D9DC85D",
    x"0D9D8AC6",
    x"0D9D4D48",
    x"0D9D0FE2",
    x"0D9CD294",
    x"0D9C955D",
    x"0D9C583F",
    x"0D9C1B38",
    x"0D9BDE4A",
    x"0D9BA173",
    x"0D9B64B4",
    x"0D9B280C",
    x"0D9AEB7C",
    x"0D9AAF04",
    x"0D9A72A4",
    x"0D9A365B",
    x"0D99FA29",
    x"0D99BE0F",
    x"0D99820D",
    x"0D994622",
    x"0D990A4E",
    x"0D98CE91",
    x"0D9892EC",
    x"0D98575F",
    x"0D981BE8",
    x"0D97E089",
    x"0D97A541",
    x"0D976A10",
    x"0D972EF6",
    x"0D96F3F3",
    x"0D96B907",
    x"0D967E32",
    x"0D964375",
    x"0D9608CE",
    x"0D95CE3E",
    x"0D9593C5",
    x"0D955962",
    x"0D951F17",
    x"0D94E4E2",
    x"0D94AAC4",
    x"0D9470BD",
    x"0D9436CC",
    x"0D93FCF2",
    x"0D93C32E",
    x"0D938981",
    x"0D934FEB",
    x"0D93166B",
    x"0D92DD01",
    x"0D92A3AE",
    x"0D926A71",
    x"0D92314B",
    x"0D91F83B",
    x"0D91BF41",
    x"0D91865D",
    x"0D914D90",
    x"0D9114D9",
    x"0D90DC38",
    x"0D90A3AD",
    x"0D906B38",
    x"0D9032D9",
    x"0D8FFA90",
    x"0D8FC25D",
    x"0D8F8A40",
    x"0D8F5239",
    x"0D8F1A48",
    x"0D8EE26D",
    x"0D8EAAA7",
    x"0D8E72F7",
    x"0D8E3B5D",
    x"0D8E03D9",
    x"0D8DCC6A",
    x"0D8D9511",
    x"0D8D5DCE",
    x"0D8D26A0",
    x"0D8CEF88",
    x"0D8CB885",
    x"0D8C8197",
    x"0D8C4AC0",
    x"0D8C13FD",
    x"0D8BDD50",
    x"0D8BA6B8",
    x"0D8B7036",
    x"0D8B39C8",
    x"0D8B0370",
    x"0D8ACD2E",
    x"0D8A9700",
    x"0D8A60E8",
    x"0D8A2AE4",
    x"0D89F4F6",
    x"0D89BF1D",
    x"0D898959",
    x"0D8953AA",
    x"0D891E10",
    x"0D88E88A",
    x"0D88B31A",
    x"0D887DBE",
    x"0D884878",
    x"0D881346",
    x"0D87DE29",
    x"0D87A920",
    x"0D87742C",
    x"0D873F4D",
    x"0D870A83",
    x"0D86D5CD",
    x"0D86A12C",
    x"0D866C9F",
    x"0D863827",
    x"0D8603C3",
    x"0D85CF74",
    x"0D859B39",
    x"0D856713",
    x"0D853301",
    x"0D84FF03",
    x"0D84CB19",
    x"0D849744",
    x"0D846383",
    x"0D842FD7",
    x"0D83FC3E",
    x"0D83C8B9",
    x"0D839549",
    x"0D8361ED",
    x"0D832EA5",
    x"0D82FB70",
    x"0D82C850",
    x"0D829544",
    x"0D82624C",
    x"0D822F67",
    x"0D81FC96",
    x"0D81C9DA",
    x"0D819731",
    x"0D81649C",
    x"0D81321A",
    x"0D80FFAC",
    x"0D80CD52",
    x"0D809B0C",
    x"0D8068D9",
    x"0D8036BA",
    x"0D8004AE",
    x"0D7FA56D",
    x"0D7F41A4",
    x"0D7EDE02",
    x"0D7E7A86",
    x"0D7E1732",
    x"0D7DB404",
    x"0D7D50FD",
    x"0D7CEE1D",
    x"0D7C8B63",
    x"0D7C28D0",
    x"0D7BC663",
    x"0D7B641D",
    x"0D7B01FD",
    x"0D7AA003",
    x"0D7A3E30",
    x"0D79DC83",
    x"0D797AFC",
    x"0D79199B",
    x"0D78B860",
    x"0D78574B",
    x"0D77F65B",
    x"0D779592",
    x"0D7734EF",
    x"0D76D471",
    x"0D767419",
    x"0D7613E6",
    x"0D75B3D9",
    x"0D7553F1",
    x"0D74F42F",
    x"0D749493",
    x"0D74351B",
    x"0D73D5C9",
    x"0D73769C",
    x"0D731794",
    x"0D72B8B2",
    x"0D7259F4",
    x"0D71FB5C",
    x"0D719CE8",
    x"0D713E99",
    x"0D70E06F",
    x"0D70826A",
    x"0D702489",
    x"0D6FC6CD",
    x"0D6F6936",
    x"0D6F0BC3",
    x"0D6EAE74",
    x"0D6E514A",
    x"0D6DF445",
    x"0D6D9764",
    x"0D6D3AA7",
    x"0D6CDE0E",
    x"0D6C8199",
    x"0D6C2549",
    x"0D6BC91C",
    x"0D6B6D13",
    x"0D6B112F",
    x"0D6AB56E",
    x"0D6A59D1",
    x"0D69FE58",
    x"0D69A302",
    x"0D6947D0",
    x"0D68ECC2",
    x"0D6891D7",
    x"0D683710",
    x"0D67DC6C",
    x"0D6781EC",
    x"0D67278F",
    x"0D66CD55",
    x"0D66733E",
    x"0D66194B",
    x"0D65BF7B",
    x"0D6565CD",
    x"0D650C43",
    x"0D64B2DC",
    x"0D645997",
    x"0D640076",
    x"0D63A777",
    x"0D634E9B",
    x"0D62F5E2",
    x"0D629D4B",
    x"0D6244D7",
    x"0D61EC85",
    x"0D619456",
    x"0D613C49",
    x"0D60E45F",
    x"0D608C97",
    x"0D6034F1",
    x"0D5FDD6D",
    x"0D5F860C",
    x"0D5F2ECD",
    x"0D5ED7AF",
    x"0D5E80B4",
    x"0D5E29DB",
    x"0D5DD323",
    x"0D5D7C8E",
    x"0D5D261A",
    x"0D5CCFC8",
    x"0D5C7998",
    x"0D5C2389",
    x"0D5BCD9C",
    x"0D5B77D0",
    x"0D5B2226",
    x"0D5ACC9E",
    x"0D5A7736",
    x"0D5A21F0",
    x"0D59CCCC",
    x"0D5977C8",
    x"0D5922E6",
    x"0D58CE25",
    x"0D587985",
    x"0D582506",
    x"0D57D0A8",
    x"0D577C6B",
    x"0D57284F",
    x"0D56D454",
    x"0D568079",
    x"0D562CBF",
    x"0D55D926",
    x"0D5585AE",
    x"0D553256",
    x"0D54DF1E",
    x"0D548C07",
    x"0D543911",
    x"0D53E63B",
    x"0D539385",
    x"0D5340EF",
    x"0D52EE7A",
    x"0D529C25",
    x"0D5249F0",
    x"0D51F7DB",
    x"0D51A5E7",
    x"0D515412",
    x"0D51025D",
    x"0D50B0C8",
    x"0D505F53",
    x"0D500DFD",
    x"0D4FBCC8",
    x"0D4F6BB2",
    x"0D4F1ABC",
    x"0D4EC9E5",
    x"0D4E792E",
    x"0D4E2896",
    x"0D4DD81E",
    x"0D4D87C5",
    x"0D4D378C",
    x"0D4CE772",
    x"0D4C9777",
    x"0D4C479C",
    x"0D4BF7DF",
    x"0D4BA842",
    x"0D4B58C4",
    x"0D4B0965",
    x"0D4ABA24",
    x"0D4A6B03",
    x"0D4A1C01",
    x"0D49CD1D",
    x"0D497E59",
    x"0D492FB3",
    x"0D48E12B",
    x"0D4892C3",
    x"0D484479",
    x"0D47F64D",
    x"0D47A840",
    x"0D475A52",
    x"0D470C82",
    x"0D46BED0",
    x"0D46713D",
    x"0D4623C7",
    x"0D45D671",
    x"0D458938",
    x"0D453C1D",
    x"0D44EF21",
    x"0D44A243",
    x"0D445582",
    x"0D4408E0",
    x"0D43BC5B",
    x"0D436FF5",
    x"0D4323AC",
    x"0D42D781",
    x"0D428B73",
    x"0D423F84",
    x"0D41F3B2",
    x"0D41A7FD",
    x"0D415C66",
    x"0D4110ED",
    x"0D40C591",
    x"0D407A53",
    x"0D402F32",
    x"0D3FE42E",
    x"0D3F9947",
    x"0D3F4E7E",
    x"0D3F03D2",
    x"0D3EB943",
    x"0D3E6ED1",
    x"0D3E247C",
    x"0D3DDA45",
    x"0D3D902A",
    x"0D3D462C",
    x"0D3CFC4B",
    x"0D3CB287",
    x"0D3C68E0",
    x"0D3C1F55",
    x"0D3BD5E7",
    x"0D3B8C96",
    x"0D3B4361",
    x"0D3AFA49",
    x"0D3AB14E",
    x"0D3A686F",
    x"0D3A1FAC",
    x"0D39D706",
    x"0D398E7C",
    x"0D39460F",
    x"0D38FDBD",
    x"0D38B588",
    x"0D386D70",
    x"0D382573",
    x"0D37DD92",
    x"0D3795CE",
    x"0D374E25",
    x"0D370699",
    x"0D36BF28",
    x"0D3677D3",
    x"0D36309A",
    x"0D35E97D",
    x"0D35A27C",
    x"0D355B96",
    x"0D3514CC",
    x"0D34CE1E",
    x"0D34878B",
    x"0D344114",
    x"0D33FAB9",
    x"0D33B478",
    x"0D336E54",
    x"0D33284A",
    x"0D32E25C",
    x"0D329C89",
    x"0D3256D2",
    x"0D321135",
    x"0D31CBB4",
    x"0D31864E",
    x"0D314103",
    x"0D30FBD3",
    x"0D30B6BF",
    x"0D3071C5",
    x"0D302CE6",
    x"0D2FE822",
    x"0D2FA378",
    x"0D2F5EEA",
    x"0D2F1A76",
    x"0D2ED61D",
    x"0D2E91DF",
    x"0D2E4DBB",
    x"0D2E09B2",
    x"0D2DC5C4",
    x"0D2D81F0",
    x"0D2D3E36",
    x"0D2CFA97",
    x"0D2CB712",
    x"0D2C73A8",
    x"0D2C3058",
    x"0D2BED22",
    x"0D2BAA07",
    x"0D2B6705",
    x"0D2B241E",
    x"0D2AE151",
    x"0D2A9E9E",
    x"0D2A5C05",
    x"0D2A1986",
    x"0D29D721",
    x"0D2994D6",
    x"0D2952A5",
    x"0D29108E",
    x"0D28CE90",
    x"0D288CAC",
    x"0D284AE2",
    x"0D280932",
    x"0D27C79B",
    x"0D27861E",
    x"0D2744BA",
    x"0D270370",
    x"0D26C23F",
    x"0D268128",
    x"0D26402A",
    x"0D25FF46",
    x"0D25BE7B",
    x"0D257DC9",
    x"0D253D31",
    x"0D24FCB1",
    x"0D24BC4B",
    x"0D247BFE",
    x"0D243BCA",
    x"0D23FBB0",
    x"0D23BBAE",
    x"0D237BC5",
    x"0D233BF5",
    x"0D22FC3E",
    x"0D22BCA0",
    x"0D227D1B",
    x"0D223DAE",
    x"0D21FE5A",
    x"0D21BF1F",
    x"0D217FFD",
    x"0D2140F3",
    x"0D210202",
    x"0D20C32A",
    x"0D20846A",
    x"0D2045C2",
    x"0D200733",
    x"0D1FC8BD",
    x"0D1F8A5F",
    x"0D1F4C19",
    x"0D1F0DEB",
    x"0D1ECFD6",
    x"0D1E91D9",
    x"0D1E53F4",
    x"0D1E1627",
    x"0D1DD873",
    x"0D1D9AD6",
    x"0D1D5D52",
    x"0D1D1FE5",
    x"0D1CE291",
    x"0D1CA554",
    x"0D1C682F",
    x"0D1C2B23",
    x"0D1BEE2E",
    x"0D1BB151",
    x"0D1B748B",
    x"0D1B37DE",
    x"0D1AFB48",
    x"0D1ABEC9",
    x"0D1A8262",
    x"0D1A4613",
    x"0D1A09DC",
    x"0D19CDBC",
    x"0D1991B3",
    x"0D1955C2",
    x"0D1919E8",
    x"0D18DE26",
    x"0D18A27A",
    x"0D1866E7",
    x"0D182B6A",
    x"0D17F005",
    x"0D17B4B6",
    x"0D17797F",
    x"0D173E60",
    x"0D170357",
    x"0D16C865",
    x"0D168D8A",
    x"0D1652C6",
    x"0D161819",
    x"0D15DD83",
    x"0D15A304",
    x"0D15689C",
    x"0D152E4B",
    x"0D14F410",
    x"0D14B9EC",
    x"0D147FDF",
    x"0D1445E8",
    x"0D140C08",
    x"0D13D23F",
    x"0D13988C",
    x"0D135EEF",
    x"0D13256A",
    x"0D12EBFA",
    x"0D12B2A1",
    x"0D12795F",
    x"0D124032",
    x"0D12071C",
    x"0D11CE1D",
    x"0D119533",
    x"0D115C60",
    x"0D1123A3",
    x"0D10EAFC",
    x"0D10B26C",
    x"0D1079F1",
    x"0D10418C",
    x"0D10093E",
    x"0D0FD105",
    x"0D0F98E2",
    x"0D0F60D6",
    x"0D0F28DF",
    x"0D0EF0FE",
    x"0D0EB933",
    x"0D0E817D",
    x"0D0E49DD",
    x"0D0E1253",
    x"0D0DDADF",
    x"0D0DA380",
    x"0D0D6C37",
    x"0D0D3504",
    x"0D0CFDE6",
    x"0D0CC6DD",
    x"0D0C8FEA",
    x"0D0C590D",
    x"0D0C2245",
    x"0D0BEB92",
    x"0D0BB4F5",
    x"0D0B7E6D",
    x"0D0B47FA",
    x"0D0B119D",
    x"0D0ADB54",
    x"0D0AA521",
    x"0D0A6F03",
    x"0D0A38FA",
    x"0D0A0307",
    x"0D09CD28",
    x"0D09975E",
    x"0D0961AA",
    x"0D092C0A",
    x"0D08F67F",
    x"0D08C10A",
    x"0D088BA9",
    x"0D08565C",
    x"0D082125",
    x"0D07EC03",
    x"0D07B6F5",
    x"0D0781FC",
    x"0D074D17",
    x"0D071847",
    x"0D06E38C",
    x"0D06AEE6",
    x"0D067A54",
    x"0D0645D6",
    x"0D06116D",
    x"0D05DD18",
    x"0D05A8D8",
    x"0D0574AC",
    x"0D054095",
    x"0D050C92",
    x"0D04D8A3",
    x"0D04A4C9",
    x"0D047102",
    x"0D043D50",
    x"0D0409B3",
    x"0D03D629",
    x"0D03A2B3",
    x"0D036F52",
    x"0D033C04",
    x"0D0308CB",
    x"0D02D5A5",
    x"0D02A294",
    x"0D026F96",
    x"0D023CAD",
    x"0D0209D7",
    x"0D01D715",
    x"0D01A467",
    x"0D0171CD",
    x"0D013F46",
    x"0D010CD3",
    x"0D00DA74",
    x"0D00A828",
    x"0D0075F1",
    x"0D0043CC",
    x"0D0011BC",
    x"0CFFBF7D",
    x"0CFF5BAA",
    x"0CFEF7FD",
    x"0CFE9478",
    x"0CFE3119",
    x"0CFDCDE1",
    x"0CFD6AD0",
    x"0CFD07E6",
    x"0CFCA522",
    x"0CFC4285",
    x"0CFBE00E",
    x"0CFB7DBE",
    x"0CFB1B94",
    x"0CFAB990",
    x"0CFA57B3",
    x"0CF9F5FC",
    x"0CF9946B",
    x"0CF93300",
    x"0CF8D1BB",
    x"0CF8709C",
    x"0CF80FA3",
    x"0CF7AED0",
    x"0CF74E22",
    x"0CF6ED9B",
    x"0CF68D39",
    x"0CF62CFC",
    x"0CF5CCE6",
    x"0CF56CF4",
    x"0CF50D28",
    x"0CF4AD82",
    x"0CF44E01",
    x"0CF3EEA5",
    x"0CF38F6E",
    x"0CF3305D",
    x"0CF2D171",
    x"0CF272A9",
    x"0CF21407",
    x"0CF1B58A",
    x"0CF15731",
    x"0CF0F8FD",
    x"0CF09AEF",
    x"0CF03D04",
    x"0CEFDF3F",
    x"0CEF819E",
    x"0CEF2422",
    x"0CEEC6CA",
    x"0CEE6996",
    x"0CEE0C87",
    x"0CEDAF9C",
    x"0CED52D6",
    x"0CECF634",
    x"0CEC99B6",
    x"0CEC3D5C",
    x"0CEBE126",
    x"0CEB8514",
    x"0CEB2926",
    x"0CEACD5C",
    x"0CEA71B5",
    x"0CEA1633",
    x"0CE9BAD4",
    x"0CE95F99",
    x"0CE90481",
    x"0CE8A98D",
    x"0CE84EBD",
    x"0CE7F410",
    x"0CE79986",
    x"0CE73F20",
    x"0CE6E4DD",
    x"0CE68ABD",
    x"0CE630C0",
    x"0CE5D6E7",
    x"0CE57D30",
    x"0CE5239D",
    x"0CE4CA2D",
    x"0CE470DF",
    x"0CE417B4",
    x"0CE3BEAC",
    x"0CE365C7",
    x"0CE30D05",
    x"0CE2B465",
    x"0CE25BE8",
    x"0CE2038D",
    x"0CE1AB55",
    x"0CE1533F",
    x"0CE0FB4C",
    x"0CE0A37B",
    x"0CE04BCC",
    x"0CDFF440",
    x"0CDF9CD6",
    x"0CDF458D",
    x"0CDEEE67",
    x"0CDE9763",
    x"0CDE4081",
    x"0CDDE9C1",
    x"0CDD9322",
    x"0CDD3CA6",
    x"0CDCE64B",
    x"0CDC9012",
    x"0CDC39FA",
    x"0CDBE404",
    x"0CDB8E30",
    x"0CDB387D",
    x"0CDAE2EC",
    x"0CDA8D7C",
    x"0CDA382D",
    x"0CD9E300",
    x"0CD98DF4",
    x"0CD93909",
    x"0CD8E43F",
    x"0CD88F97",
    x"0CD83B0F",
    x"0CD7E6A9",
    x"0CD79263",
    x"0CD73E3E",
    x"0CD6EA3A",
    x"0CD69657",
    x"0CD64295",
    x"0CD5EEF3",
    x"0CD59B72",
    x"0CD54812",
    x"0CD4F4D2",
    x"0CD4A1B3",
    x"0CD44EB4",
    x"0CD3FBD5",
    x"0CD3A917",
    x"0CD35679",
    x"0CD303FB",
    x"0CD2B19E",
    x"0CD25F60",
    x"0CD20D43",
    x"0CD1BB46",
    x"0CD16969",
    x"0CD117AC",
    x"0CD0C60E",
    x"0CD07491",
    x"0CD02333",
    x"0CCFD1F5",
    x"0CCF80D7",
    x"0CCF2FD9",
    x"0CCEDEFA",
    x"0CCE8E3B",
    x"0CCE3D9B",
    x"0CCDED1A",
    x"0CCD9CBA",
    x"0CCD4C78",
    x"0CCCFC56",
    x"0CCCAC53",
    x"0CCC5C6F",
    x"0CCC0CAB",
    x"0CCBBD05",
    x"0CCB6D7F",
    x"0CCB1E18",
    x"0CCACECF",
    x"0CCA7FA6",
    x"0CCA309C",
    x"0CC9E1B0",
    x"0CC992E3",
    x"0CC94435",
    x"0CC8F5A6",
    x"0CC8A735",
    x"0CC858E3",
    x"0CC80AB0",
    x"0CC7BC9B",
    x"0CC76EA5",
    x"0CC720CD",
    x"0CC6D313",
    x"0CC68578",
    x"0CC637FB",
    x"0CC5EA9C",
    x"0CC59D5B",
    x"0CC55039",
    x"0CC50335",
    x"0CC4B64E",
    x"0CC46986",
    x"0CC41CDC",
    x"0CC3D050",
    x"0CC383E1",
    x"0CC33791",
    x"0CC2EB5E",
    x"0CC29F49",
    x"0CC25351",
    x"0CC20778",
    x"0CC1BBBB",
    x"0CC1701D",
    x"0CC1249C",
    x"0CC0D938",
    x"0CC08DF2",
    x"0CC042C9",
    x"0CBFF7BE",
    x"0CBFACD0",
    x"0CBF61FF",
    x"0CBF174B",
    x"0CBECCB5",
    x"0CBE823B",
    x"0CBE37DF",
    x"0CBDEDA0",
    x"0CBDA37D",
    x"0CBD5978",
    x"0CBD0F8F",
    x"0CBCC5C4",
    x"0CBC7C15",
    x"0CBC3283",
    x"0CBBE90D",
    x"0CBB9FB5",
    x"0CBB5679",
    x"0CBB0D59",
    x"0CBAC456",
    x"0CBA7B70",
    x"0CBA32A6",
    x"0CB9E9F8",
    x"0CB9A167",
    x"0CB958F2",
    x"0CB91099",
    x"0CB8C85D",
    x"0CB8803D",
    x"0CB83839",
    x"0CB7F051",
    x"0CB7A885",
    x"0CB760D5",
    x"0CB71941",
    x"0CB6D1CA",
    x"0CB68A6E",
    x"0CB6432D",
    x"0CB5FC09",
    x"0CB5B500",
    x"0CB56E14",
    x"0CB52742",
    x"0CB4E08D",
    x"0CB499F3",
    x"0CB45375",
    x"0CB40D12",
    x"0CB3C6CA",
    x"0CB3809E",
    x"0CB33A8E",
    x"0CB2F499",
    x"0CB2AEBF",
    x"0CB26900",
    x"0CB2235D",
    x"0CB1DDD5",
    x"0CB19867",
    x"0CB15315",
    x"0CB10DDF",
    x"0CB0C8C3",
    x"0CB083C2",
    x"0CB03EDC",
    x"0CAFFA11",
    x"0CAFB560",
    x"0CAF70CB",
    x"0CAF2C50",
    x"0CAEE7F0",
    x"0CAEA3AB",
    x"0CAE5F80",
    x"0CAE1B70",
    x"0CADD77B",
    x"0CAD93A0",
    x"0CAD4FE0",
    x"0CAD0C3A",
    x"0CACC8AE",
    x"0CAC853D",
    x"0CAC41E6",
    x"0CABFEA9",
    x"0CABBB87",
    x"0CAB787F",
    x"0CAB3591",
    x"0CAAF2BD",
    x"0CAAB003",
    x"0CAA6D63",
    x"0CAA2ADE",
    x"0CA9E872",
    x"0CA9A620",
    x"0CA963E8",
    x"0CA921CA",
    x"0CA8DFC6",
    x"0CA89DDB",
    x"0CA85C0A",
    x"0CA81A53",
    x"0CA7D8B6",
    x"0CA79732",
    x"0CA755C8",
    x"0CA71477",
    x"0CA6D340",
    x"0CA69222",
    x"0CA6511D",
    x"0CA61032",
    x"0CA5CF61",
    x"0CA58EA8",
    x"0CA54E09",
    x"0CA50D83",
    x"0CA4CD17",
    x"0CA48CC3",
    x"0CA44C89",
    x"0CA40C67",
    x"0CA3CC5F",
    x"0CA38C70",
    x"0CA34C99",
    x"0CA30CDC",
    x"0CA2CD37",
    x"0CA28DAB",
    x"0CA24E39",
    x"0CA20EDE",
    x"0CA1CF9D",
    x"0CA19074",
    x"0CA15164",
    x"0CA1126D",
    x"0CA0D38E",
    x"0CA094C7",
    x"0CA05619",
    x"0CA01784",
    x"0C9FD907",
    x"0C9F9AA2",
    x"0C9F5C56",
    x"0C9F1E22",
    x"0C9EE007",
    x"0C9EA203",
    x"0C9E6418",
    x"0C9E2645",
    x"0C9DE88A",
    x"0C9DAAE7",
    x"0C9D6D5D",
    x"0C9D2FEA",
    x"0C9CF28F",
    x"0C9CB54C",
    x"0C9C7821",
    x"0C9C3B0E",
    x"0C9BFE13",
    x"0C9BC130",
    x"0C9B8464",
    x"0C9B47B1",
    x"0C9B0B14",
    x"0C9ACE90",
    x"0C9A9223",
    x"0C9A55CE",
    x"0C9A1990",
    x"0C99DD6A",
    x"0C99A15B",
    x"0C996564",
    x"0C992984",
    x"0C98EDBB",
    x"0C98B20A",
    x"0C987670",
    x"0C983AED",
    x"0C97FF82",
    x"0C97C42E",
    x"0C9788F1",
    x"0C974DCB",
    x"0C9712BC",
    x"0C96D7C4",
    x"0C969CE3",
    x"0C96621A",
    x"0C962767",
    x"0C95ECCB",
    x"0C95B246",
    x"0C9577D8",
    x"0C953D80",
    x"0C95033F",
    x"0C94C916",
    x"0C948F02",
    x"0C945506",
    x"0C941B20",
    x"0C93E151",
    x"0C93A798",
    x"0C936DF6",
    x"0C93346A",
    x"0C92FAF5",
    x"0C92C196",
    x"0C92884D",
    x"0C924F1B",
    x"0C921600",
    x"0C91DCFA",
    x"0C91A40B",
    x"0C916B32",
    x"0C91326F",
    x"0C90F9C3",
    x"0C90C12C",
    x"0C9088AC",
    x"0C905041",
    x"0C9017ED",
    x"0C8FDFAF",
    x"0C8FA786",
    x"0C8F6F74",
    x"0C8F3777",
    x"0C8EFF90",
    x"0C8EC7BF",
    x"0C8E9004",
    x"0C8E585F",
    x"0C8E20CF",
    x"0C8DE955",
    x"0C8DB1F1",
    x"0C8D7AA2",
    x"0C8D4369",
    x"0C8D0C46",
    x"0C8CD538",
    x"0C8C9E3F",
    x"0C8C675C",
    x"0C8C308E",
    x"0C8BF9D6",
    x"0C8BC333",
    x"0C8B8CA5",
    x"0C8B562D",
    x"0C8B1FCA",
    x"0C8AE97C",
    x"0C8AB344",
    x"0C8A7D20",
    x"0C8A4712",
    x"0C8A1119",
    x"0C89DB35",
    x"0C89A565",
    x"0C896FAB",
    x"0C893A06",
    x"0C890476",
    x"0C88CEFB",
    x"0C889994",
    x"0C886443",
    x"0C882F06",
    x"0C87F9DE",
    x"0C87C4CB",
    x"0C878FCC",
    x"0C875AE2",
    x"0C87260D",
    x"0C86F14D",
    x"0C86BCA1",
    x"0C868809",
    x"0C865386",
    x"0C861F18",
    x"0C85EABE",
    x"0C85B679",
    x"0C858248",
    x"0C854E2B",
    x"0C851A22",
    x"0C84E62E",
    x"0C84B24F",
    x"0C847E83",
    x"0C844ACC",
    x"0C841729",
    x"0C83E39A",
    x"0C83B01F",
    x"0C837CB8",
    x"0C834965",
    x"0C831627",
    x"0C82E2FC",
    x"0C82AFE5",
    x"0C827CE3",
    x"0C8249F4",
    x"0C821719",
    x"0C81E452",
    x"0C81B19E",
    x"0C817EFF",
    x"0C814C73",
    x"0C8119FB",
    x"0C80E797",
    x"0C80B546",
    x"0C808309",
    x"0C8050E0",
    x"0C801ECA",
    x"0C7FD990",
    x"0C7F75B2",
    x"0C7F11FC",
    x"0C7EAE6C",
    x"0C7E4B03",
    x"0C7DE7C1",
    x"0C7D84A6",
    x"0C7D21B2",
    x"0C7CBEE4",
    x"0C7C5C3D",
    x"0C7BF9BC",
    x"0C7B9762",
    x"0C7B352E",
    x"0C7AD320",
    x"0C7A7139",
    x"0C7A0F77",
    x"0C79ADDD",
    x"0C794C68",
    x"0C78EB19",
    x"0C7889F0",
    x"0C7828ED",
    x"0C77C810",
    x"0C776759",
    x"0C7706C7",
    x"0C76A65B",
    x"0C764615",
    x"0C75E5F5",
    x"0C7585FA",
    x"0C752624",
    x"0C74C674",
    x"0C7466E9",
    x"0C740783",
    x"0C73A843",
    x"0C734928",
    x"0C72EA32",
    x"0C728B61",
    x"0C722CB5",
    x"0C71CE2E",
    x"0C716FCC",
    x"0C71118F",
    x"0C70B376",
    x"0C705582",
    x"0C6FF7B3",
    x"0C6F9A09",
    x"0C6F3C83",
    x"0C6EDF22",
    x"0C6E81E5",
    x"0C6E24CC",
    x"0C6DC7D8",
    x"0C6D6B08",
    x"0C6D0E5C",
    x"0C6CB1D5",
    x"0C6C5571",
    x"0C6BF932",
    x"0C6B9D17",
    x"0C6B411F",
    x"0C6AE54C",
    x"0C6A899C",
    x"0C6A2E10",
    x"0C69D2A8",
    x"0C697763",
    x"0C691C43",
    x"0C68C145",
    x"0C68666C",
    x"0C680BB5",
    x"0C67B122",
    x"0C6756B3",
    x"0C66FC67",
    x"0C66A23E",
    x"0C664838",
    x"0C65EE55",
    x"0C659496",
    x"0C653AF9",
    x"0C64E180",
    x"0C648829",
    x"0C642EF5",
    x"0C63D5E4",
    x"0C637CF6",
    x"0C63242B",
    x"0C62CB82",
    x"0C6272FC",
    x"0C621A98",
    x"0C61C257",
    x"0C616A38",
    x"0C61123C",
    x"0C60BA62",
    x"0C6062AA",
    x"0C600B15",
    x"0C5FB3A2",
    x"0C5F5C50",
    x"0C5F0521",
    x"0C5EAE14",
    x"0C5E5729",
    x"0C5E0060",
    x"0C5DA9B9",
    x"0C5D5334",
    x"0C5CFCD0",
    x"0C5CA68E",
    x"0C5C506E",
    x"0C5BFA6F",
    x"0C5BA492",
    x"0C5B4ED7",
    x"0C5AF93D",
    x"0C5AA3C4",
    x"0C5A4E6D",
    x"0C59F937",
    x"0C59A422",
    x"0C594F2E",
    x"0C58FA5C",
    x"0C58A5AB",
    x"0C58511B",
    x"0C57FCAB",
    x"0C57A85D",
    x"0C575430",
    x"0C570023",
    x"0C56AC38",
    x"0C56586D",
    x"0C5604C3",
    x"0C55B139",
    x"0C555DD0",
    x"0C550A88",
    x"0C54B760",
    x"0C546459",
    x"0C541172",
    x"0C53BEAB",
    x"0C536C05",
    x"0C53197F",
    x"0C52C719",
    x"0C5274D3",
    x"0C5222AD",
    x"0C51D0A8",
    x"0C517EC2",
    x"0C512CFD",
    x"0C50DB57",
    x"0C5089D1",
    x"0C50386C",
    x"0C4FE725",
    x"0C4F95FF",
    x"0C4F44F8",
    x"0C4EF411",
    x"0C4EA349",
    x"0C4E52A1",
    x"0C4E0219",
    x"0C4DB1B0",
    x"0C4D6166",
    x"0C4D113C",
    x"0C4CC131",
    x"0C4C7145",
    x"0C4C2178",
    x"0C4BD1CB",
    x"0C4B823C",
    x"0C4B32CD",
    x"0C4AE37C",
    x"0C4A944B",
    x"0C4A4539",
    x"0C49F645",
    x"0C49A770",
    x"0C4958BA",
    x"0C490A23",
    x"0C48BBAA",
    x"0C486D50",
    x"0C481F15",
    x"0C47D0F8",
    x"0C4782FA",
    x"0C47351A",
    x"0C46E758",
    x"0C4699B5",
    x"0C464C30",
    x"0C45FEC9",
    x"0C45B181",
    x"0C456457",
    x"0C45174A",
    x"0C44CA5C",
    x"0C447D8C",
    x"0C4430DA",
    x"0C43E446",
    x"0C4397D0",
    x"0C434B78",
    x"0C42FF3D",
    x"0C42B320",
    x"0C426721",
    x"0C421B40",
    x"0C41CF7C",
    x"0C4183D5",
    x"0C41384D",
    x"0C40ECE1",
    x"0C40A194",
    x"0C405663",
    x"0C400B50",
    x"0C3FC05A",
    x"0C3F7582",
    x"0C3F2AC6",
    x"0C3EE028",
    x"0C3E95A7",
    x"0C3E4B43",
    x"0C3E00FD",
    x"0C3DB6D3",
    x"0C3D6CC6",
    x"0C3D22D6",
    x"0C3CD902",
    x"0C3C8F4C",
    x"0C3C45B3",
    x"0C3BFC36",
    x"0C3BB2D5",
    x"0C3B6992",
    x"0C3B206B",
    x"0C3AD761",
    x"0C3A8E73",
    x"0C3A45A1",
    x"0C39FCEC",
    x"0C39B454",
    x"0C396BD7",
    x"0C392377",
    x"0C38DB34",
    x"0C38930C",
    x"0C384B01",
    x"0C380312",
    x"0C37BB3E",
    x"0C377387",
    x"0C372BEC",
    x"0C36E46D",
    x"0C369D0A",
    x"0C3655C2",
    x"0C360E97",
    x"0C35C787",
    x"0C358093",
    x"0C3539BA",
    x"0C34F2FE",
    x"0C34AC5C",
    x"0C3465D7",
    x"0C341F6D",
    x"0C33D91E",
    x"0C3392EB",
    x"0C334CD4",
    x"0C3306D7",
    x"0C32C0F6",
    x"0C327B30",
    x"0C323586",
    x"0C31EFF7",
    x"0C31AA82",
    x"0C316529",
    x"0C311FEB",
    x"0C30DAC8",
    x"0C3095C0",
    x"0C3050D3",
    x"0C300C01",
    x"0C2FC74A",
    x"0C2F82AE",
    x"0C2F3E2C",
    x"0C2EF9C5",
    x"0C2EB579",
    x"0C2E7147",
    x"0C2E2D30",
    x"0C2DE934",
    x"0C2DA552",
    x"0C2D618B",
    x"0C2D1DDE",
    x"0C2CDA4B",
    x"0C2C96D3",
    x"0C2C5376",
    x"0C2C1032",
    x"0C2BCD09",
    x"0C2B89FA",
    x"0C2B4705",
    x"0C2B042A",
    x"0C2AC16A",
    x"0C2A7EC3",
    x"0C2A3C37",
    x"0C29F9C4",
    x"0C29B76C",
    x"0C29752D",
    x"0C293308",
    x"0C28F0FD",
    x"0C28AF0C",
    x"0C286D34",
    x"0C282B76",
    x"0C27E9D2",
    x"0C27A848",
    x"0C2766D7",
    x"0C27257F",
    x"0C26E442",
    x"0C26A31D",
    x"0C266212",
    x"0C262120",
    x"0C25E048",
    x"0C259F89",
    x"0C255EE4",
    x"0C251E57",
    x"0C24DDE4",
    x"0C249D8A",
    x"0C245D49",
    x"0C241D21",
    x"0C23DD12",
    x"0C239D1C",
    x"0C235D3F",
    x"0C231D7B",
    x"0C22DDD0",
    x"0C229E3E",
    x"0C225EC5",
    x"0C221F64",
    x"0C21E01C",
    x"0C21A0ED",
    x"0C2161D6",
    x"0C2122D8",
    x"0C20E3F3",
    x"0C20A526",
    x"0C206672",
    x"0C2027D6",
    x"0C1FE953",
    x"0C1FAAE8",
    x"0C1F6C95",
    x"0C1F2E5B",
    x"0C1EF039",
    x"0C1EB22F",
    x"0C1E743E",
    x"0C1E3665",
    x"0C1DF8A3",
    x"0C1DBAFA",
    x"0C1D7D69",
    x"0C1D3FF0",
    x"0C1D028F",
    x"0C1CC546",
    x"0C1C8815",
    x"0C1C4AFC",
    x"0C1C0DFB",
    x"0C1BD111",
    x"0C1B943F",
    x"0C1B5785",
    x"0C1B1AE3",
    x"0C1ADE58",
    x"0C1AA1E5",
    x"0C1A658A",
    x"0C1A2946",
    x"0C19ED19",
    x"0C19B105",
    x"0C197507",
    x"0C193921",
    x"0C18FD52",
    x"0C18C19B",
    x"0C1885FB",
    x"0C184A72",
    x"0C180F01",
    x"0C17D3A7",
    x"0C179864",
    x"0C175D38",
    x"0C172223",
    x"0C16E725",
    x"0C16AC3E",
    x"0C16716E",
    x"0C1636B6",
    x"0C15FC14",
    x"0C15C189",
    x"0C158714",
    x"0C154CB7",
    x"0C151271",
    x"0C14D841",
    x"0C149E28",
    x"0C146425",
    x"0C142A39",
    x"0C13F064",
    x"0C13B6A5",
    x"0C137CFD",
    x"0C13436C",
    x"0C1309F1",
    x"0C12D08C",
    x"0C12973E",
    x"0C125E06",
    x"0C1224E4",
    x"0C11EBD9",
    x"0C11B2E4",
    x"0C117A05",
    x"0C11413D",
    x"0C11088A",
    x"0C10CFEE",
    x"0C109768",
    x"0C105EF8",
    x"0C10269E",
    x"0C0FEE5A",
    x"0C0FB62B",
    x"0C0F7E13",
    x"0C0F4611",
    x"0C0F0E24",
    x"0C0ED64E",
    x"0C0E9E8D",
    x"0C0E66E2",
    x"0C0E2F4D",
    x"0C0DF7CD",
    x"0C0DC063",
    x"0C0D890F",
    x"0C0D51D0",
    x"0C0D1AA7",
    x"0C0CE393",
    x"0C0CAC95",
    x"0C0C75AC",
    x"0C0C3ED9",
    x"0C0C081B",
    x"0C0BD173",
    x"0C0B9AE0",
    x"0C0B6462",
    x"0C0B2DF9",
    x"0C0AF7A6",
    x"0C0AC168",
    x"0C0A8B3F",
    x"0C0A552B",
    x"0C0A1F2C",
    x"0C09E942",
    x"0C09B36E",
    x"0C097DAE",
    x"0C094804",
    x"0C09126E",
    x"0C08DCED",
    x"0C08A781",
    x"0C08722A",
    x"0C083CE8",
    x"0C0807BB",
    x"0C07D2A2",
    x"0C079D9E",
    x"0C0768AF",
    x"0C0733D4",
    x"0C06FF0E",
    x"0C06CA5D",
    x"0C0695C0",
    x"0C066138",
    x"0C062CC4",
    x"0C05F865",
    x"0C05C41A",
    x"0C058FE4",
    x"0C055BC2",
    x"0C0527B4",
    x"0C04F3BB",
    x"0C04BFD6",
    x"0C048C05",
    x"0C045848",
    x"0C0424A0",
    x"0C03F10C",
    x"0C03BD8C",
    x"0C038A20",
    x"0C0356C8",
    x"0C032384",
    x"0C02F054",
    x"0C02BD38",
    x"0C028A30",
    x"0C02573C",
    x"0C02245C",
    x"0C01F190",
    x"0C01BED7",
    x"0C018C33",
    x"0C0159A2",
    x"0C012725",
    x"0C00F4BB",
    x"0C00C265",
    x"0C009023",
    x"0C005DF5",
    x"0C002BDA",
    x"0BFFF3A5",
    x"0BFF8FBD",
    x"0BFF2BFD",
    x"0BFEC863",
    x"0BFE64F0",
    x"0BFE01A4",
    x"0BFD9E7F",
    x"0BFD3B80",
    x"0BFCD8A8",
    x"0BFC75F7",
    x"0BFC136C",
    x"0BFBB108",
    x"0BFB4ECA",
    x"0BFAECB2",
    x"0BFA8AC1",
    x"0BFA28F6",
    x"0BF9C751",
    x"0BF965D2",
    x"0BF90479",
    x"0BF8A347",
    x"0BF8423A",
    x"0BF7E153",
    x"0BF78092",
    x"0BF71FF6",
    x"0BF6BF81",
    x"0BF65F31",
    x"0BF5FF06",
    x"0BF59F01",
    x"0BF53F22",
    x"0BF4DF68",
    x"0BF47FD3",
    x"0BF42064",
    x"0BF3C11A",
    x"0BF361F5",
    x"0BF302F6",
    x"0BF2A41B",
    x"0BF24565",
    x"0BF1E6D5",
    x"0BF18869",
    x"0BF12A22",
    x"0BF0CC00",
    x"0BF06E03",
    x"0BF0102A",
    x"0BEFB276",
    x"0BEF54E7",
    x"0BEEF77C",
    x"0BEE9A35",
    x"0BEE3D13",
    x"0BEDE016",
    x"0BED833C",
    x"0BED2687",
    x"0BECC9F6",
    x"0BEC6D89",
    x"0BEC1140",
    x"0BEBB51C",
    x"0BEB591B",
    x"0BEAFD3E",
    x"0BEAA185",
    x"0BEA45F0",
    x"0BE9EA7E",
    x"0BE98F31",
    x"0BE93407",
    x"0BE8D900",
    x"0BE87E1D",
    x"0BE8235D",
    x"0BE7C8C1",
    x"0BE76E49",
    x"0BE713F3",
    x"0BE6B9C1",
    x"0BE65FB2",
    x"0BE605C6",
    x"0BE5ABFE",
    x"0BE55258",
    x"0BE4F8D5",
    x"0BE49F75",
    x"0BE44639",
    x"0BE3ED1F",
    x"0BE39427",
    x"0BE33B53",
    x"0BE2E2A1",
    x"0BE28A12",
    x"0BE231A5",
    x"0BE1D95B",
    x"0BE18133",
    x"0BE1292E",
    x"0BE0D14B",
    x"0BE0798A",
    x"0BE021EC",
    x"0BDFCA70",
    x"0BDF7316",
    x"0BDF1BDE",
    x"0BDEC4C8",
    x"0BDE6DD4",
    x"0BDE1702",
    x"0BDDC052",
    x"0BDD69C4",
    x"0BDD1358",
    x"0BDCBD0D",
    x"0BDC66E4",
    x"0BDC10DC",
    x"0BDBBAF7",
    x"0BDB6532",
    x"0BDB0F90",
    x"0BDABA0E",
    x"0BDA64AE",
    x"0BDA0F70",
    x"0BD9BA52",
    x"0BD96556",
    x"0BD9107B",
    x"0BD8BBC1",
    x"0BD86728",
    x"0BD812B0",
    x"0BD7BE5A",
    x"0BD76A24",
    x"0BD7160F",
    x"0BD6C21B",
    x"0BD66E47",
    x"0BD61A94",
    x"0BD5C702",
    x"0BD57391",
    x"0BD52040",
    x"0BD4CD10",
    x"0BD47A00",
    x"0BD42710",
    x"0BD3D441",
    x"0BD38192",
    x"0BD32F04",
    x"0BD2DC96",
    x"0BD28A48",
    x"0BD2381A",
    x"0BD1E60C",
    x"0BD1941E",
    x"0BD14250",
    x"0BD0F0A2",
    x"0BD09F14",
    x"0BD04DA6",
    x"0BCFFC57",
    x"0BCFAB29",
    x"0BCF5A1A",
    x"0BCF092A",
    x"0BCEB85A",
    x"0BCE67AA",
    x"0BCE1719",
    x"0BCDC6A8",
    x"0BCD7656",
    x"0BCD2624",
    x"0BCCD610",
    x"0BCC861C",
    x"0BCC3648",
    x"0BCBE692",
    x"0BCB96FB",
    x"0BCB4784",
    x"0BCAF82C",
    x"0BCAA8F2",
    x"0BCA59D8",
    x"0BCA0ADC",
    x"0BC9BBFF",
    x"0BC96D41",
    x"0BC91EA2",
    x"0BC8D021",
    x"0BC881BF",
    x"0BC8337C",
    x"0BC7E557",
    x"0BC79751",
    x"0BC74969",
    x"0BC6FB9F",
    x"0BC6ADF4",
    x"0BC66067",
    x"0BC612F9",
    x"0BC5C5A8",
    x"0BC57876",
    x"0BC52B62",
    x"0BC4DE6C",
    x"0BC49194",
    x"0BC444DB",
    x"0BC3F83F",
    x"0BC3ABC1",
    x"0BC35F60",
    x"0BC3131E",
    x"0BC2C6FA",
    x"0BC27AF3",
    x"0BC22F09",
    x"0BC1E33E",
    x"0BC19790",
    x"0BC14BFF",
    x"0BC1008D",
    x"0BC0B537",
    x"0BC069FF",
    x"0BC01EE4",
    x"0BBFD3E7",
    x"0BBF8907",
    x"0BBF3E44",
    x"0BBEF39E",
    x"0BBEA915",
    x"0BBE5EAA",
    x"0BBE145B",
    x"0BBDCA2A",
    x"0BBD8015",
    x"0BBD361E",
    x"0BBCEC43",
    x"0BBCA285",
    x"0BBC58E4",
    x"0BBC0F60",
    x"0BBBC5F8",
    x"0BBB7CAD",
    x"0BBB337F",
    x"0BBAEA6D",
    x"0BBAA178",
    x"0BBA589F",
    x"0BBA0FE2",
    x"0BB9C742",
    x"0BB97EBF",
    x"0BB93657",
    x"0BB8EE0C",
    x"0BB8A5DD",
    x"0BB85DCB",
    x"0BB815D4",
    x"0BB7CDFA",
    x"0BB7863B",
    x"0BB73E99",
    x"0BB6F712",
    x"0BB6AFA8",
    x"0BB66859",
    x"0BB62126",
    x"0BB5DA0F",
    x"0BB59314",
    x"0BB54C34",
    x"0BB50570",
    x"0BB4BEC8",
    x"0BB4783B",
    x"0BB431CA",
    x"0BB3EB74",
    x"0BB3A53A",
    x"0BB35F1B",
    x"0BB31918",
    x"0BB2D32F",
    x"0BB28D63",
    x"0BB247B1",
    x"0BB2021B",
    x"0BB1BC9F",
    x"0BB1773F",
    x"0BB131FA",
    x"0BB0ECD0",
    x"0BB0A7C1",
    x"0BB062CD",
    x"0BB01DF4",
    x"0BAFD936",
    x"0BAF9492",
    x"0BAF500A",
    x"0BAF0B9C",
    x"0BAEC748",
    x"0BAE8310",
    x"0BAE3EF2",
    x"0BADFAEF",
    x"0BADB706",
    x"0BAD7338",
    x"0BAD2F84",
    x"0BACEBEB",
    x"0BACA86C",
    x"0BAC6507",
    x"0BAC21BD",
    x"0BABDE8D",
    x"0BAB9B77",
    x"0BAB587B",
    x"0BAB159A",
    x"0BAAD2D2",
    x"0BAA9025",
    x"0BAA4D92",
    x"0BAA0B18",
    x"0BA9C8B9",
    x"0BA98674",
    x"0BA94448",
    x"0BA90236",
    x"0BA8C03E",
    x"0BA87E60",
    x"0BA83C9B",
    x"0BA7FAF1",
    x"0BA7B95F",
    x"0BA777E8",
    x"0BA7368A",
    x"0BA6F545",
    x"0BA6B41A",
    x"0BA67308",
    x"0BA63210",
    x"0BA5F131",
    x"0BA5B06C",
    x"0BA56FBF",
    x"0BA52F2C",
    x"0BA4EEB3",
    x"0BA4AE52",
    x"0BA46E0A",
    x"0BA42DDC",
    x"0BA3EDC7",
    x"0BA3ADCA",
    x"0BA36DE7",
    x"0BA32E1C",
    x"0BA2EE6B",
    x"0BA2AED2",
    x"0BA26F52",
    x"0BA22FEB",
    x"0BA1F09D",
    x"0BA1B167",
    x"0BA1724A",
    x"0BA13346",
    x"0BA0F45A",
    x"0BA0B587",
    x"0BA076CC",
    x"0BA0382A",
    x"0B9FF9A0",
    x"0B9FBB2F",
    x"0B9F7CD6",
    x"0B9F3E95",
    x"0B9F006D",
    x"0B9EC25D",
    x"0B9E8465",
    x"0B9E4686",
    x"0B9E08BE",
    x"0B9DCB0F",
    x"0B9D8D78",
    x"0B9D4FF8",
    x"0B9D1291",
    x"0B9CD542",
    x"0B9C980A",
    x"0B9C5AEB",
    x"0B9C1DE3",
    x"0B9BE0F4",
    x"0B9BA41C",
    x"0B9B675B",
    x"0B9B2AB3",
    x"0B9AEE22",
    x"0B9AB1A9",
    x"0B9A7547",
    x"0B9A38FD",
    x"0B99FCCB",
    x"0B99C0B0",
    x"0B9984AC",
    x"0B9948C0",
    x"0B990CEB",
    x"0B98D12E",
    x"0B989588",
    x"0B9859F9",
    x"0B981E82",
    x"0B97E321",
    x"0B97A7D8",
    x"0B976CA6",
    x"0B97318B",
    x"0B96F687",
    x"0B96BB9B",
    x"0B9680C5",
    x"0B964606",
    x"0B960B5E",
    x"0B95D0CD",
    x"0B959653",
    x"0B955BF0",
    x"0B9521A3",
    x"0B94E76D",
    x"0B94AD4E",
    x"0B947346",
    x"0B943954",
    x"0B93FF79",
    x"0B93C5B5",
    x"0B938C07",
    x"0B93526F",
    x"0B9318EE",
    x"0B92DF84",
    x"0B92A630",
    x"0B926CF2",
    x"0B9233CB",
    x"0B91FAB9",
    x"0B91C1BF",
    x"0B9188DA",
    x"0B91500C",
    x"0B911754",
    x"0B90DEB1",
    x"0B90A626",
    x"0B906DB0",
    x"0B903550",
    x"0B8FFD06",
    x"0B8FC4D2",
    x"0B8F8CB4",
    x"0B8F54AC",
    x"0B8F1CBA",
    x"0B8EE4DE",
    x"0B8EAD17",
    x"0B8E7566",
    x"0B8E3DCB",
    x"0B8E0646",
    x"0B8DCED7",
    x"0B8D977D",
    x"0B8D6038",
    x"0B8D2909",
    x"0B8CF1F0",
    x"0B8CBAEC",
    x"0B8C83FE",
    x"0B8C4D25",
    x"0B8C1662",
    x"0B8BDFB4",
    x"0B8BA91B",
    x"0B8B7298",
    x"0B8B3C2A",
    x"0B8B05D1",
    x"0B8ACF8D",
    x"0B8A995E",
    x"0B8A6345",
    x"0B8A2D41",
    x"0B89F752",
    x"0B89C178",
    x"0B898BB3",
    x"0B895603",
    x"0B892067",
    x"0B88EAE1",
    x"0B88B570",
    x"0B888013",
    x"0B884ACC",
    x"0B881599",
    x"0B87E07B",
    x"0B87AB72",
    x"0B87767D",
    x"0B87419D",
    x"0B870CD2",
    x"0B86D81B",
    x"0B86A379",
    x"0B866EEB",
    x"0B863A72",
    x"0B86060E",
    x"0B85D1BD",
    x"0B859D82",
    x"0B85695A",
    x"0B853547",
    x"0B850149",
    x"0B84CD5E",
    x"0B849988",
    x"0B8465C6",
    x"0B843219",
    x"0B83FE7F",
    x"0B83CAFA",
    x"0B839789",
    x"0B83642C",
    x"0B8330E2",
    x"0B82FDAD",
    x"0B82CA8C",
    x"0B82977F",
    x"0B826486",
    x"0B8231A1",
    x"0B81FECF",
    x"0B81CC11",
    x"0B819968",
    x"0B8166D2",
    x"0B81344F",
    x"0B8101E1",
    x"0B80CF86",
    x"0B809D3F",
    x"0B806B0B",
    x"0B8038EB",
    x"0B8006DF",
    x"0B7FA9CB",
    x"0B7F4600",
    x"0B7EE25C",
    x"0B7E7EE0",
    x"0B7E1B89",
    x"0B7DB85A",
    x"0B7D5551",
    x"0B7CF26F",
    x"0B7C8FB4",
    x"0B7C2D1F",
    x"0B7BCAB1",
    x"0B7B6869",
    x"0B7B0647",
    x"0B7AA44C",
    x"0B7A4277",
    x"0B79E0C8",
    x"0B797F3F",
    x"0B791DDC",
    x"0B78BCA0",
    x"0B785B89",
    x"0B77FA98",
    x"0B7799CD",
    x"0B773928",
    x"0B76D8A8",
    x"0B76784F",
    x"0B76181A",
    x"0B75B80C",
    x"0B755823",
    x"0B74F85F",
    x"0B7498C1",
    x"0B743948",
    x"0B73D9F4",
    x"0B737AC5",
    x"0B731BBC",
    x"0B72BCD8",
    x"0B725E18",
    x"0B71FF7E",
    x"0B71A109",
    x"0B7142B8",
    x"0B70E48D",
    x"0B708686",
    x"0B7028A3",
    x"0B6FCAE6",
    x"0B6F6D4D",
    x"0B6F0FD9",
    x"0B6EB289",
    x"0B6E555D",
    x"0B6DF856",
    x"0B6D9B73",
    x"0B6D3EB4",
    x"0B6CE21A",
    x"0B6C85A4",
    x"0B6C2952",
    x"0B6BCD23",
    x"0B6B7119",
    x"0B6B1533",
    x"0B6AB971",
    x"0B6A5DD2",
    x"0B6A0257",
    x"0B69A700",
    x"0B694BCD",
    x"0B68F0BD",
    x"0B6895D1",
    x"0B683B08",
    x"0B67E063",
    x"0B6785E1",
    x"0B672B82",
    x"0B66D147",
    x"0B66772F",
    x"0B661D3A",
    x"0B65C368",
    x"0B6569B9",
    x"0B65102D",
    x"0B64B6C4",
    x"0B645D7E",
    x"0B64045B",
    x"0B63AB5B",
    x"0B63527D",
    x"0B62F9C2",
    x"0B62A12A",
    x"0B6248B4",
    x"0B61F061",
    x"0B619831",
    x"0B614022",
    x"0B60E837",
    x"0B60906D",
    x"0B6038C6",
    x"0B5FE141",
    x"0B5F89DE",
    x"0B5F329D",
    x"0B5EDB7E",
    x"0B5E8481",
    x"0B5E2DA7",
    x"0B5DD6EE",
    x"0B5D8057",
    x"0B5D29E1",
    x"0B5CD38E",
    x"0B5C7D5C",
    x"0B5C274C",
    x"0B5BD15D",
    x"0B5B7B90",
    x"0B5B25E5",
    x"0B5AD05B",
    x"0B5A7AF2",
    x"0B5A25AB",
    x"0B59D085",
    x"0B597B80",
    x"0B59269C",
    x"0B58D1DA",
    x"0B587D38",
    x"0B5828B8",
    x"0B57D458",
    x"0B57801A",
    x"0B572BFC",
    x"0B56D7FF",
    x"0B568423",
    x"0B563068",
    x"0B55DCCE",
    x"0B558954",
    x"0B5535FA",
    x"0B54E2C1",
    x"0B548FA9",
    x"0B543CB1",
    x"0B53E9DA",
    x"0B539723",
    x"0B53448C",
    x"0B52F215",
    x"0B529FBE",
    x"0B524D88",
    x"0B51FB72",
    x"0B51A97C",
    x"0B5157A5",
    x"0B5105EF",
    x"0B50B459",
    x"0B5062E2",
    x"0B50118C",
    x"0B4FC055",
    x"0B4F6F3D",
    x"0B4F1E46",
    x"0B4ECD6E",
    x"0B4E7CB5",
    x"0B4E2C1C",
    x"0B4DDBA3",
    x"0B4D8B49",
    x"0B4D3B0E",
    x"0B4CEAF2",
    x"0B4C9AF6",
    x"0B4C4B19",
    x"0B4BFB5C",
    x"0B4BABBD",
    x"0B4B5C3D",
    x"0B4B0CDD",
    x"0B4ABD9B",
    x"0B4A6E79",
    x"0B4A1F75",
    x"0B49D090",
    x"0B4981CA",
    x"0B493323",
    x"0B48E49A",
    x"0B489630",
    x"0B4847E5",
    x"0B47F9B8",
    x"0B47ABAA",
    x"0B475DBA",
    x"0B470FE8",
    x"0B46C235",
    x"0B4674A1",
    x"0B46272A",
    x"0B45D9D2",
    x"0B458C98",
    x"0B453F7C",
    x"0B44F27E",
    x"0B44A59F",
    x"0B4458DD",
    x"0B440C39",
    x"0B43BFB3",
    x"0B43734B",
    x"0B432701",
    x"0B42DAD5",
    x"0B428EC6",
    x"0B4242D5",
    x"0B41F702",
    x"0B41AB4C",
    x"0B415FB4",
    x"0B41143A",
    x"0B40C8DC",
    x"0B407D9D",
    x"0B40327A",
    x"0B3FE775",
    x"0B3F9C8D",
    x"0B3F51C3",
    x"0B3F0716",
    x"0B3EBC85",
    x"0B3E7212",
    x"0B3E27BC",
    x"0B3DDD83",
    x"0B3D9367",
    x"0B3D4968",
    x"0B3CFF86",
    x"0B3CB5C0",
    x"0B3C6C18",
    x"0B3C228C",
    x"0B3BD91D",
    x"0B3B8FCA",
    x"0B3B4694",
    x"0B3AFD7B",
    x"0B3AB47E",
    x"0B3A6B9E",
    x"0B3A22DA",
    x"0B39DA33",
    x"0B3991A8",
    x"0B394939",
    x"0B3900E7",
    x"0B38B8B0",
    x"0B387096",
    x"0B382898",
    x"0B37E0B7",
    x"0B3798F1",
    x"0B375147",
    x"0B3709B9",
    x"0B36C247",
    x"0B367AF2",
    x"0B3633B7",
    x"0B35EC99",
    x"0B35A597",
    x"0B355EB0",
    x"0B3517E5",
    x"0B34D135",
    x"0B348AA1",
    x"0B344429",
    x"0B33FDCC",
    x"0B33B78A",
    x"0B337164",
    x"0B332B5A",
    x"0B32E56B",
    x"0B329F97",
    x"0B3259DE",
    x"0B321440",
    x"0B31CEBE",
    x"0B318957",
    x"0B31440B",
    x"0B30FEDA",
    x"0B30B9C4",
    x"0B3074C9",
    x"0B302FE8",
    x"0B2FEB23",
    x"0B2FA679",
    x"0B2F61E9",
    x"0B2F1D74",
    x"0B2ED91A",
    x"0B2E94DB",
    x"0B2E50B6",
    x"0B2E0CAB",
    x"0B2DC8BC",
    x"0B2D84E7",
    x"0B2D412C",
    x"0B2CFD8C",
    x"0B2CBA06",
    x"0B2C769A",
    x"0B2C3349",
    x"0B2BF012",
    x"0B2BACF6",
    x"0B2B69F3",
    x"0B2B270B",
    x"0B2AE43D",
    x"0B2AA188",
    x"0B2A5EEE",
    x"0B2A1C6E",
    x"0B29DA08",
    x"0B2997BC",
    x"0B29558A",
    x"0B291371",
    x"0B28D172",
    x"0B288F8D",
    x"0B284DC2",
    x"0B280C11",
    x"0B27CA79",
    x"0B2788FB",
    x"0B274796",
    x"0B27064B",
    x"0B26C519",
    x"0B268401",
    x"0B264302",
    x"0B26021C",
    x"0B25C150",
    x"0B25809D",
    x"0B254004",
    x"0B24FF83",
    x"0B24BF1C",
    x"0B247ECE",
    x"0B243E99",
    x"0B23FE7D",
    x"0B23BE7A",
    x"0B237E90",
    x"0B233EBF",
    x"0B22FF07",
    x"0B22BF68",
    x"0B227FE2",
    x"0B224074",
    x"0B22011F",
    x"0B21C1E3",
    x"0B2182C0",
    x"0B2143B5",
    x"0B2104C3",
    x"0B20C5E9",
    x"0B208728",
    x"0B204880",
    x"0B2009EF",
    x"0B1FCB78",
    x"0B1F8D19",
    x"0B1F4ED2",
    x"0B1F10A3",
    x"0B1ED28D",
    x"0B1E948E",
    x"0B1E56A8",
    x"0B1E18DB",
    x"0B1DDB25",
    x"0B1D9D87",
    x"0B1D6002",
    x"0B1D2294",
    x"0B1CE53F",
    x"0B1CA801",
    x"0B1C6ADC",
    x"0B1C2DCE",
    x"0B1BF0D8",
    x"0B1BB3FA",
    x"0B1B7733",
    x"0B1B3A85",
    x"0B1AFDEE",
    x"0B1AC16E",
    x"0B1A8506",
    x"0B1A48B6",
    x"0B1A0C7E",
    x"0B19D05C",
    x"0B199453",
    x"0B195861",
    x"0B191C86",
    x"0B18E0C2",
    x"0B18A516",
    x"0B186981",
    x"0B182E04",
    x"0B17F29D",
    x"0B17B74E",
    x"0B177C16",
    x"0B1740F5",
    x"0B1705EB",
    x"0B16CAF9",
    x"0B16901D",
    x"0B165558",
    x"0B161AAA",
    x"0B15E013",
    x"0B15A593",
    x"0B156B2A",
    x"0B1530D7",
    x"0B14F69C",
    x"0B14BC77",
    x"0B148268",
    x"0B144871",
    x"0B140E90",
    x"0B13D4C5",
    x"0B139B11",
    x"0B136174",
    x"0B1327ED",
    x"0B12EE7D",
    x"0B12B523",
    x"0B127BDF",
    x"0B1242B2",
    x"0B12099B",
    x"0B11D09B",
    x"0B1197B0",
    x"0B115EDC",
    x"0B11261E",
    x"0B10ED76",
    x"0B10B4E5",
    x"0B107C69",
    x"0B104403",
    x"0B100BB4",
    x"0B0FD37A",
    x"0B0F9B57",
    x"0B0F6349",
    x"0B0F2B51",
    x"0B0EF36F",
    x"0B0EBBA3",
    x"0B0E83EC",
    x"0B0E4C4C",
    x"0B0E14C1",
    x"0B0DDD4C",
    x"0B0DA5EC",
    x"0B0D6EA2",
    x"0B0D376E",
    x"0B0D004F",
    x"0B0CC945",
    x"0B0C9251",
    x"0B0C5B73",
    x"0B0C24AA",
    x"0B0BEDF6",
    x"0B0BB758",
    x"0B0B80CF",
    x"0B0B4A5B",
    x"0B0B13FD",
    x"0B0ADDB4",
    x"0B0AA780",
    x"0B0A7161",
    x"0B0A3B57",
    x"0B0A0563",
    x"0B09CF83",
    x"0B0999B8",
    x"0B096403",
    x"0B092E62",
    x"0B08F8D7",
    x"0B08C360",
    x"0B088DFE",
    x"0B0858B1",
    x"0B082379",
    x"0B07EE55",
    x"0B07B946",
    x"0B07844C",
    x"0B074F67",
    x"0B071A96",
    x"0B06E5DA",
    x"0B06B133",
    x"0B067CA0",
    x"0B064821",
    x"0B0613B7",
    x"0B05DF62",
    x"0B05AB21",
    x"0B0576F4",
    x"0B0542DC",
    x"0B050ED8",
    x"0B04DAE8",
    x"0B04A70D",
    x"0B047346",
    x"0B043F93",
    x"0B040BF4",
    x"0B03D86A",
    x"0B03A4F3",
    x"0B037191",
    x"0B033E42",
    x"0B030B08",
    x"0B02D7E2",
    x"0B02A4CF",
    x"0B0271D1",
    x"0B023EE6",
    x"0B020C10",
    x"0B01D94D",
    x"0B01A69E",
    x"0B017403",
    x"0B01417B",
    x"0B010F08",
    x"0B00DCA8",
    x"0B00AA5B",
    x"0B007823",
    x"0B0045FD",
    x"0B0013EC",
    x"0AFFC3DC",
    x"0AFF6007",
    x"0AFEFC59",
    x"0AFE98D2",
    x"0AFE3571",
    x"0AFDD238",
    x"0AFD6F25",
    x"0AFD0C39",
    x"0AFCA973",
    x"0AFC46D5",
    x"0AFBE45C",
    x"0AFB820A",
    x"0AFB1FDE",
    x"0AFABDD9",
    x"0AFA5BFA",
    x"0AF9FA41",
    x"0AF998AF",
    x"0AF93742",
    x"0AF8D5FB",
    x"0AF874DB",
    x"0AF813E0",
    x"0AF7B30B",
    x"0AF7525C",
    x"0AF6F1D3",
    x"0AF6916F",
    x"0AF63131",
    x"0AF5D119",
    x"0AF57126",
    x"0AF51158",
    x"0AF4B1B0",
    x"0AF4522E",
    x"0AF3F2D0",
    x"0AF39398",
    x"0AF33485",
    x"0AF2D597",
    x"0AF276CE",
    x"0AF2182A",
    x"0AF1B9AB",
    x"0AF15B51",
    x"0AF0FD1C",
    x"0AF09F0B",
    x"0AF0411F",
    x"0AEFE358",
    x"0AEF85B6",
    x"0AEF2838",
    x"0AEECADE",
    x"0AEE6DA9",
    x"0AEE1099",
    x"0AEDB3AC",
    x"0AED56E4",
    x"0AECFA40",
    x"0AEC9DC1",
    x"0AEC4165",
    x"0AEBE52E",
    x"0AEB891A",
    x"0AEB2D2A",
    x"0AEAD15F",
    x"0AEA75B7",
    x"0AEA1A33",
    x"0AE9BED2",
    x"0AE96396",
    x"0AE9087D",
    x"0AE8AD87",
    x"0AE852B5",
    x"0AE7F806",
    x"0AE79D7B",
    x"0AE74313",
    x"0AE6E8CF",
    x"0AE68EAD",
    x"0AE634AF",
    x"0AE5DAD4",
    x"0AE5811C",
    x"0AE52787",
    x"0AE4CE15",
    x"0AE474C6",
    x"0AE41B9A",
    x"0AE3C291",
    x"0AE369AA",
    x"0AE310E6",
    x"0AE2B845",
    x"0AE25FC6",
    x"0AE2076A",
    x"0AE1AF30",
    x"0AE15719",
    x"0AE0FF24",
    x"0AE0A752",
    x"0AE04FA2",
    x"0ADFF814",
    x"0ADFA0A8",
    x"0ADF495E",
    x"0ADEF236",
    x"0ADE9B31",
    x"0ADE444D",
    x"0ADDED8B",
    x"0ADD96EC",
    x"0ADD406E",
    x"0ADCEA11",
    x"0ADC93D7",
    x"0ADC3DBE",
    x"0ADBE7C6",
    x"0ADB91F1",
    x"0ADB3C3C",
    x"0ADAE6AA",
    x"0ADA9138",
    x"0ADA3BE8",
    x"0AD9E6B9",
    x"0AD991AC",
    x"0AD93CBF",
    x"0AD8E7F4",
    x"0AD8934A",
    x"0AD83EC1",
    x"0AD7EA59",
    x"0AD79612",
    x"0AD741EC",
    x"0AD6EDE7",
    x"0AD69A02",
    x"0AD6463E",
    x"0AD5F29B",
    x"0AD59F19",
    x"0AD54BB7",
    x"0AD4F876",
    x"0AD4A555",
    x"0AD45254",
    x"0AD3FF74",
    x"0AD3ACB5",
    x"0AD35A15",
    x"0AD30796",
    x"0AD2B538",
    x"0AD262F9",
    x"0AD210DA",
    x"0AD1BEDC",
    x"0AD16CFD",
    x"0AD11B3E",
    x"0AD0C9A0",
    x"0AD07821",
    x"0AD026C2",
    x"0ACFD583",
    x"0ACF8463",
    x"0ACF3363",
    x"0ACEE283",
    x"0ACE91C2",
    x"0ACE4121",
    x"0ACDF09F",
    x"0ACDA03D",
    x"0ACD4FFA",
    x"0ACCFFD7",
    x"0ACCAFD2",
    x"0ACC5FED",
    x"0ACC1027",
    x"0ACBC081",
    x"0ACB70F9",
    x"0ACB2190",
    x"0ACAD247",
    x"0ACA831C",
    x"0ACA3410",
    x"0AC9E523",
    x"0AC99655",
    x"0AC947A6",
    x"0AC8F915",
    x"0AC8AAA3",
    x"0AC85C50",
    x"0AC80E1B",
    x"0AC7C005",
    x"0AC7720D",
    x"0AC72434",
    x"0AC6D679",
    x"0AC688DC",
    x"0AC63B5E",
    x"0AC5EDFE",
    x"0AC5A0BC",
    x"0AC55398",
    x"0AC50693",
    x"0AC4B9AB",
    x"0AC46CE1",
    x"0AC42036",
    x"0AC3D3A8",
    x"0AC38739",
    x"0AC33AE7",
    x"0AC2EEB2",
    x"0AC2A29C",
    x"0AC256A3",
    x"0AC20AC8",
    x"0AC1BF0B",
    x"0AC1736B",
    x"0AC127E9",
    x"0AC0DC84",
    x"0AC0913D",
    x"0AC04612",
    x"0ABFFB06",
    x"0ABFB016",
    x"0ABF6544",
    x"0ABF1A8F",
    x"0ABECFF7",
    x"0ABE857D",
    x"0ABE3B1F",
    x"0ABDF0DF",
    x"0ABDA6BB",
    x"0ABD5CB4",
    x"0ABD12CA",
    x"0ABCC8FE",
    x"0ABC7F4D",
    x"0ABC35BA",
    x"0ABBEC43",
    x"0ABBA2E9",
    x"0ABB59AC",
    x"0ABB108B",
    x"0ABAC787",
    x"0ABA7EA0",
    x"0ABA35D4",
    x"0AB9ED25",
    x"0AB9A493",
    x"0AB95C1D",
    x"0AB913C3",
    x"0AB8CB85",
    x"0AB88364",
    x"0AB83B5F",
    x"0AB7F376",
    x"0AB7ABA9",
    x"0AB763F7",
    x"0AB71C62",
    x"0AB6D4E9",
    x"0AB68D8C",
    x"0AB6464B",
    x"0AB5FF25",
    x"0AB5B81B",
    x"0AB5712D",
    x"0AB52A5B",
    x"0AB4E3A4",
    x"0AB49D09",
    x"0AB45689",
    x"0AB41025",
    x"0AB3C9DD",
    x"0AB383B0",
    x"0AB33D9E",
    x"0AB2F7A8",
    x"0AB2B1CC",
    x"0AB26C0D",
    x"0AB22668",
    x"0AB1E0DF",
    x"0AB19B70",
    x"0AB1561D",
    x"0AB110E5",
    x"0AB0CBC8",
    x"0AB086C6",
    x"0AB041DF",
    x"0AAFFD12",
    x"0AAFB861",
    x"0AAF73CA",
    x"0AAF2F4E",
    x"0AAEEAED",
    x"0AAEA6A7",
    x"0AAE627B",
    x"0AAE1E6A",
    x"0AADDA73",
    x"0AAD9697",
    x"0AAD52D6",
    x"0AAD0F2F",
    x"0AACCBA2",
    x"0AAC882F",
    x"0AAC44D7",
    x"0AAC019A",
    x"0AABBE76",
    x"0AAB7B6D",
    x"0AAB387E",
    x"0AAAF5A9",
    x"0AAAB2EE",
    x"0AAA704D",
    x"0AAA2DC6",
    x"0AA9EB59",
    x"0AA9A906",
    x"0AA966CD",
    x"0AA924AE",
    x"0AA8E2A8",
    x"0AA8A0BD",
    x"0AA85EEB",
    x"0AA81D33",
    x"0AA7DB94",
    x"0AA79A0F",
    x"0AA758A4",
    x"0AA71752",
    x"0AA6D619",
    x"0AA694FA",
    x"0AA653F5",
    x"0AA61309",
    x"0AA5D236",
    x"0AA5917D",
    x"0AA550DC",
    x"0AA51055",
    x"0AA4CFE8",
    x"0AA48F93",
    x"0AA44F57",
    x"0AA40F35",
    x"0AA3CF2C",
    x"0AA38F3B",
    x"0AA34F64",
    x"0AA30FA5",
    x"0AA2CFFF",
    x"0AA29073",
    x"0AA250FF",
    x"0AA211A3",
    x"0AA1D261",
    x"0AA19337",
    x"0AA15426",
    x"0AA1152D",
    x"0AA0D64D",
    x"0AA09786",
    x"0AA058D7",
    x"0AA01A40",
    x"0A9FDBC2",
    x"0A9F9D5D",
    x"0A9F5F0F",
    x"0A9F20DA",
    x"0A9EE2BE",
    x"0A9EA4B9",
    x"0A9E66CD",
    x"0A9E28F9",
    x"0A9DEB3D",
    x"0A9DAD99",
    x"0A9D700D",
    x"0A9D329A",
    x"0A9CF53E",
    x"0A9CB7FA",
    x"0A9C7ACE",
    x"0A9C3DBA",
    x"0A9C00BE",
    x"0A9BC3D9",
    x"0A9B870D",
    x"0A9B4A58",
    x"0A9B0DBB",
    x"0A9AD135",
    x"0A9A94C7",
    x"0A9A5871",
    x"0A9A1C32",
    x"0A99E00B",
    x"0A99A3FB",
    x"0A996803",
    x"0A992C22",
    x"0A98F058",
    x"0A98B4A6",
    x"0A98790B",
    x"0A983D87",
    x"0A98021B",
    x"0A97C6C6",
    x"0A978B88",
    x"0A975061",
    x"0A971551",
    x"0A96DA58",
    x"0A969F76",
    x"0A9664AB",
    x"0A9629F8",
    x"0A95EF5B",
    x"0A95B4D5",
    x"0A957A65",
    x"0A95400D",
    x"0A9505CB",
    x"0A94CBA0",
    x"0A94918C",
    x"0A94578F",
    x"0A941DA8",
    x"0A93E3D8",
    x"0A93AA1E",
    x"0A93707B",
    x"0A9336EE",
    x"0A92FD78",
    x"0A92C418",
    x"0A928ACE",
    x"0A92519B",
    x"0A92187F",
    x"0A91DF78",
    x"0A91A688",
    x"0A916DAE",
    x"0A9134EA",
    x"0A90FC3D",
    x"0A90C3A5",
    x"0A908B24",
    x"0A9052B9",
    x"0A901A63",
    x"0A8FE224",
    x"0A8FA9FB",
    x"0A8F71E7",
    x"0A8F39EA",
    x"0A8F0202",
    x"0A8ECA30",
    x"0A8E9274",
    x"0A8E5ACE",
    x"0A8E233D",
    x"0A8DEBC2",
    x"0A8DB45D",
    x"0A8D7D0D",
    x"0A8D45D3",
    x"0A8D0EAF",
    x"0A8CD7A0",
    x"0A8CA0A6",
    x"0A8C69C2",
    x"0A8C32F4",
    x"0A8BFC3A",
    x"0A8BC596",
    x"0A8B8F08",
    x"0A8B588F",
    x"0A8B222B",
    x"0A8AEBDC",
    x"0A8AB5A2",
    x"0A8A7F7E",
    x"0A8A496F",
    x"0A8A1375",
    x"0A89DD90",
    x"0A89A7C0",
    x"0A897205",
    x"0A893C5F",
    x"0A8906CD",
    x"0A88D151",
    x"0A889BEA",
    x"0A886697",
    x"0A88315A",
    x"0A87FC31",
    x"0A87C71D",
    x"0A87921D",
    x"0A875D32",
    x"0A87285C",
    x"0A86F39B",
    x"0A86BEEE",
    x"0A868A56",
    x"0A8655D2",
    x"0A862163",
    x"0A85ED08",
    x"0A85B8C2",
    x"0A858490",
    x"0A855072",
    x"0A851C69",
    x"0A84E874",
    x"0A84B493",
    x"0A8480C7",
    x"0A844D0E",
    x"0A84196A",
    x"0A83E5DB",
    x"0A83B25F",
    x"0A837EF7",
    x"0A834BA4",
    x"0A831864",
    x"0A82E539",
    x"0A82B221",
    x"0A827F1D",
    x"0A824C2E",
    x"0A821952",
    x"0A81E68A",
    x"0A81B3D6",
    x"0A818135",
    x"0A814EA9",
    x"0A811C30",
    x"0A80E9CB",
    x"0A80B779",
    x"0A80853B",
    x"0A805311",
    x"0A8020FB",
    x"0A7FDDEF",
    x"0A7F7A10",
    x"0A7F1658",
    x"0A7EB2C6",
    x"0A7E4F5C",
    x"0A7DEC18",
    x"0A7D88FB",
    x"0A7D2605",
    x"0A7CC336",
    x"0A7C608D",
    x"0A7BFE0A",
    x"0A7B9BAE",
    x"0A7B3979",
    x"0A7AD769",
    x"0A7A7580",
    x"0A7A13BD",
    x"0A79B221",
    x"0A7950AA",
    x"0A78EF5A",
    x"0A788E2F",
    x"0A782D2B",
    x"0A77CC4C",
    x"0A776B93",
    x"0A770B00",
    x"0A76AA92",
    x"0A764A4B",
    x"0A75EA28",
    x"0A758A2C",
    x"0A752A54",
    x"0A74CAA3",
    x"0A746B16",
    x"0A740BAF",
    x"0A73AC6D",
    x"0A734D50",
    x"0A72EE58",
    x"0A728F86",
    x"0A7230D8",
    x"0A71D250",
    x"0A7173EC",
    x"0A7115AD",
    x"0A70B793",
    x"0A70599E",
    x"0A6FFBCD",
    x"0A6F9E21",
    x"0A6F4099",
    x"0A6EE336",
    x"0A6E85F8",
    x"0A6E28DE",
    x"0A6DCBE8",
    x"0A6D6F16",
    x"0A6D1269",
    x"0A6CB5E0",
    x"0A6C597B",
    x"0A6BFD3A",
    x"0A6BA11D",
    x"0A6B4524",
    x"0A6AE94F",
    x"0A6A8D9E",
    x"0A6A3211",
    x"0A69D6A7",
    x"0A697B61",
    x"0A69203E",
    x"0A68C540",
    x"0A686A64",
    x"0A680FAC",
    x"0A67B518",
    x"0A675AA7",
    x"0A670059",
    x"0A66A62F",
    x"0A664C27",
    x"0A65F243",
    x"0A659882",
    x"0A653EE4",
    x"0A64E569",
    x"0A648C11",
    x"0A6432DB",
    x"0A63D9C9",
    x"0A6380D9",
    x"0A63280C",
    x"0A62CF62",
    x"0A6276DA",
    x"0A621E75",
    x"0A61C632",
    x"0A616E12",
    x"0A611614",
    x"0A60BE39",
    x"0A606680",
    x"0A600EE9",
    x"0A5FB774",
    x"0A5F6022",
    x"0A5F08F1",
    x"0A5EB1E3",
    x"0A5E5AF6",
    x"0A5E042B",
    x"0A5DAD83",
    x"0A5D56FC",
    x"0A5D0097",
    x"0A5CAA53",
    x"0A5C5432",
    x"0A5BFE32",
    x"0A5BA853",
    x"0A5B5296",
    x"0A5AFCFB",
    x"0A5AA780",
    x"0A5A5228",
    x"0A59FCF0",
    x"0A59A7DA",
    x"0A5952E5",
    x"0A58FE11",
    x"0A58A95F",
    x"0A5854CD",
    x"0A58005C",
    x"0A57AC0D",
    x"0A5757DE",
    x"0A5703D0",
    x"0A56AFE3",
    x"0A565C17",
    x"0A56086B",
    x"0A55B4E0",
    x"0A556176",
    x"0A550E2C",
    x"0A54BB03",
    x"0A5467FA",
    x"0A541511",
    x"0A53C249",
    x"0A536FA2",
    x"0A531D1A",
    x"0A52CAB3",
    x"0A52786C",
    x"0A522645",
    x"0A51D43E",
    x"0A518257",
    x"0A513090",
    x"0A50DEE9",
    x"0A508D62",
    x"0A503BFA",
    x"0A4FEAB3",
    x"0A4F998B",
    x"0A4F4883",
    x"0A4EF79A",
    x"0A4EA6D1",
    x"0A4E5628",
    x"0A4E059E",
    x"0A4DB534",
    x"0A4D64E9",
    x"0A4D14BD",
    x"0A4CC4B0",
    x"0A4C74C3",
    x"0A4C24F5",
    x"0A4BD546",
    x"0A4B85B6",
    x"0A4B3646",
    x"0A4AE6F4",
    x"0A4A97C1",
    x"0A4A48AD",
    x"0A49F9B8",
    x"0A49AAE2",
    x"0A495C2B",
    x"0A490D92",
    x"0A48BF18",
    x"0A4870BD",
    x"0A482280",
    x"0A47D462",
    x"0A478662",
    x"0A473881",
    x"0A46EABE",
    x"0A469D1A",
    x"0A464F93",
    x"0A46022B",
    x"0A45B4E2",
    x"0A4567B6",
    x"0A451AA9",
    x"0A44CDB9",
    x"0A4480E8",
    x"0A443435",
    x"0A43E79F",
    x"0A439B28",
    x"0A434ECE",
    x"0A430292",
    x"0A42B674",
    x"0A426A73",
    x"0A421E91",
    x"0A41D2CC",
    x"0A418724",
    x"0A413B9A",
    x"0A40F02D",
    x"0A40A4DE",
    x"0A4059AD",
    x"0A400E98",
    x"0A3FC3A1",
    x"0A3F78C7",
    x"0A3F2E0B",
    x"0A3EE36B",
    x"0A3E98E9",
    x"0A3E4E84",
    x"0A3E043C",
    x"0A3DBA11",
    x"0A3D7002",
    x"0A3D2611",
    x"0A3CDC3D",
    x"0A3C9285",
    x"0A3C48EA",
    x"0A3BFF6C",
    x"0A3BB60B",
    x"0A3B6CC6",
    x"0A3B239E",
    x"0A3ADA92",
    x"0A3A91A3",
    x"0A3A48D0",
    x"0A3A001A",
    x"0A39B780",
    x"0A396F03",
    x"0A3926A1",
    x"0A38DE5C",
    x"0A389634",
    x"0A384E27",
    x"0A380637",
    x"0A37BE62",
    x"0A3776AA",
    x"0A372F0D",
    x"0A36E78D",
    x"0A36A028",
    x"0A3658E0",
    x"0A3611B3",
    x"0A35CAA2",
    x"0A3583AD",
    x"0A353CD3",
    x"0A34F615",
    x"0A34AF73",
    x"0A3468EC",
    x"0A342281",
    x"0A33DC31",
    x"0A3395FD",
    x"0A334FE4",
    x"0A3309E6",
    x"0A32C404",
    x"0A327E3D",
    x"0A323892",
    x"0A31F301",
    x"0A31AD8C",
    x"0A316831",
    x"0A3122F2",
    x"0A30DDCE",
    x"0A3098C5",
    x"0A3053D7",
    x"0A300F03",
    x"0A2FCA4B",
    x"0A2F85AD",
    x"0A2F412B",
    x"0A2EFCC2",
    x"0A2EB875",
    x"0A2E7442",
    x"0A2E302A",
    x"0A2DEC2D",
    x"0A2DA84A",
    x"0A2D6481",
    x"0A2D20D3",
    x"0A2CDD40",
    x"0A2C99C6",
    x"0A2C5667",
    x"0A2C1323",
    x"0A2BCFF8",
    x"0A2B8CE8",
    x"0A2B49F2",
    x"0A2B0717",
    x"0A2AC455",
    x"0A2A81AD",
    x"0A2A3F1F",
    x"0A29FCAC",
    x"0A29BA52",
    x"0A297812",
    x"0A2935EC",
    x"0A28F3E0",
    x"0A28B1EE",
    x"0A287015",
    x"0A282E56",
    x"0A27ECB1",
    x"0A27AB25",
    x"0A2769B3",
    x"0A27285B",
    x"0A26E71C",
    x"0A26A5F6",
    x"0A2664EA",
    x"0A2623F7",
    x"0A25E31E",
    x"0A25A25E",
    x"0A2561B7",
    x"0A252129",
    x"0A24E0B5",
    x"0A24A05A",
    x"0A246018",
    x"0A241FEF",
    x"0A23DFDF",
    x"0A239FE8",
    x"0A23600A",
    x"0A232045",
    x"0A22E099",
    x"0A22A105",
    x"0A22618B",
    x"0A222229",
    x"0A21E2E0",
    x"0A21A3B0",
    x"0A216498",
    x"0A212599",
    x"0A20E6B3",
    x"0A20A7E5",
    x"0A206930",
    x"0A202A93",
    x"0A1FEC0E",
    x"0A1FADA2",
    x"0A1F6F4F",
    x"0A1F3113",
    x"0A1EF2F0",
    x"0A1EB4E6",
    x"0A1E76F3",
    x"0A1E3919",
    x"0A1DFB56",
    x"0A1DBDAC",
    x"0A1D801A",
    x"0A1D42A0",
    x"0A1D053E",
    x"0A1CC7F4",
    x"0A1C8AC2",
    x"0A1C4DA8",
    x"0A1C10A5",
    x"0A1BD3BB",
    x"0A1B96E8",
    x"0A1B5A2D",
    x"0A1B1D89",
    x"0A1AE0FE",
    x"0A1AA48A",
    x"0A1A682D",
    x"0A1A2BE8",
    x"0A19EFBB",
    x"0A19B3A5",
    x"0A1977A6",
    x"0A193BBF",
    x"0A18FFF0",
    x"0A18C437",
    x"0A188896",
    x"0A184D0D",
    x"0A18119A",
    x"0A17D63F",
    x"0A179AFB",
    x"0A175FCE",
    x"0A1724B8",
    x"0A16E9B9",
    x"0A16AED1",
    x"0A167401",
    x"0A163947",
    x"0A15FEA4",
    x"0A15C418",
    x"0A1589A3",
    x"0A154F44",
    x"0A1514FD",
    x"0A14DACC",
    x"0A14A0B2",
    x"0A1466AE",
    x"0A142CC1",
    x"0A13F2EB",
    x"0A13B92C",
    x"0A137F83",
    x"0A1345F0",
    x"0A130C74",
    x"0A12D30E",
    x"0A1299BF",
    x"0A126086",
    x"0A122764",
    x"0A11EE57",
    x"0A11B561",
    x"0A117C82",
    x"0A1143B8",
    x"0A110B05",
    x"0A10D268",
    x"0A1099E0",
    x"0A10616F",
    x"0A102914",
    x"0A0FF0CF",
    x"0A0FB8A0",
    x"0A0F8087",
    x"0A0F4884",
    x"0A0F1096",
    x"0A0ED8BF",
    x"0A0EA0FD",
    x"0A0E6951",
    x"0A0E31BB",
    x"0A0DFA3A",
    x"0A0DC2CF",
    x"0A0D8B7A",
    x"0A0D543A",
    x"0A0D1D10",
    x"0A0CE5FB",
    x"0A0CAEFC",
    x"0A0C7813",
    x"0A0C413F",
    x"0A0C0A80",
    x"0A0BD3D6",
    x"0A0B9D42",
    x"0A0B66C3",
    x"0A0B305A",
    x"0A0AFA06",
    x"0A0AC3C7",
    x"0A0A8D9D",
    x"0A0A5788",
    x"0A0A2188",
    x"0A09EB9E",
    x"0A09B5C8",
    x"0A098008",
    x"0A094A5C",
    x"0A0914C6",
    x"0A08DF44",
    x"0A08A9D7",
    x"0A08747F",
    x"0A083F3C",
    x"0A080A0E",
    x"0A07D4F4",
    x"0A079FEF",
    x"0A076AFF",
    x"0A073624",
    x"0A07015D",
    x"0A06CCAB",
    x"0A06980D",
    x"0A066384",
    x"0A062F0F",
    x"0A05FAAF",
    x"0A05C664",
    x"0A05922C",
    x"0A055E09",
    x"0A0529FB",
    x"0A04F600",
    x"0A04C21B",
    x"0A048E49",
    x"0A045A8B",
    x"0A0426E2",
    x"0A03F34D",
    x"0A03BFCC",
    x"0A038C5F",
    x"0A035906",
    x"0A0325C2",
    x"0A02F291",
    x"0A02BF74",
    x"0A028C6B",
    x"0A025976",
    x"0A022695",
    x"0A01F3C8",
    x"0A01C10F",
    x"0A018E69",
    x"0A015BD8",
    x"0A01295A",
    x"0A00F6EF",
    x"0A00C499",
    x"0A009256",
    x"0A006026",
    x"0A002E0B",
    x"09FFF805",
    x"09FF941B",
    x"09FF3059",
    x"09FECCBE",
    x"09FE6949",
    x"09FE05FB",
    x"09FDA2D4",
    x"09FD3FD4",
    x"09FCDCFA",
    x"09FC7A47",
    x"09FC17BB",
    x"09FBB555",
    x"09FB5315",
    x"09FAF0FC",
    x"09FA8F09",
    x"09FA2D3C",
    x"09F9CB96",
    x"09F96A15",
    x"09F908BB",
    x"09F8A786",
    x"09F84678",
    x"09F7E58F",
    x"09F784CC",
    x"09F7242F",
    x"09F6C3B8",
    x"09F66366",
    x"09F6033A",
    x"09F5A334",
    x"09F54353",
    x"09F4E397",
    x"09F48401",
    x"09F42490",
    x"09F3C544",
    x"09F3661E",
    x"09F3071D",
    x"09F2A840",
    x"09F24989",
    x"09F1EAF7",
    x"09F18C8A",
    x"09F12E41",
    x"09F0D01D",
    x"09F0721F",
    x"09F01444",
    x"09EFB68F",
    x"09EF58FE",
    x"09EEFB91",
    x"09EE9E49",
    x"09EE4125",
    x"09EDE426",
    x"09ED874B",
    x"09ED2A94",
    x"09ECCE02",
    x"09EC7194",
    x"09EC1549",
    x"09EBB923",
    x"09EB5D21",
    x"09EB0142",
    x"09EAA588",
    x"09EA49F1",
    x"09E9EE7E",
    x"09E9932E",
    x"09E93803",
    x"09E8DCFB",
    x"09E88216",
    x"09E82755",
    x"09E7CCB7",
    x"09E7723D",
    x"09E717E6",
    x"09E6BDB2",
    x"09E663A2",
    x"09E609B5",
    x"09E5AFEA",
    x"09E55643",
    x"09E4FCBF",
    x"09E4A35E",
    x"09E44A1F",
    x"09E3F104",
    x"09E3980B",
    x"09E33F35",
    x"09E2E681",
    x"09E28DF1",
    x"09E23583",
    x"09E1DD37",
    x"09E1850E",
    x"09E12D07",
    x"09E0D523",
    x"09E07D60",
    x"09E025C1",
    x"09DFCE43",
    x"09DF76E7",
    x"09DF1FAE",
    x"09DEC897",
    x"09DE71A1",
    x"09DE1ACE",
    x"09DDC41C",
    x"09DD6D8D",
    x"09DD171F",
    x"09DCC0D3",
    x"09DC6AA8",
    x"09DC149F",
    x"09DBBEB8",
    x"09DB68F2",
    x"09DB134E",
    x"09DABDCB",
    x"09DA686A",
    x"09DA132A",
    x"09D9BE0B",
    x"09D9690D",
    x"09D91431",
    x"09D8BF75",
    x"09D86ADB",
    x"09D81662",
    x"09D7C209",
    x"09D76DD2",
    x"09D719BC",
    x"09D6C5C6",
    x"09D671F1",
    x"09D61E3D",
    x"09D5CAA9",
    x"09D57737",
    x"09D523E4",
    x"09D4D0B3",
    x"09D47DA1",
    x"09D42AB0",
    x"09D3D7E0",
    x"09D38530",
    x"09D332A0",
    x"09D2E030",
    x"09D28DE1",
    x"09D23BB1",
    x"09D1E9A2",
    x"09D197B3",
    x"09D145E3",
    x"09D0F434",
    x"09D0A2A5",
    x"09D05135",
    x"09CFFFE5",
    x"09CFAEB5",
    x"09CF5DA5",
    x"09CF0CB4",
    x"09CEBBE3",
    x"09CE6B31",
    x"09CE1A9F",
    x"09CDCA2C",
    x"09CD79D9",
    x"09CD29A5",
    x"09CCD991",
    x"09CC899B",
    x"09CC39C5",
    x"09CBEA0E",
    x"09CB9A76",
    x"09CB4AFD",
    x"09CAFBA4",
    x"09CAAC69",
    x"09CA5D4D",
    x"09CA0E50",
    x"09C9BF72",
    x"09C970B2",
    x"09C92212",
    x"09C8D390",
    x"09C8852C",
    x"09C836E8",
    x"09C7E8C1",
    x"09C79ABA",
    x"09C74CD0",
    x"09C6FF06",
    x"09C6B159",
    x"09C663CB",
    x"09C6165B",
    x"09C5C90A",
    x"09C57BD6",
    x"09C52EC1",
    x"09C4E1CA",
    x"09C494F0",
    x"09C44835",
    x"09C3FB98",
    x"09C3AF19",
    x"09C362B7",
    x"09C31674",
    x"09C2CA4E",
    x"09C27E45",
    x"09C2325B",
    x"09C1E68E",
    x"09C19ADF",
    x"09C14F4D",
    x"09C103D9",
    x"09C0B882",
    x"09C06D49",
    x"09C0222D",
    x"09BFD72E",
    x"09BF8C4D",
    x"09BF4188",
    x"09BEF6E1",
    x"09BEAC57",
    x"09BE61EB",
    x"09BE179B",
    x"09BDCD68",
    x"09BD8352",
    x"09BD395A",
    x"09BCEF7E",
    x"09BCA5BF",
    x"09BC5C1C",
    x"09BC1297",
    x"09BBC92E",
    x"09BB7FE1",
    x"09BB36B2",
    x"09BAED9F",
    x"09BAA4A8",
    x"09BA5BCE",
    x"09BA1310",
    x"09B9CA6F",
    x"09B981EA",
    x"09B93982",
    x"09B8F135",
    x"09B8A905",
    x"09B860F1",
    x"09B818F9",
    x"09B7D11E",
    x"09B7895E",
    x"09B741BA",
    x"09B6FA33",
    x"09B6B2C7",
    x"09B66B77",
    x"09B62443",
    x"09B5DD2B",
    x"09B5962E",
    x"09B54F4D",
    x"09B50888",
    x"09B4C1DF",
    x"09B47B51",
    x"09B434DE",
    x"09B3EE87",
    x"09B3A84C",
    x"09B3622C",
    x"09B31C27",
    x"09B2D63E",
    x"09B29070",
    x"09B24ABD",
    x"09B20525",
    x"09B1BFA9",
    x"09B17A48",
    x"09B13501",
    x"09B0EFD6",
    x"09B0AAC6",
    x"09B065D1",
    x"09B020F6",
    x"09AFDC37",
    x"09AF9792",
    x"09AF5309",
    x"09AF0E99",
    x"09AECA45",
    x"09AE860B",
    x"09AE41EC",
    x"09ADFDE8",
    x"09ADB9FE",
    x"09AD762F",
    x"09AD327A",
    x"09ACEEDF",
    x"09ACAB5F",
    x"09AC67F9",
    x"09AC24AE",
    x"09ABE17D",
    x"09AB9E66",
    x"09AB5B69",
    x"09AB1886",
    x"09AAD5BE",
    x"09AA930F",
    x"09AA507B",
    x"09AA0E00",
    x"09A9CBA0",
    x"09A98959",
    x"09A9472C",
    x"09A9051A",
    x"09A8C320",
    x"09A88141",
    x"09A83F7B",
    x"09A7FDCF",
    x"09A7BC3D",
    x"09A77AC4",
    x"09A73965",
    x"09A6F820",
    x"09A6B6F3",
    x"09A675E1",
    x"09A634E7",
    x"09A5F407",
    x"09A5B341",
    x"09A57293",
    x"09A531FF",
    x"09A4F184",
    x"09A4B122",
    x"09A470DA",
    x"09A430AA",
    x"09A3F094",
    x"09A3B096",
    x"09A370B2",
    x"09A330E6",
    x"09A2F134",
    x"09A2B19A",
    x"09A27219",
    x"09A232B1",
    x"09A1F361",
    x"09A1B42A",
    x"09A1750C",
    x"09A13607",
    x"09A0F71A",
    x"09A0B846",
    x"09A0798A",
    x"09A03AE7",
    x"099FFC5C",
    x"099FBDEA",
    x"099F7F90",
    x"099F414E",
    x"099F0325",
    x"099EC514",
    x"099E871B",
    x"099E493A",
    x"099E0B72",
    x"099DCDC1",
    x"099D9029",
    x"099D52A8",
    x"099D1540",
    x"099CD7F0",
    x"099C9AB7",
    x"099C5D97",
    x"099C208E",
    x"099BE39E",
    x"099BA6C5",
    x"099B6A03",
    x"099B2D5A",
    x"099AF0C8",
    x"099AB44E",
    x"099A77EB",
    x"099A3BA0",
    x"0999FF6C",
    x"0999C350",
    x"0999874C",
    x"09994B5F",
    x"09990F89",
    x"0998D3CA",
    x"09989823",
    x"09985C94",
    x"0998211B",
    x"0997E5BA",
    x"0997AA70",
    x"09976F3D",
    x"09973421",
    x"0996F91C",
    x"0996BE2E",
    x"09968357",
    x"09964897",
    x"09960DEE",
    x"0995D35C",
    x"099598E1",
    x"09955E7D",
    x"09952430",
    x"0994E9F9",
    x"0994AFD9",
    x"099475CF",
    x"09943BDD",
    x"09940201",
    x"0993C83B",
    x"09938E8C",
    x"099354F4",
    x"09931B72",
    x"0992E206",
    x"0992A8B1",
    x"09926F72",
    x"0992364A",
    x"0991FD38",
    x"0991C43C",
    x"09918B57",
    x"09915287",
    x"099119CE",
    x"0990E12B",
    x"0990A89E",
    x"09907027",
    x"099037C7",
    x"098FFF7C",
    x"098FC747",
    x"098F8F28",
    x"098F571F",
    x"098F1F2C",
    x"098EE74F",
    x"098EAF87",
    x"098E77D6",
    x"098E403A",
    x"098E08B4",
    x"098DD143",
    x"098D99E8",
    x"098D62A3",
    x"098D2B73",
    x"098CF459",
    x"098CBD54",
    x"098C8665",
    x"098C4F8B",
    x"098C18C7",
    x"098BE218",
    x"098BAB7E",
    x"098B74FA",
    x"098B3E8B",
    x"098B0831",
    x"098AD1EC",
    x"098A9BBD",
    x"098A65A3",
    x"098A2F9D",
    x"0989F9AD",
    x"0989C3D2",
    x"09898E0C",
    x"0989585B",
    x"098922BF",
    x"0988ED38",
    x"0988B7C6",
    x"09888269",
    x"09884D20",
    x"098817EC",
    x"0987E2CD",
    x"0987ADC3",
    x"098778CE",
    x"098743ED",
    x"09870F21",
    x"0986DA69",
    x"0986A5C6",
    x"09867137",
    x"09863CBD",
    x"09860858",
    x"0985D407",
    x"09859FCA",
    x"09856BA2",
    x"0985378E",
    x"0985038F",
    x"0984CFA3",
    x"09849BCC",
    x"0984680A",
    x"0984345B",
    x"098400C1",
    x"0983CD3B",
    x"098399C8",
    x"0983666A",
    x"09833320",
    x"0982FFEA",
    x"0982CCC8",
    x"098299BA",
    x"098266C0",
    x"098233DA",
    x"09820108",
    x"0981CE49",
    x"09819B9F",
    x"09816908",
    x"09813685",
    x"09810415",
    x"0980D1B9",
    x"09809F71",
    x"09806D3D",
    x"09803B1C",
    x"0980090F",
    x"097FAE2A",
    x"097F4A5D",
    x"097EE6B8",
    x"097E8339",
    x"097E1FE1",
    x"097DBCB0",
    x"097D59A6",
    x"097CF6C2",
    x"097C9405",
    x"097C316E",
    x"097BCEFE",
    x"097B6CB4",
    x"097B0A91",
    x"097AA894",
    x"097A46BD",
    x"0979E50D",
    x"09798382",
    x"0979221E",
    x"0978C0E0",
    x"09785FC7",
    x"0977FED5",
    x"09779E08",
    x"09773D61",
    x"0976DCE0",
    x"09767C85",
    x"09761C4F",
    x"0975BC3F",
    x"09755C54",
    x"0974FC8F",
    x"09749CEF",
    x"09743D74",
    x"0973DE1F",
    x"09737EEE",
    x"09731FE3",
    x"0972C0FE",
    x"0972623D",
    x"097203A1",
    x"0971A52A",
    x"097146D8",
    x"0970E8AA",
    x"09708AA2",
    x"09702CBE",
    x"096FCEFF",
    x"096F7164",
    x"096F13EE",
    x"096EB69D",
    x"096E5970",
    x"096DFC67",
    x"096D9F82",
    x"096D42C2",
    x"096CE626",
    x"096C89AE",
    x"096C2D5B",
    x"096BD12B",
    x"096B751F",
    x"096B1937",
    x"096ABD74",
    x"096A61D3",
    x"096A0657",
    x"0969AAFE",
    x"09694FC9",
    x"0968F4B8",
    x"096899CA",
    x"09683F00",
    x"0967E459",
    x"096789D6",
    x"09672F75",
    x"0966D538",
    x"09667B1F",
    x"09662128",
    x"0965C755",
    x"09656DA4",
    x"09651417",
    x"0964BAAD",
    x"09646165",
    x"09640841",
    x"0963AF3F",
    x"09635660",
    x"0962FDA3",
    x"0962A50A",
    x"09624C92",
    x"0961F43E",
    x"09619C0C",
    x"096143FC",
    x"0960EC0E",
    x"09609443",
    x"09603C9B",
    x"095FE514",
    x"095F8DB0",
    x"095F366D",
    x"095EDF4D",
    x"095E884F",
    x"095E3173",
    x"095DDAB8",
    x"095D8420",
    x"095D2DA9",
    x"095CD754",
    x"095C8121",
    x"095C2B0F",
    x"095BD51F",
    x"095B7F51",
    x"095B29A4",
    x"095AD418",
    x"095A7EAE",
    x"095A2965",
    x"0959D43D",
    x"09597F37",
    x"09592A52",
    x"0958D58E",
    x"095880EB",
    x"09582C69",
    x"0957D808",
    x"095783C9",
    x"09572FAA",
    x"0956DBAB",
    x"095687CE",
    x"09563411",
    x"0955E075",
    x"09558CFA",
    x"0955399F",
    x"0954E665",
    x"0954934B",
    x"09544052",
    x"0953ED79",
    x"09539AC0",
    x"09534828",
    x"0952F5B0",
    x"0952A358",
    x"09525120",
    x"0951FF08",
    x"0951AD11",
    x"09515B39",
    x"09510982",
    x"0950B7EA",
    x"09506672",
    x"0950151A",
    x"094FC3E1",
    x"094F72C9",
    x"094F21D0",
    x"094ED0F6",
    x"094E803C",
    x"094E2FA2",
    x"094DDF27",
    x"094D8ECC",
    x"094D3E90",
    x"094CEE73",
    x"094C9E75",
    x"094C4E97",
    x"094BFED8",
    x"094BAF38",
    x"094B5FB7",
    x"094B1055",
    x"094AC112",
    x"094A71EE",
    x"094A22E9",
    x"0949D403",
    x"0949853C",
    x"09493693",
    x"0948E809",
    x"0948999E",
    x"09484B51",
    x"0947FD23",
    x"0947AF13",
    x"09476122",
    x"0947134F",
    x"0946C59B",
    x"09467805",
    x"09462A8D",
    x"0945DD34",
    x"09458FF8",
    x"094542DB",
    x"0944F5DC",
    x"0944A8FB",
    x"09445C38",
    x"09440F93",
    x"0943C30C",
    x"094376A3",
    x"09432A57",
    x"0942DE29",
    x"09429219",
    x"09424627",
    x"0941FA53",
    x"0941AE9C",
    x"09416302",
    x"09411786",
    x"0940CC28",
    x"094080E7",
    x"094035C3",
    x"093FEABD",
    x"093F9FD4",
    x"093F5508",
    x"093F0A59",
    x"093EBFC8",
    x"093E7553",
    x"093E2AFC",
    x"093DE0C2",
    x"093D96A5",
    x"093D4CA4",
    x"093D02C1",
    x"093CB8FA",
    x"093C6F50",
    x"093C25C3",
    x"093BDC53",
    x"093B92FF",
    x"093B49C8",
    x"093B00AD",
    x"093AB7AF",
    x"093A6ECE",
    x"093A2609",
    x"0939DD60",
    x"093994D4",
    x"09394C64",
    x"09390410",
    x"0938BBD8",
    x"093873BD",
    x"09382BBE",
    x"0937E3DB",
    x"09379C14",
    x"09375469",
    x"09370CDA",
    x"0936C567",
    x"09367E10",
    x"093636D4",
    x"0935EFB5",
    x"0935A8B1",
    x"093561C9",
    x"09351AFD",
    x"0934D44C",
    x"09348DB7",
    x"0934473D",
    x"093400DF",
    x"0933BA9D",
    x"09337475",
    x"09332E6A",
    x"0932E879",
    x"0932A2A4",
    x"09325CEA",
    x"0932174B",
    x"0931D1C8",
    x"09318C60",
    x"09314712",
    x"093101E0",
    x"0930BCC9",
    x"093077CC",
    x"093032EB",
    x"092FEE25",
    x"092FA979",
    x"092F64E8",
    x"092F2072",
    x"092EDC17",
    x"092E97D6",
    x"092E53B0",
    x"092E0FA5",
    x"092DCBB4",
    x"092D87DE",
    x"092D4422",
    x"092D0080",
    x"092CBCF9",
    x"092C798D",
    x"092C363A",
    x"092BF302",
    x"092BAFE5",
    x"092B6CE1",
    x"092B29F8",
    x"092AE728",
    x"092AA473",
    x"092A61D8",
    x"092A1F56",
    x"0929DCEF",
    x"09299AA2",
    x"0929586E",
    x"09291655",
    x"0928D455",
    x"0928926F",
    x"092850A3",
    x"09280EF0",
    x"0927CD57",
    x"09278BD7",
    x"09274A72",
    x"09270925",
    x"0926C7F2",
    x"092686D9",
    x"092645D9",
    x"092604F2",
    x"0925C425",
    x"09258371",
    x"092542D6",
    x"09250255",
    x"0924C1ED",
    x"0924819D",
    x"09244167",
    x"0924014A",
    x"0923C146",
    x"0923815B",
    x"09234189",
    x"092301D0",
    x"0922C230",
    x"092282A8",
    x"0922433A",
    x"092203E4",
    x"0921C4A7",
    x"09218582",
    x"09214676",
    x"09210783",
    x"0920C8A9",
    x"092089E6",
    x"09204B3D",
    x"09200CAC",
    x"091FCE33",
    x"091F8FD2",
    x"091F518A",
    x"091F135B",
    x"091ED543",
    x"091E9744",
    x"091E595D",
    x"091E1B8E",
    x"091DDDD8",
    x"091DA039",
    x"091D62B2",
    x"091D2544",
    x"091CE7ED",
    x"091CAAAF",
    x"091C6D88",
    x"091C3079",
    x"091BF382",
    x"091BB6A3",
    x"091B79DB",
    x"091B3D2C",
    x"091B0094",
    x"091AC413",
    x"091A87AA",
    x"091A4B59",
    x"091A0F1F",
    x"0919D2FD",
    x"091996F3",
    x"09195AFF",
    x"09191F24",
    x"0918E35F",
    x"0918A7B2",
    x"09186C1C",
    x"0918309D",
    x"0917F536",
    x"0917B9E6",
    x"09177EAD",
    x"0917438B",
    x"09170880",
    x"0916CD8C",
    x"091692AF",
    x"091657EA",
    x"09161D3B",
    x"0915E2A3",
    x"0915A822",
    x"09156DB7",
    x"09153364",
    x"0914F927",
    x"0914BF01",
    x"091484F2",
    x"09144AF9",
    x"09141117",
    x"0913D74C",
    x"09139D97",
    x"091363F9",
    x"09132A71",
    x"0912F100",
    x"0912B7A5",
    x"09127E60",
    x"09124532",
    x"09120C1A",
    x"0911D319",
    x"09119A2D",
    x"09116158",
    x"09112899",
    x"0910EFF0",
    x"0910B75E",
    x"09107EE1",
    x"0910467B",
    x"09100E2A",
    x"090FD5F0",
    x"090F9DCB",
    x"090F65BC",
    x"090F2DC3",
    x"090EF5E0",
    x"090EBE13",
    x"090E865C",
    x"090E4EBA",
    x"090E172E",
    x"090DDFB8",
    x"090DA858",
    x"090D710D",
    x"090D39D7",
    x"090D02B7",
    x"090CCBAD",
    x"090C94B8",
    x"090C5DD9",
    x"090C270F",
    x"090BF05A",
    x"090BB9BB",
    x"090B8331",
    x"090B4CBD",
    x"090B165D",
    x"090AE013",
    x"090AA9DE",
    x"090A73BF",
    x"090A3DB4",
    x"090A07BE",
    x"0909D1DE",
    x"09099C12",
    x"0909665C",
    x"090930BA",
    x"0908FB2E",
    x"0908C5B6",
    x"09089053",
    x"09085B05",
    x"090825CC",
    x"0907F0A8",
    x"0907BB98",
    x"0907869D",
    x"090751B7",
    x"09071CE5",
    x"0906E828",
    x"0906B380",
    x"09067EEC",
    x"09064A6D",
    x"09061602",
    x"0905E1AC",
    x"0905AD6A",
    x"0905793C",
    x"09054523",
    x"0905111E",
    x"0904DD2E",
    x"0904A951",
    x"09047589",
    x"090441D5",
    x"09040E36",
    x"0903DAAA",
    x"0903A733",
    x"090373D0",
    x"09034081",
    x"09030D45",
    x"0902DA1E",
    x"0902A70B",
    x"0902740C",
    x"09024120",
    x"09020E49",
    x"0901DB85",
    x"0901A8D5",
    x"09017639",
    x"090143B1",
    x"0901113C",
    x"0900DEDB",
    x"0900AC8E",
    x"09007A55",
    x"0900482F",
    x"0900161C",
    x"08FFC83B",
    x"08FF6464",
    x"08FF00B4",
    x"08FE9D2B",
    x"08FE39C9",
    x"08FDD68E",
    x"08FD737A",
    x"08FD108C",
    x"08FCADC5",
    x"08FC4B24",
    x"08FBE8AA",
    x"08FB8656",
    x"08FB2429",
    x"08FAC222",
    x"08FA6041",
    x"08F9FE87",
    x"08F99CF3",
    x"08F93B84",
    x"08F8DA3C",
    x"08F8791A",
    x"08F8181D",
    x"08F7B747",
    x"08F75696",
    x"08F6F60B",
    x"08F695A6",
    x"08F63566",
    x"08F5D54C",
    x"08F57558",
    x"08F51588",
    x"08F4B5DF",
    x"08F4565A",
    x"08F3F6FB",
    x"08F397C1",
    x"08F338AD",
    x"08F2D9BD",
    x"08F27AF3",
    x"08F21C4D",
    x"08F1BDCC",
    x"08F15F71",
    x"08F1013A",
    x"08F0A328",
    x"08F0453A",
    x"08EFE772",
    x"08EF89CE",
    x"08EF2C4E",
    x"08EECEF3",
    x"08EE71BC",
    x"08EE14AA",
    x"08EDB7BC",
    x"08ED5AF2",
    x"08ECFE4D",
    x"08ECA1CC",
    x"08EC456F",
    x"08EBE936",
    x"08EB8D20",
    x"08EB312F",
    x"08EAD562",
    x"08EA79B9",
    x"08EA1E33",
    x"08E9C2D1",
    x"08E96793",
    x"08E90C78",
    x"08E8B181",
    x"08E856AD",
    x"08E7FBFD",
    x"08E7A170",
    x"08E74707",
    x"08E6ECC1",
    x"08E6929E",
    x"08E6389E",
    x"08E5DEC2",
    x"08E58508",
    x"08E52B72",
    x"08E4D1FE",
    x"08E478AE",
    x"08E41F80",
    x"08E3C675",
    x"08E36D8D",
    x"08E314C8",
    x"08E2BC25",
    x"08E263A5",
    x"08E20B47",
    x"08E1B30C",
    x"08E15AF3",
    x"08E102FD",
    x"08E0AB29",
    x"08E05377",
    x"08DFFBE7",
    x"08DFA47A",
    x"08DF4D2F",
    x"08DEF606",
    x"08DE9EFF",
    x"08DE481A",
    x"08DDF156",
    x"08DD9AB5",
    x"08DD4435",
    x"08DCEDD8",
    x"08DC979C",
    x"08DC4181",
    x"08DBEB88",
    x"08DB95B1",
    x"08DB3FFB",
    x"08DAEA67",
    x"08DA94F4",
    x"08DA3FA3",
    x"08D9EA73",
    x"08D99564",
    x"08D94076",
    x"08D8EBA9",
    x"08D896FE",
    x"08D84273",
    x"08D7EE0A",
    x"08D799C1",
    x"08D7459A",
    x"08D6F193",
    x"08D69DAD",
    x"08D649E8",
    x"08D5F643",
    x"08D5A2BF",
    x"08D54F5C",
    x"08D4FC19",
    x"08D4A8F7",
    x"08D455F5",
    x"08D40314",
    x"08D3B053",
    x"08D35DB2",
    x"08D30B32",
    x"08D2B8D1",
    x"08D26691",
    x"08D21471",
    x"08D1C271",
    x"08D17091",
    x"08D11ED1",
    x"08D0CD31",
    x"08D07BB1",
    x"08D02A50",
    x"08CFD910",
    x"08CF87EF",
    x"08CF36EE",
    x"08CEE60C",
    x"08CE954A",
    x"08CE44A7",
    x"08CDF424",
    x"08CDA3C1",
    x"08CD537C",
    x"08CD0357",
    x"08CCB352",
    x"08CC636B",
    x"08CC13A4",
    x"08CBC3FC",
    x"08CB7473",
    x"08CB2509",
    x"08CAD5BE",
    x"08CA8692",
    x"08CA3785",
    x"08C9E896",
    x"08C999C7",
    x"08C94B16",
    x"08C8FC84",
    x"08C8AE11",
    x"08C85FBC",
    x"08C81186",
    x"08C7C36F",
    x"08C77576",
    x"08C7279B",
    x"08C6D9DF",
    x"08C68C41",
    x"08C63EC1",
    x"08C5F160",
    x"08C5A41C",
    x"08C556F7",
    x"08C509F0",
    x"08C4BD08",
    x"08C4703D",
    x"08C42390",
    x"08C3D701",
    x"08C38A90",
    x"08C33E3D",
    x"08C2F207",
    x"08C2A5F0",
    x"08C259F6",
    x"08C20E19",
    x"08C1C25B",
    x"08C176B9",
    x"08C12B36",
    x"08C0DFD0",
    x"08C09487",
    x"08C0495C",
    x"08BFFE4E",
    x"08BFB35D",
    x"08BF6889",
    x"08BF1DD3",
    x"08BED33A",
    x"08BE88BE",
    x"08BE3E5F",
    x"08BDF41D",
    x"08BDA9F9",
    x"08BD5FF1",
    x"08BD1606",
    x"08BCCC37",
    x"08BC8286",
    x"08BC38F1",
    x"08BBEF7A",
    x"08BBA61E",
    x"08BB5CE0",
    x"08BB13BE",
    x"08BACAB8",
    x"08BA81CF",
    x"08BA3903",
    x"08B9F053",
    x"08B9A7BF",
    x"08B95F48",
    x"08B916ED",
    x"08B8CEAE",
    x"08B8868B",
    x"08B83E85",
    x"08B7F69A",
    x"08B7AECC",
    x"08B7671A",
    x"08B71F83",
    x"08B6D809",
    x"08B690AB",
    x"08B64968",
    x"08B60241",
    x"08B5BB36",
    x"08B57447",
    x"08B52D73",
    x"08B4E6BC",
    x"08B4A01F",
    x"08B4599E",
    x"08B41339",
    x"08B3CCEF",
    x"08B386C1",
    x"08B340AE",
    x"08B2FAB6",
    x"08B2B4DA",
    x"08B26F19",
    x"08B22973",
    x"08B1E3E9",
    x"08B19E79",
    x"08B15925",
    x"08B113EC",
    x"08B0CECD",
    x"08B089CA",
    x"08B044E2",
    x"08B00014",
    x"08AFBB62",
    x"08AF76CA",
    x"08AF324D",
    x"08AEEDEB",
    x"08AEA9A3",
    x"08AE6576",
    x"08AE2164",
    x"08ADDD6C",
    x"08AD998F",
    x"08AD55CC",
    x"08AD1224",
    x"08ACCE96",
    x"08AC8B22",
    x"08AC47C9",
    x"08AC048A",
    x"08ABC165",
    x"08AB7E5B",
    x"08AB3B6B",
    x"08AAF895",
    x"08AAB5D9",
    x"08AA7336",
    x"08AA30AE",
    x"08A9EE40",
    x"08A9ABEC",
    x"08A969B2",
    x"08A92792",
    x"08A8E58B",
    x"08A8A39E",
    x"08A861CB",
    x"08A82012",
    x"08A7DE72",
    x"08A79CEC",
    x"08A75B80",
    x"08A71A2D",
    x"08A6D8F3",
    x"08A697D3",
    x"08A656CD",
    x"08A615DF",
    x"08A5D50B",
    x"08A59451",
    x"08A553B0",
    x"08A51328",
    x"08A4D2B9",
    x"08A49263",
    x"08A45226",
    x"08A41203",
    x"08A3D1F8",
    x"08A39207",
    x"08A3522E",
    x"08A3126E",
    x"08A2D2C8",
    x"08A2933A",
    x"08A253C5",
    x"08A21468",
    x"08A1D525",
    x"08A195FA",
    x"08A156E7",
    x"08A117EE",
    x"08A0D90D",
    x"08A09A44",
    x"08A05B94",
    x"08A01CFD",
    x"089FDE7E",
    x"089FA017",
    x"089F61C9",
    x"089F2392",
    x"089EE575",
    x"089EA76F",
    x"089E6982",
    x"089E2BAD",
    x"089DEDF0",
    x"089DB04B",
    x"089D72BE",
    x"089D3549",
    x"089CF7EC",
    x"089CBAA7",
    x"089C7D7B",
    x"089C4065",
    x"089C0368",
    x"089BC683",
    x"089B89B5",
    x"089B4CFF",
    x"089B1061",
    x"089AD3DA",
    x"089A976B",
    x"089A5B14",
    x"089A1ED4",
    x"0899E2AC",
    x"0899A69B",
    x"08996AA2",
    x"08992EC0",
    x"0898F2F5",
    x"0898B742",
    x"08987BA6",
    x"08984021",
    x"089804B4",
    x"0897C95E",
    x"08978E1F",
    x"089752F7",
    x"089717E6",
    x"0896DCEC",
    x"0896A209",
    x"0896673D",
    x"08962C89",
    x"0895F1EB",
    x"0895B764",
    x"08957CF3",
    x"0895429A",
    x"08950857",
    x"0894CE2B",
    x"08949416",
    x"08945A18",
    x"08942030",
    x"0893E65F",
    x"0893ACA4",
    x"08937300",
    x"08933972",
    x"0892FFFB",
    x"0892C69A",
    x"08928D50",
    x"0892541C",
    x"08921AFE",
    x"0891E1F6",
    x"0891A905",
    x"0891702A",
    x"08913766",
    x"0890FEB7",
    x"0890C61F",
    x"08908D9C",
    x"08905530",
    x"08901CDA",
    x"088FE499",
    x"088FAC6F",
    x"088F745B",
    x"088F3C5C",
    x"088F0474",
    x"088ECCA1",
    x"088E94E4",
    x"088E5D3C",
    x"088E25AB",
    x"088DEE2F",
    x"088DB6C9",
    x"088D7F78",
    x"088D483D",
    x"088D1118",
    x"088CDA08",
    x"088CA30D",
    x"088C6C28",
    x"088C3559",
    x"088BFE9F",
    x"088BC7FA",
    x"088B916A",
    x"088B5AF0",
    x"088B248B",
    x"088AEE3C",
    x"088AB801",
    x"088A81DC",
    x"088A4BCC",
    x"088A15D1",
    x"0889DFEB",
    x"0889AA1A",
    x"0889745E",
    x"08893EB7",
    x"08890925",
    x"0888D3A8",
    x"08889E3F",
    x"088868EC",
    x"088833AD",
    x"0887FE84",
    x"0887C96F",
    x"0887946E",
    x"08875F83",
    x"08872AAC",
    x"0886F5E9",
    x"0886C13C",
    x"08868CA2",
    x"0886581E",
    x"088623AD",
    x"0885EF52",
    x"0885BB0B",
    x"088586D8",
    x"088552B9",
    x"08851EAF",
    x"0884EAB9",
    x"0884B6D8",
    x"0884830A",
    x"08844F51",
    x"08841BAC",
    x"0883E81C",
    x"0883B49F",
    x"08838136",
    x"08834DE2",
    x"08831AA2",
    x"0882E775",
    x"0882B45D",
    x"08828158",
    x"08824E68",
    x"08821B8B",
    x"0881E8C2",
    x"0881B60D",
    x"0881836C",
    x"088150DF",
    x"08811E65",
    x"0880EBFF",
    x"0880B9AC",
    x"0880876E",
    x"08805543",
    x"0880232B",
    x"087FE24E",
    x"087F7E6D",
    x"087F1AB3",
    x"087EB720",
    x"087E53B4",
    x"087DF06F",
    x"087D8D50",
    x"087D2A59",
    x"087CC787",
    x"087C64DD",
    x"087C0259",
    x"087B9FFB",
    x"087B3DC4",
    x"087ADBB3",
    x"087A79C8",
    x"087A1803",
    x"0879B665",
    x"087954ED",
    x"0878F39B",
    x"0878926F",
    x"08783168",
    x"0877D088",
    x"08776FCD",
    x"08770F39",
    x"0876AEC9",
    x"08764E80",
    x"0875EE5C",
    x"08758E5E",
    x"08752E85",
    x"0874CED1",
    x"08746F43",
    x"08740FDA",
    x"0873B097",
    x"08735178",
    x"0872F27F",
    x"087293AB",
    x"087234FC",
    x"0871D672",
    x"0871780C",
    x"087119CC",
    x"0870BBB0",
    x"08705DB9",
    x"086FFFE7",
    x"086FA239",
    x"086F44B0",
    x"086EE74C",
    x"086E8A0B",
    x"086E2CF0",
    x"086DCFF8",
    x"086D7325",
    x"086D1676",
    x"086CB9EC",
    x"086C5D85",
    x"086C0143",
    x"086BA524",
    x"086B4929",
    x"086AED53",
    x"086A91A0",
    x"086A3611",
    x"0869DAA6",
    x"08697F5E",
    x"0869243A",
    x"0868C93A",
    x"08686E5D",
    x"086813A4",
    x"0867B90E",
    x"08675E9B",
    x"0867044C",
    x"0866AA20",
    x"08665017",
    x"0865F631",
    x"08659C6E",
    x"086542CF",
    x"0864E952",
    x"08648FF9",
    x"086436C2",
    x"0863DDAE",
    x"086384BD",
    x"08632BEE",
    x"0862D342",
    x"08627AB9",
    x"08622252",
    x"0861CA0E",
    x"086171EC",
    x"086119ED",
    x"0860C210",
    x"08606A56",
    x"086012BD",
    x"085FBB47",
    x"085F63F3",
    x"085F0CC1",
    x"085EB5B1",
    x"085E5EC3",
    x"085E07F7",
    x"085DB14D",
    x"085D5AC4",
    x"085D045E",
    x"085CAE19",
    x"085C57F6",
    x"085C01F4",
    x"085BAC14",
    x"085B5656",
    x"085B00B9",
    x"085AAB3D",
    x"085A55E3",
    x"085A00AA",
    x"0859AB92",
    x"0859569C",
    x"085901C7",
    x"0858AD12",
    x"0858587F",
    x"0858040D",
    x"0857AFBC",
    x"08575B8C",
    x"0857077D",
    x"0856B38E",
    x"08565FC0",
    x"08560C13",
    x"0855B887",
    x"0855651B",
    x"085511D0",
    x"0854BEA5",
    x"08546B9B",
    x"085418B1",
    x"0853C5E8",
    x"0853733E",
    x"085320B6",
    x"0852CE4D",
    x"08527C04",
    x"085229DC",
    x"0851D7D4",
    x"085185EB",
    x"08513423",
    x"0850E27B",
    x"085090F2",
    x"08503F89",
    x"084FEE40",
    x"084F9D17",
    x"084F4C0E",
    x"084EFB24",
    x"084EAA59",
    x"084E59AF",
    x"084E0923",
    x"084DB8B8",
    x"084D686B",
    x"084D183E",
    x"084CC830",
    x"084C7842",
    x"084C2872",
    x"084BD8C2",
    x"084B8931",
    x"084B39BF",
    x"084AEA6C",
    x"084A9B38",
    x"084A4C22",
    x"0849FD2C",
    x"0849AE55",
    x"08495F9C",
    x"08491102",
    x"0848C287",
    x"0848742A",
    x"084825EC",
    x"0847D7CC",
    x"084789CB",
    x"08473BE9",
    x"0846EE24",
    x"0846A07E",
    x"084652F7",
    x"0846058E",
    x"0845B843",
    x"08456B16",
    x"08451E07",
    x"0844D116",
    x"08448444",
    x"0844378F",
    x"0843EAF8",
    x"08439E7F",
    x"08435224",
    x"084305E7",
    x"0842B9C8",
    x"08426DC6",
    x"084221E2",
    x"0841D61B",
    x"08418A73",
    x"08413EE7",
    x"0840F379",
    x"0840A829",
    x"08405CF6",
    x"084011E0",
    x"083FC6E8",
    x"083F7C0D",
    x"083F314F",
    x"083EE6AE",
    x"083E9C2B",
    x"083E51C4",
    x"083E077B",
    x"083DBD4F",
    x"083D733F",
    x"083D294D",
    x"083CDF77",
    x"083C95BE",
    x"083C4C22",
    x"083C02A2",
    x"083BB940",
    x"083B6FFA",
    x"083B26D0",
    x"083ADDC3",
    x"083A94D3",
    x"083A4BFF",
    x"083A0348",
    x"0839BAAC",
    x"0839722E",
    x"083929CB",
    x"0838E185",
    x"0838995B",
    x"0838514D",
    x"0838095C",
    x"0837C186",
    x"083779CC",
    x"0837322F",
    x"0836EAAD",
    x"0836A347",
    x"08365BFE",
    x"083614D0",
    x"0835CDBD",
    x"083586C7",
    x"08353FEC",
    x"0834F92D",
    x"0834B289",
    x"08346C01",
    x"08342595",
    x"0833DF44",
    x"0833990E",
    x"083352F4",
    x"08330CF6",
    x"0832C712",
    x"0832814A",
    x"08323B9D",
    x"0831F60B",
    x"0831B095",
    x"08316B3A",
    x"083125F9",
    x"0830E0D4",
    x"08309BCA",
    x"083056DA",
    x"08301206",
    x"082FCD4C",
    x"082F88AD",
    x"082F4429",
    x"082EFFC0",
    x"082EBB71",
    x"082E773E",
    x"082E3324",
    x"082DEF26",
    x"082DAB41",
    x"082D6778",
    x"082D23C9",
    x"082CE034",
    x"082C9CB9",
    x"082C5959",
    x"082C1614",
    x"082BD2E8",
    x"082B8FD7",
    x"082B4CE0",
    x"082B0A03",
    x"082AC740",
    x"082A8497",
    x"082A4208",
    x"0829FF93",
    x"0829BD39",
    x"08297AF8",
    x"082938D0",
    x"0828F6C3",
    x"0828B4D0",
    x"082872F6",
    x"08283136",
    x"0827EF8F",
    x"0827AE03",
    x"08276C90",
    x"08272B36",
    x"0826E9F6",
    x"0826A8CF",
    x"082667C2",
    x"082626CE",
    x"0825E5F4",
    x"0825A532",
    x"0825648A",
    x"082523FC",
    x"0824E386",
    x"0824A32A",
    x"082462E7",
    x"082422BD",
    x"0823E2AC",
    x"0823A2B4",
    x"082362D5",
    x"0823230E",
    x"0822E361",
    x"0822A3CD",
    x"08226451",
    x"082224EE",
    x"0821E5A4",
    x"0821A673",
    x"0821675A",
    x"0821285A",
    x"0820E973",
    x"0820AAA4",
    x"08206BED",
    x"08202D4F",
    x"081FEECA",
    x"081FB05D",
    x"081F7208",
    x"081F33CC",
    x"081EF5A8",
    x"081EB79C",
    x"081E79A8",
    x"081E3BCD",
    x"081DFE0A",
    x"081DC05E",
    x"081D82CB",
    x"081D4550",
    x"081D07ED",
    x"081CCAA2",
    x"081C8D6F",
    x"081C5053",
    x"081C1350",
    x"081BD664",
    x"081B9990",
    x"081B5CD4",
    x"081B2030",
    x"081AE3A3",
    x"081AA72E",
    x"081A6AD1",
    x"081A2E8B",
    x"0819F25C",
    x"0819B645",
    x"08197A46",
    x"08193E5E",
    x"0819028D",
    x"0818C6D4",
    x"08188B32",
    x"08184FA7",
    x"08181433",
    x"0817D8D7",
    x"08179D92",
    x"08176264",
    x"0817274D",
    x"0816EC4D",
    x"0816B165",
    x"08167693",
    x"08163BD8",
    x"08160134",
    x"0815C6A7",
    x"08158C31",
    x"081551D1",
    x"08151789",
    x"0814DD57",
    x"0814A33C",
    x"08146937",
    x"08142F4A",
    x"0813F573",
    x"0813BBB2",
    x"08138208",
    x"08134874",
    x"08130EF7",
    x"0812D591",
    x"08129C40",
    x"08126307",
    x"081229E3",
    x"0811F0D6",
    x"0811B7DF",
    x"08117EFE",
    x"08114634",
    x"08110D7F",
    x"0810D4E1",
    x"08109C59",
    x"081063E7",
    x"08102B8B",
    x"080FF345",
    x"080FBB15",
    x"080F82FB",
    x"080F4AF6",
    x"080F1308",
    x"080EDB30",
    x"080EA36D",
    x"080E6BC0",
    x"080E3429",
    x"080DFCA7",
    x"080DC53B",
    x"080D8DE5",
    x"080D56A4",
    x"080D1F79",
    x"080CE864",
    x"080CB164",
    x"080C7A79",
    x"080C43A4",
    x"080C0CE4",
    x"080BD63A",
    x"080B9FA5",
    x"080B6925",
    x"080B32BB",
    x"080AFC66",
    x"080AC626",
    x"080A8FFB",
    x"080A59E5",
    x"080A23E5",
    x"0809EDF9",
    x"0809B823",
    x"08098261",
    x"08094CB5",
    x"0809171D",
    x"0808E19B",
    x"0808AC2D",
    x"080876D4",
    x"08084190",
    x"08080C61",
    x"0807D747",
    x"0807A241",
    x"08076D50",
    x"08073873",
    x"080703AC",
    x"0806CEF8",
    x"08069A5A",
    x"080665D0",
    x"0806315A",
    x"0805FCF9",
    x"0805C8AD",
    x"08059475",
    x"08056051",
    x"08052C41",
    x"0804F846",
    x"0804C45F",
    x"0804908D",
    x"08045CCE",
    x"08042924",
    x"0803F58E",
    x"0803C20C",
    x"08038E9F",
    x"08035B45",
    x"080327FF",
    x"0802F4CE",
    x"0802C1B0",
    x"08028EA6",
    x"08025BB1",
    x"080228CF",
    x"0801F601",
    x"0801C347",
    x"080190A0",
    x"08015E0E",
    x"08012B8F",
    x"0800F923",
    x"0800C6CC",
    x"08009488",
    x"08006258",
    x"0800303B",
    x"07FFFC64",
    x"07FF9879",
    x"07FF34B5",
    x"07FED118",
    x"07FE6DA2",
    x"07FE0A53",
    x"07FDA72A",
    x"07FD4428",
    x"07FCE14D",
    x"07FC7E98",
    x"07FC1C0A",
    x"07FBB9A2",
    x"07FB5761",
    x"07FAF546",
    x"07FA9351",
    x"07FA3183",
    x"07F9CFDA",
    x"07F96E58",
    x"07F90CFC",
    x"07F8ABC6",
    x"07F84AB6",
    x"07F7E9CC",
    x"07F78907",
    x"07F72869",
    x"07F6C7F0",
    x"07F6679C",
    x"07F6076F",
    x"07F5A766",
    x"07F54784",
    x"07F4E7C7",
    x"07F4882F",
    x"07F428BC",
    x"07F3C96F",
    x"07F36A47",
    x"07F30B44",
    x"07F2AC66",
    x"07F24DAD",
    x"07F1EF19",
    x"07F190AA",
    x"07F13260",
    x"07F0D43B",
    x"07F0763A",
    x"07F0185F",
    x"07EFBAA7",
    x"07EF5D15",
    x"07EEFFA7",
    x"07EEA25D",
    x"07EE4538",
    x"07EDE837",
    x"07ED8B5A",
    x"07ED2EA2",
    x"07ECD20E",
    x"07EC759E",
    x"07EC1952",
    x"07EBBD2A",
    x"07EB6126",
    x"07EB0546",
    x"07EAA98A",
    x"07EA4DF2",
    x"07E9F27D",
    x"07E9972C",
    x"07E93BFF",
    x"07E8E0F5",
    x"07E8860F",
    x"07E82B4D",
    x"07E7D0AD",
    x"07E77632",
    x"07E71BD9",
    x"07E6C1A4",
    x"07E66792",
    x"07E60DA3",
    x"07E5B3D7",
    x"07E55A2E",
    x"07E500A9",
    x"07E4A746",
    x"07E44E06",
    x"07E3F4E9",
    x"07E39BEF",
    x"07E34317",
    x"07E2EA62",
    x"07E291D0",
    x"07E23960",
    x"07E1E113",
    x"07E188E8",
    x"07E130E0",
    x"07E0D8FA",
    x"07E08136",
    x"07E02995",
    x"07DFD216",
    x"07DF7AB9",
    x"07DF237E",
    x"07DECC65",
    x"07DE756E",
    x"07DE1E99",
    x"07DDC7E6",
    x"07DD7155",
    x"07DD1AE6",
    x"07DCC498",
    x"07DC6E6C",
    x"07DC1862",
    x"07DBC279",
    x"07DB6CB2",
    x"07DB170C",
    x"07DAC188",
    x"07DA6C25",
    x"07DA16E4",
    x"07D9C1C3",
    x"07D96CC4",
    x"07D917E6",
    x"07D8C329",
    x"07D86E8E",
    x"07D81A13",
    x"07D7C5B9",
    x"07D77181",
    x"07D71D69",
    x"07D6C972",
    x"07D6759B",
    x"07D621E6",
    x"07D5CE51",
    x"07D57ADC",
    x"07D52789",
    x"07D4D456",
    x"07D48143",
    x"07D42E51",
    x"07D3DB7F",
    x"07D388CD",
    x"07D3363C",
    x"07D2E3CB",
    x"07D2917A",
    x"07D23F49",
    x"07D1ED38",
    x"07D19B48",
    x"07D14977",
    x"07D0F7C6",
    x"07D0A635",
    x"07D054C4",
    x"07D00373",
    x"07CFB242",
    x"07CF6130",
    x"07CF103E",
    x"07CEBF6B",
    x"07CE6EB8",
    x"07CE1E25",
    x"07CDCDB1",
    x"07CD7D5C",
    x"07CD2D27",
    x"07CCDD11",
    x"07CC8D1A",
    x"07CC3D42",
    x"07CBED8A",
    x"07CB9DF1",
    x"07CB4E77",
    x"07CAFF1B",
    x"07CAAFDF",
    x"07CA60C2",
    x"07CA11C4",
    x"07C9C2E4",
    x"07C97423",
    x"07C92581",
    x"07C8D6FE",
    x"07C88899",
    x"07C83A53",
    x"07C7EC2C",
    x"07C79E23",
    x"07C75038",
    x"07C7026C",
    x"07C6B4BE",
    x"07C6672F",
    x"07C619BE",
    x"07C5CC6B",
    x"07C57F36",
    x"07C5321F",
    x"07C4E527",
    x"07C4984C",
    x"07C44B90",
    x"07C3FEF1",
    x"07C3B271",
    x"07C3660E",
    x"07C319C9",
    x"07C2CDA2",
    x"07C28198",
    x"07C235AD",
    x"07C1E9DE",
    x"07C19E2E",
    x"07C1529B",
    x"07C10725",
    x"07C0BBCD",
    x"07C07092",
    x"07C02575",
    x"07BFDA75",
    x"07BF8F93",
    x"07BF44CD",
    x"07BEFA25",
    x"07BEAF9A",
    x"07BE652C",
    x"07BE1ADB",
    x"07BDD0A7",
    x"07BD8690",
    x"07BD3C95",
    x"07BCF2B8",
    x"07BCA8F8",
    x"07BC5F54",
    x"07BC15CD",
    x"07BBCC63",
    x"07BB8316",
    x"07BB39E5",
    x"07BAF0D0",
    x"07BAA7D9",
    x"07BA5EFD",
    x"07BA163E",
    x"07B9CD9C",
    x"07B98516",
    x"07B93CAC",
    x"07B8F45E",
    x"07B8AC2D",
    x"07B86418",
    x"07B81C1F",
    x"07B7D442",
    x"07B78C81",
    x"07B744DC",
    x"07B6FD53",
    x"07B6B5E6",
    x"07B66E95",
    x"07B62760",
    x"07B5E046",
    x"07B59948",
    x"07B55266",
    x"07B50BA0",
    x"07B4C4F5",
    x"07B47E66",
    x"07B437F3",
    x"07B3F19A",
    x"07B3AB5E",
    x"07B3653D",
    x"07B31F37",
    x"07B2D94C",
    x"07B2937D",
    x"07B24DC9",
    x"07B20830",
    x"07B1C2B2",
    x"07B17D50",
    x"07B13809",
    x"07B0F2DC",
    x"07B0ADCB",
    x"07B068D4",
    x"07B023F9",
    x"07AFDF38",
    x"07AF9A92",
    x"07AF5607",
    x"07AF1197",
    x"07AECD42",
    x"07AE8907",
    x"07AE44E7",
    x"07AE00E1",
    x"07ADBCF6",
    x"07AD7925",
    x"07AD356F",
    x"07ACF1D4",
    x"07ACAE52",
    x"07AC6AEB",
    x"07AC279F",
    x"07ABE46C",
    x"07ABA154",
    x"07AB5E56",
    x"07AB1B73",
    x"07AAD8A9",
    x"07AA95F9",
    x"07AA5364",
    x"07AA10E8",
    x"07A9CE87",
    x"07A98C3F",
    x"07A94A11",
    x"07A907FD",
    x"07A8C603",
    x"07A88422",
    x"07A8425B",
    x"07A800AE",
    x"07A7BF1B",
    x"07A77DA1",
    x"07A73C41",
    x"07A6FAFA",
    x"07A6B9CD",
    x"07A678B9",
    x"07A637BE",
    x"07A5F6DD",
    x"07A5B615",
    x"07A57567",
    x"07A534D2",
    x"07A4F456",
    x"07A4B3F3",
    x"07A473A9",
    x"07A43378",
    x"07A3F361",
    x"07A3B362",
    x"07A3737D",
    x"07A333B0",
    x"07A2F3FC",
    x"07A2B461",
    x"07A274DF",
    x"07A23576",
    x"07A1F626",
    x"07A1B6EE",
    x"07A177CF",
    x"07A138C8",
    x"07A0F9DA",
    x"07A0BB05",
    x"07A07C48",
    x"07A03DA4",
    x"079FFF18",
    x"079FC0A5",
    x"079F824A",
    x"079F4407",
    x"079F05DC",
    x"079EC7CA",
    x"079E89D0",
    x"079E4BEF",
    x"079E0E25",
    x"079DD073",
    x"079D92DA",
    x"079D5559",
    x"079D17EF",
    x"079CDA9E",
    x"079C9D65",
    x"079C6043",
    x"079C2339",
    x"079BE648",
    x"079BA96D",
    x"079B6CAB",
    x"079B3001",
    x"079AF36E",
    x"079AB6F2",
    x"079A7A8F",
    x"079A3E43",
    x"079A020E",
    x"0799C5F1",
    x"079989EB",
    x"07994DFD",
    x"07991226",
    x"0798D667",
    x"07989ABF",
    x"07985F2E",
    x"079823B5",
    x"0797E852",
    x"0797AD07",
    x"079771D3",
    x"079736B6",
    x"0796FBB0",
    x"0796C0C1",
    x"079685EA",
    x"07964B29",
    x"0796107F",
    x"0795D5EC",
    x"07959B70",
    x"0795610A",
    x"079526BC",
    x"0794EC84",
    x"0794B263",
    x"07947859",
    x"07943E65",
    x"07940488",
    x"0793CAC2",
    x"07939112",
    x"07935778",
    x"07931DF5",
    x"0792E489",
    x"0792AB33",
    x"079271F3",
    x"079238CA",
    x"0791FFB7",
    x"0791C6BA",
    x"07918DD3",
    x"07915503",
    x"07911C49",
    x"0790E3A5",
    x"0790AB17",
    x"0790729F",
    x"07903A3E",
    x"079001F2",
    x"078FC9BC",
    x"078F919C",
    x"078F5992",
    x"078F219E",
    x"078EE9C0",
    x"078EB1F8",
    x"078E7A45",
    x"078E42A8",
    x"078E0B21",
    x"078DD3AF",
    x"078D9C53",
    x"078D650D",
    x"078D2DDD",
    x"078CF6C1",
    x"078CBFBC",
    x"078C88CC",
    x"078C51F1",
    x"078C1B2C",
    x"078BE47C",
    x"078BADE1",
    x"078B775C",
    x"078B40EC",
    x"078B0A91",
    x"078AD44B",
    x"078A9E1B",
    x"078A6800",
    x"078A31FA",
    x"0789FC09",
    x"0789C62D",
    x"07899066",
    x"07895AB4",
    x"07892517",
    x"0788EF8F",
    x"0788BA1C",
    x"078884BE",
    x"07884F74",
    x"07881A40",
    x"0787E520",
    x"0787B015",
    x"07877B1E",
    x"0787463C",
    x"0787116F",
    x"0786DCB7",
    x"0786A813",
    x"07867384",
    x"07863F09",
    x"07860AA2",
    x"0785D650",
    x"0785A213",
    x"07856DEA",
    x"078539D5",
    x"078505D5",
    x"0784D1E8",
    x"07849E11",
    x"07846A4D",
    x"0784369D",
    x"07840302",
    x"0783CF7B",
    x"07839C08",
    x"078368A9",
    x"0783355E",
    x"07830227",
    x"0782CF05",
    x"07829BF6",
    x"078268FB",
    x"07823614",
    x"07820341",
    x"0781D081",
    x"07819DD6",
    x"07816B3E",
    x"078138BA",
    x"0781064A",
    x"0780D3ED",
    x"0780A1A4",
    x"07806F6F",
    x"07803D4D",
    x"07800B3F",
    x"077FB288",
    x"077F4EBA",
    x"077EEB13",
    x"077E8792",
    x"077E2439",
    x"077DC106",
    x"077D5DFA",
    x"077CFB14",
    x"077C9856",
    x"077C35BD",
    x"077BD34C",
    x"077B7100",
    x"077B0EDB",
    x"077AACDD",
    x"077A4B04",
    x"0779E952",
    x"077987C6",
    x"07792660",
    x"0778C520",
    x"07786406",
    x"07780312",
    x"0777A244",
    x"0777419B",
    x"0776E118",
    x"077680BB",
    x"07762084",
    x"0775C072",
    x"07756085",
    x"077500BE",
    x"0774A11D",
    x"077441A0",
    x"0773E249",
    x"07738318",
    x"0773240B",
    x"0772C523",
    x"07726661",
    x"077207C3",
    x"0771A94B",
    x"07714AF7",
    x"0770ECC8",
    x"07708EBE",
    x"077030D9",
    x"076FD318",
    x"076F757C",
    x"076F1804",
    x"076EBAB1",
    x"076E5D82",
    x"076E0078",
    x"076DA392",
    x"076D46D0",
    x"076CEA33",
    x"076C8DB9",
    x"076C3164",
    x"076BD533",
    x"076B7925",
    x"076B1D3C",
    x"076AC176",
    x"076A65D5",
    x"076A0A57",
    x"0769AEFD",
    x"076953C6",
    x"0768F8B3",
    x"07689DC4",
    x"076842F8",
    x"0767E84F",
    x"07678DCA",
    x"07673369",
    x"0766D92A",
    x"07667F0F",
    x"07662517",
    x"0765CB42",
    x"07657190",
    x"07651801",
    x"0764BE95",
    x"0764654C",
    x"07640C26",
    x"0763B323",
    x"07635A42",
    x"07630184",
    x"0762A8E9",
    x"07625070",
    x"0761F81A",
    x"07619FE7",
    x"076147D5",
    x"0760EFE6",
    x"0760981A",
    x"07604070",
    x"075FE8E7",
    x"075F9182",
    x"075F3A3E",
    x"075EE31C",
    x"075E8C1C",
    x"075E353F",
    x"075DDE83",
    x"075D87E9",
    x"075D3170",
    x"075CDB1A",
    x"075C84E5",
    x"075C2ED2",
    x"075BD8E1",
    x"075B8311",
    x"075B2D62",
    x"075AD7D5",
    x"075A826A",
    x"075A2D1F",
    x"0759D7F6",
    x"075982EF",
    x"07592E08",
    x"0758D943",
    x"0758849E",
    x"0758301B",
    x"0757DBB9",
    x"07578777",
    x"07573357",
    x"0756DF57",
    x"07568B78",
    x"075637BA",
    x"0755E41D",
    x"075590A0",
    x"07553D44",
    x"0754EA08",
    x"075496ED",
    x"075443F2",
    x"0753F118",
    x"07539E5E",
    x"07534BC4",
    x"0752F94B",
    x"0752A6F1",
    x"075254B8",
    x"0752029F",
    x"0751B0A6",
    x"07515ECD",
    x"07510D14",
    x"0750BB7B",
    x"07506A02",
    x"075018A8",
    x"074FC76E",
    x"074F7654",
    x"074F255A",
    x"074ED47F",
    x"074E83C4",
    x"074E3328",
    x"074DE2AC",
    x"074D924F",
    x"074D4212",
    x"074CF1F3",
    x"074CA1F4",
    x"074C5215",
    x"074C0254",
    x"074BB2B3",
    x"074B6331",
    x"074B13CD",
    x"074AC489",
    x"074A7564",
    x"074A265D",
    x"0749D776",
    x"074988AD",
    x"07493A03",
    x"0748EB78",
    x"07489D0B",
    x"07484EBD",
    x"0748008E",
    x"0747B27D",
    x"0747648A",
    x"074716B6",
    x"0746C900",
    x"07467B69",
    x"07462DF0",
    x"0745E095",
    x"07459359",
    x"0745463A",
    x"0744F93A",
    x"0744AC57",
    x"07445F93",
    x"074412ED",
    x"0743C664",
    x"074379FA",
    x"07432DAD",
    x"0742E17E",
    x"0742956D",
    x"07424979",
    x"0741FDA3",
    x"0741B1EB",
    x"07416650",
    x"07411AD3",
    x"0740CF73",
    x"07408431",
    x"0740390C",
    x"073FEE04",
    x"073FA31A",
    x"073F584D",
    x"073F0D9D",
    x"073EC30A",
    x"073E7895",
    x"073E2E3C",
    x"073DE400",
    x"073D99E2",
    x"073D4FE0",
    x"073D05FB",
    x"073CBC34",
    x"073C7288",
    x"073C28FA",
    x"073BDF88",
    x"073B9633",
    x"073B4CFB",
    x"073B03DF",
    x"073ABAE0",
    x"073A71FD",
    x"073A2937",
    x"0739E08D",
    x"07399800",
    x"07394F8E",
    x"07390739",
    x"0738BF01",
    x"073876E4",
    x"07382EE4",
    x"0737E6FF",
    x"07379F37",
    x"0737578B",
    x"07370FFB",
    x"0736C887",
    x"0736812E",
    x"073639F2",
    x"0735F2D1",
    x"0735ABCC",
    x"073564E3",
    x"07351E15",
    x"0734D763",
    x"073490CD",
    x"07344A52",
    x"073403F3",
    x"0733BDAF",
    x"07337787",
    x"0733317A",
    x"0732EB88",
    x"0732A5B1",
    x"07325FF6",
    x"07321A56",
    x"0731D4D2",
    x"07318F68",
    x"07314A1A",
    x"073104E6",
    x"0730BFCE",
    x"07307AD0",
    x"073035EE",
    x"072FF126",
    x"072FAC7A",
    x"072F67E8",
    x"072F2370",
    x"072EDF14",
    x"072E9AD2",
    x"072E56AB",
    x"072E129E",
    x"072DCEAC",
    x"072D8AD5",
    x"072D4718",
    x"072D0375",
    x"072CBFED",
    x"072C7C7F",
    x"072C392C",
    x"072BF5F3",
    x"072BB2D4",
    x"072B6FCF",
    x"072B2CE4",
    x"072AEA14",
    x"072AA75D",
    x"072A64C1",
    x"072A223F",
    x"0729DFD6",
    x"07299D88",
    x"07295B53",
    x"07291938",
    x"0728D738",
    x"07289550",
    x"07285383",
    x"072811CF",
    x"0727D035",
    x"07278EB4",
    x"07274D4D",
    x"07270C00",
    x"0726CACC",
    x"072689B2",
    x"072648B0",
    x"072607C9",
    x"0725C6FA",
    x"07258645",
    x"072545A9",
    x"07250527",
    x"0724C4BD",
    x"0724846D",
    x"07244436",
    x"07240418",
    x"0723C413",
    x"07238427",
    x"07234453",
    x"07230499",
    x"0722C4F8",
    x"0722856F",
    x"07224600",
    x"072206A9",
    x"0721C76A",
    x"07218845",
    x"07214938",
    x"07210A44",
    x"0720CB68",
    x"07208CA5",
    x"07204DFA",
    x"07200F68",
    x"071FD0EE",
    x"071F928D",
    x"071F5443",
    x"071F1613",
    x"071ED7FA",
    x"071E99FA",
    x"071E5C12",
    x"071E1E42",
    x"071DE08A",
    x"071DA2EB",
    x"071D6563",
    x"071D27F3",
    x"071CEA9C",
    x"071CAD5C",
    x"071C7034",
    x"071C3324",
    x"071BF62C",
    x"071BB94C",
    x"071B7C84",
    x"071B3FD3",
    x"071B033A",
    x"071AC6B8",
    x"071A8A4E",
    x"071A4DFC",
    x"071A11C1",
    x"0719D59E",
    x"07199993",
    x"07195D9E",
    x"071921C1",
    x"0718E5FC",
    x"0718AA4E",
    x"07186EB7",
    x"07183337",
    x"0717F7CF",
    x"0717BC7E",
    x"07178144",
    x"07174621",
    x"07170B15",
    x"0716D020",
    x"07169542",
    x"07165A7B",
    x"07161FCB",
    x"0715E532",
    x"0715AAB0",
    x"07157045",
    x"071535F1",
    x"0714FBB3",
    x"0714C18C",
    x"0714877C",
    x"07144D82",
    x"0714139F",
    x"0713D9D3",
    x"0713A01D",
    x"0713667E",
    x"07132CF5",
    x"0712F383",
    x"0712BA27",
    x"071280E1",
    x"071247B2",
    x"07120E99",
    x"0711D597",
    x"07119CAA",
    x"071163D4",
    x"07112B14",
    x"0710F26A",
    x"0710B9D7",
    x"07108159",
    x"071048F2",
    x"071010A0",
    x"070FD865",
    x"070FA03F",
    x"070F6830",
    x"070F3036",
    x"070EF852",
    x"070EC084",
    x"070E88CB",
    x"070E5129",
    x"070E199C",
    x"070DE225",
    x"070DAAC3",
    x"070D7377",
    x"070D3C41",
    x"070D0520",
    x"070CCE15",
    x"070C971F",
    x"070C603F",
    x"070C2974",
    x"070BF2BF",
    x"070BBC1E",
    x"070B8594",
    x"070B4F1E",
    x"070B18BE",
    x"070AE273",
    x"070AAC3D",
    x"070A761C",
    x"070A4011",
    x"070A0A1A",
    x"0709D439",
    x"07099E6C",
    x"070968B5",
    x"07093313",
    x"0708FD85",
    x"0708C80C",
    x"070892A9",
    x"07085D5A",
    x"07082820",
    x"0707F2FB",
    x"0707BDEA",
    x"070788EE",
    x"07075407",
    x"07071F34",
    x"0706EA77",
    x"0706B5CD",
    x"07068139",
    x"07064CB8",
    x"0706184D",
    x"0705E3F5",
    x"0705AFB2",
    x"07057B84",
    x"0705476A",
    x"07051364",
    x"0704DF73",
    x"0704AB96",
    x"070477CD",
    x"07044418",
    x"07041078",
    x"0703DCEB",
    x"0703A973",
    x"0703760F",
    x"070342BF",
    x"07030F83",
    x"0702DC5B",
    x"0702A946",
    x"07027646",
    x"0702435A",
    x"07021082",
    x"0701DDBD",
    x"0701AB0C",
    x"07017870",
    x"070145E6",
    x"07011371",
    x"0700E10F",
    x"0700AEC1",
    x"07007C87",
    x"07004A60",
    x"0700184C",
    x"06FFCC9A",
    x"06FF68C1",
    x"06FF0510",
    x"06FEA185",
    x"06FE3E21",
    x"06FDDAE5",
    x"06FD77CE",
    x"06FD14DF",
    x"06FCB216",
    x"06FC4F74",
    x"06FBECF8",
    x"06FB8AA3",
    x"06FB2874",
    x"06FAC66B",
    x"06FA6489",
    x"06FA02CC",
    x"06F9A136",
    x"06F93FC7",
    x"06F8DE7D",
    x"06F87D59",
    x"06F81C5B",
    x"06F7BB83",
    x"06F75AD0",
    x"06F6FA44",
    x"06F699DD",
    x"06F6399B",
    x"06F5D980",
    x"06F57989",
    x"06F519B9",
    x"06F4BA0D",
    x"06F45A87",
    x"06F3FB27",
    x"06F39BEB",
    x"06F33CD5",
    x"06F2DDE3",
    x"06F27F17",
    x"06F22070",
    x"06F1C1EE",
    x"06F16391",
    x"06F10558",
    x"06F0A744",
    x"06F04955",
    x"06EFEB8B",
    x"06EF8DE5",
    x"06EF3064",
    x"06EED308",
    x"06EE75CF",
    x"06EE18BC",
    x"06EDBBCC",
    x"06ED5F01",
    x"06ED025A",
    x"06ECA5D7",
    x"06EC4978",
    x"06EBED3E",
    x"06EB9127",
    x"06EB3534",
    x"06EAD965",
    x"06EA7DBA",
    x"06EA2233",
    x"06E9C6D0",
    x"06E96B90",
    x"06E91073",
    x"06E8B57B",
    x"06E85AA6",
    x"06E7FFF4",
    x"06E7A566",
    x"06E74AFB",
    x"06E6F0B3",
    x"06E6968F",
    x"06E63C8D",
    x"06E5E2AF",
    x"06E588F4",
    x"06E52F5C",
    x"06E4D5E7",
    x"06E47C95",
    x"06E42366",
    x"06E3CA5A",
    x"06E37170",
    x"06E318A9",
    x"06E2C005",
    x"06E26783",
    x"06E20F24",
    x"06E1B6E7",
    x"06E15ECD",
    x"06E106D5",
    x"06E0AEFF",
    x"06E0574C",
    x"06DFFFBB",
    x"06DFA84C",
    x"06DF5100",
    x"06DEF9D5",
    x"06DEA2CD",
    x"06DE4BE6",
    x"06DDF521",
    x"06DD9E7E",
    x"06DD47FD",
    x"06DCF19E",
    x"06DC9B61",
    x"06DC4545",
    x"06DBEF4A",
    x"06DB9972",
    x"06DB43BB",
    x"06DAEE25",
    x"06DA98B1",
    x"06DA435E",
    x"06D9EE2C",
    x"06D9991B",
    x"06D9442C",
    x"06D8EF5E",
    x"06D89AB1",
    x"06D84625",
    x"06D7F1BA",
    x"06D79D70",
    x"06D74947",
    x"06D6F53F",
    x"06D6A158",
    x"06D64D91",
    x"06D5F9EB",
    x"06D5A666",
    x"06D55301",
    x"06D4FFBD",
    x"06D4AC99",
    x"06D45996",
    x"06D406B3",
    x"06D3B3F1",
    x"06D3614F",
    x"06D30ECD",
    x"06D2BC6B",
    x"06D26A2A",
    x"06D21808",
    x"06D1C607",
    x"06D17425",
    x"06D12264",
    x"06D0D0C3",
    x"06D07F41",
    x"06D02DDF",
    x"06CFDC9D",
    x"06CF8B7B",
    x"06CF3A78",
    x"06CEE995",
    x"06CE98D2",
    x"06CE482E",
    x"06CDF7A9",
    x"06CDA744",
    x"06CD56FF",
    x"06CD06D8",
    x"06CCB6D1",
    x"06CC66E9",
    x"06CC1721",
    x"06CBC777",
    x"06CB77ED",
    x"06CB2882",
    x"06CAD935",
    x"06CA8A08",
    x"06CA3AF9",
    x"06C9EC0A",
    x"06C99D39",
    x"06C94E87",
    x"06C8FFF4",
    x"06C8B17F",
    x"06C86329",
    x"06C814F1",
    x"06C7C6D9",
    x"06C778DE",
    x"06C72B02",
    x"06C6DD44",
    x"06C68FA5",
    x"06C64224",
    x"06C5F4C2",
    x"06C5A77D",
    x"06C55A57",
    x"06C50D4E",
    x"06C4C064",
    x"06C47398",
    x"06C426EA",
    x"06C3DA5A",
    x"06C38DE7",
    x"06C34193",
    x"06C2F55C",
    x"06C2A943",
    x"06C25D48",
    x"06C2116A",
    x"06C1C5AA",
    x"06C17A08",
    x"06C12E83",
    x"06C0E31B",
    x"06C097D1",
    x"06C04CA5",
    x"06C00196",
    x"06BFB6A4",
    x"06BF6BCF",
    x"06BF2117",
    x"06BED67D",
    x"06BE8C00",
    x"06BE41A0",
    x"06BDF75C",
    x"06BDAD36",
    x"06BD632D",
    x"06BD1941",
    x"06BCCF71",
    x"06BC85BF",
    x"06BC3C29",
    x"06BBF2B0",
    x"06BBA953",
    x"06BB6013",
    x"06BB16F0",
    x"06BACDE9",
    x"06BA84FF",
    x"06BA3C32",
    x"06B9F380",
    x"06B9AAEB",
    x"06B96273",
    x"06B91A16",
    x"06B8D1D6",
    x"06B889B2",
    x"06B841AB",
    x"06B7F9BF",
    x"06B7B1F0",
    x"06B76A3C",
    x"06B722A5",
    x"06B6DB29",
    x"06B693C9",
    x"06B64C86",
    x"06B6055E",
    x"06B5BE51",
    x"06B57761",
    x"06B5308C",
    x"06B4E9D3",
    x"06B4A335",
    x"06B45CB3",
    x"06B4164D",
    x"06B3D002",
    x"06B389D2",
    x"06B343BE",
    x"06B2FDC5",
    x"06B2B7E8",
    x"06B27226",
    x"06B22C7F",
    x"06B1E6F3",
    x"06B1A182",
    x"06B15C2D",
    x"06B116F2",
    x"06B0D1D3",
    x"06B08CCE",
    x"06B047E5",
    x"06B00316",
    x"06AFBE62",
    x"06AF79C9",
    x"06AF354B",
    x"06AEF0E8",
    x"06AEAC9F",
    x"06AE6871",
    x"06AE245D",
    x"06ADE064",
    x"06AD9C86",
    x"06AD58C2",
    x"06AD1519",
    x"06ACD18A",
    x"06AC8E15",
    x"06AC4ABB",
    x"06AC077B",
    x"06ABC455",
    x"06AB8149",
    x"06AB3E58",
    x"06AAFB81",
    x"06AAB8C3",
    x"06AA7620",
    x"06AA3397",
    x"06A9F128",
    x"06A9AED3",
    x"06A96C97",
    x"06A92A76",
    x"06A8E86E",
    x"06A8A680",
    x"06A864AC",
    x"06A822F1",
    x"06A7E151",
    x"06A79FC9",
    x"06A75E5C",
    x"06A71D08",
    x"06A6DBCD",
    x"06A69AAC",
    x"06A659A4",
    x"06A618B6",
    x"06A5D7E1",
    x"06A59725",
    x"06A55683",
    x"06A515FA",
    x"06A4D58A",
    x"06A49533",
    x"06A454F5",
    x"06A414D0",
    x"06A3D4C5",
    x"06A394D2",
    x"06A354F9",
    x"06A31538",
    x"06A2D590",
    x"06A29601",
    x"06A2568B",
    x"06A2172D",
    x"06A1D7E9",
    x"06A198BD",
    x"06A159A9",
    x"06A11AAF",
    x"06A0DBCC",
    x"06A09D03",
    x"06A05E52",
    x"06A01FB9",
    x"069FE139",
    x"069FA2D1",
    x"069F6482",
    x"069F264B",
    x"069EE82C",
    x"069EAA25",
    x"069E6C37",
    x"069E2E61",
    x"069DF0A3",
    x"069DB2FD",
    x"069D756F",
    x"069D37F9",
    x"069CFA9B",
    x"069CBD55",
    x"069C8027",
    x"069C4311",
    x"069C0613",
    x"069BC92C",
    x"069B8C5E",
    x"069B4FA7",
    x"069B1307",
    x"069AD680",
    x"069A9A10",
    x"069A5DB7",
    x"069A2176",
    x"0699E54D",
    x"0699A93B",
    x"06996D41",
    x"0699315E",
    x"0698F592",
    x"0698B9DE",
    x"06987E41",
    x"069842BB",
    x"0698074D",
    x"0697CBF6",
    x"069790B6",
    x"0697558D",
    x"06971A7B",
    x"0696DF80",
    x"0696A49C",
    x"069669CF",
    x"06962F19",
    x"0695F47B",
    x"0695B9F2",
    x"06957F81",
    x"06954527",
    x"06950AE3",
    x"0694D0B6",
    x"069496A0",
    x"06945CA1",
    x"069422B8",
    x"0693E8E6",
    x"0693AF2A",
    x"06937585",
    x"06933BF6",
    x"0693027E",
    x"0692C91C",
    x"06928FD1",
    x"0692569C",
    x"06921D7D",
    x"0691E475",
    x"0691AB83",
    x"069172A7",
    x"069139E1",
    x"06910131",
    x"0690C898",
    x"06909015",
    x"069057A7",
    x"06901F50",
    x"068FE70F",
    x"068FAEE4",
    x"068F76CE",
    x"068F3ECF",
    x"068F06E5",
    x"068ECF11",
    x"068E9753",
    x"068E5FAB",
    x"068E2819",
    x"068DF09C",
    x"068DB935",
    x"068D81E3",
    x"068D4AA7",
    x"068D1381",
    x"068CDC70",
    x"068CA575",
    x"068C6E8F",
    x"068C37BE",
    x"068C0103",
    x"068BCA5D",
    x"068B93CD",
    x"068B5D52",
    x"068B26EC",
    x"068AF09C",
    x"068ABA60",
    x"068A843A",
    x"068A4E29",
    x"068A182D",
    x"0689E246",
    x"0689AC74",
    x"068976B7",
    x"0689410F",
    x"06890B7C",
    x"0688D5FE",
    x"0688A095",
    x"06886B41",
    x"06883601",
    x"068800D7",
    x"0687CBC1",
    x"068796BF",
    x"068761D3",
    x"06872CFB",
    x"0686F838",
    x"0686C389",
    x"06868EEF",
    x"06865A69",
    x"068625F8",
    x"0685F19C",
    x"0685BD54",
    x"06858920",
    x"06855500",
    x"068520F5",
    x"0684ECFF",
    x"0684B91C",
    x"0684854E",
    x"06845194",
    x"06841DEE",
    x"0683EA5D",
    x"0683B6DF",
    x"06838376",
    x"06835020",
    x"06831CDF",
    x"0682E9B2",
    x"0682B699",
    x"06828393",
    x"068250A2",
    x"06821DC4",
    x"0681EAFB",
    x"0681B845",
    x"068185A3",
    x"06815314",
    x"0681209A",
    x"0680EE33",
    x"0680BBE0",
    x"068089A0",
    x"06805774",
    x"0680255C",
    x"067FE6AE",
    x"067F82CB",
    x"067F1F0F",
    x"067EBB7B",
    x"067E580D",
    x"067DF4C6",
    x"067D91A6",
    x"067D2EAC",
    x"067CCBD9",
    x"067C692D",
    x"067C06A7",
    x"067BA448",
    x"067B420F",
    x"067ADFFC",
    x"067A7E10",
    x"067A1C49",
    x"0679BAAA",
    x"06795930",
    x"0678F7DC",
    x"067896AE",
    x"067835A6",
    x"0677D4C4",
    x"06777408",
    x"06771371",
    x"0676B301",
    x"067652B6",
    x"0675F290",
    x"06759290",
    x"067532B5",
    x"0674D300",
    x"06747371",
    x"06741406",
    x"0673B4C1",
    x"067355A1",
    x"0672F6A6",
    x"067297D0",
    x"0672391F",
    x"0671DA94",
    x"06717C2D",
    x"06711DEB",
    x"0670BFCD",
    x"067061D5",
    x"06700401",
    x"066FA652",
    x"066F48C7",
    x"066EEB61",
    x"066E8E1F",
    x"066E3102",
    x"066DD409",
    x"066D7734",
    x"066D1A83",
    x"066CBDF7",
    x"066C618F",
    x"066C054B",
    x"066BA92B",
    x"066B4D2F",
    x"066AF157",
    x"066A95A2",
    x"066A3A12",
    x"0669DEA5",
    x"0669835C",
    x"06692836",
    x"0668CD34",
    x"06687256",
    x"0668179B",
    x"0667BD03",
    x"0667628F",
    x"0667083E",
    x"0666AE11",
    x"06665406",
    x"0665FA1F",
    x"0665A05B",
    x"066546BA",
    x"0664ED3C",
    x"066493E0",
    x"06643AA8",
    x"0663E193",
    x"066388A0",
    x"06632FD0",
    x"0662D723",
    x"06627E98",
    x"06622630",
    x"0661CDEA",
    x"066175C7",
    x"06611DC6",
    x"0660C5E7",
    x"06606E2B",
    x"06601691",
    x"065FBF1A",
    x"065F67C4",
    x"065F1091",
    x"065EB97F",
    x"065E6290",
    x"065E0BC2",
    x"065DB516",
    x"065D5E8D",
    x"065D0825",
    x"065CB1DE",
    x"065C5BBA",
    x"065C05B7",
    x"065BAFD5",
    x"065B5A15",
    x"065B0477",
    x"065AAEFA",
    x"065A599E",
    x"065A0464",
    x"0659AF4A",
    x"06595A53",
    x"0659057C",
    x"0658B0C6",
    x"06585C32",
    x"065807BE",
    x"0657B36C",
    x"06575F3A",
    x"06570B29",
    x"0656B739",
    x"0656636A",
    x"06560FBC",
    x"0655BC2E",
    x"065568C1",
    x"06551574",
    x"0654C248",
    x"06546F3C",
    x"06541C51",
    x"0653C986",
    x"065376DB",
    x"06532451",
    x"0652D1E7",
    x"06527F9D",
    x"06522D73",
    x"0651DB6A",
    x"06518980",
    x"065137B6",
    x"0650E60C",
    x"06509482",
    x"06504318",
    x"064FF1CE",
    x"064FA0A3",
    x"064F4F99",
    x"064EFEAD",
    x"064EADE2",
    x"064E5D35",
    x"064E0CA9",
    x"064DBC3B",
    x"064D6BEE",
    x"064D1BBF",
    x"064CCBB0",
    x"064C7BC0",
    x"064C2BEF",
    x"064BDC3E",
    x"064B8CAB",
    x"064B3D38",
    x"064AEDE3",
    x"064A9EAE",
    x"064A4F97",
    x"064A00A0",
    x"0649B1C7",
    x"0649630D",
    x"06491471",
    x"0648C5F5",
    x"06487797",
    x"06482957",
    x"0647DB36",
    x"06478D34",
    x"06473F50",
    x"0646F18B",
    x"0646A3E3",
    x"0646565B",
    x"064608F0",
    x"0645BBA4",
    x"06456E75",
    x"06452165",
    x"0644D473",
    x"0644879F",
    x"06443AE9",
    x"0643EE51",
    x"0643A1D7",
    x"0643557B",
    x"0643093C",
    x"0642BD1C",
    x"06427118",
    x"06422533",
    x"0641D96B",
    x"06418DC1",
    x"06414235",
    x"0640F6C6",
    x"0640AB74",
    x"06406040",
    x"06401529",
    x"063FCA2F",
    x"063F7F53",
    x"063F3494",
    x"063EE9F2",
    x"063E9F6D",
    x"063E5505",
    x"063E0ABA",
    x"063DC08D",
    x"063D767C",
    x"063D2C88",
    x"063CE2B1",
    x"063C98F7",
    x"063C4F5A",
    x"063C05D9",
    x"063BBC75",
    x"063B732E",
    x"063B2A03",
    x"063AE0F5",
    x"063A9803",
    x"063A4F2E",
    x"063A0675",
    x"0639BDD9",
    x"06397559",
    x"06392CF5",
    x"0638E4AE",
    x"06389C83",
    x"06385474",
    x"06380C81",
    x"0637C4AA",
    x"06377CEF",
    x"06373550",
    x"0636EDCD",
    x"0636A666",
    x"06365F1B",
    x"063617EC",
    x"0635D0D9",
    x"063589E1",
    x"06354305",
    x"0634FC45",
    x"0634B5A0",
    x"06346F17",
    x"063428A9",
    x"0633E257",
    x"06339C20",
    x"06335605",
    x"06331005",
    x"0632CA20",
    x"06328457",
    x"06323EA9",
    x"0631F916",
    x"0631B39E",
    x"06316E42",
    x"06312900",
    x"0630E3DA",
    x"06309ECE",
    x"063059DE",
    x"06301508",
    x"062FD04D",
    x"062F8BAD",
    x"062F4728",
    x"062F02BE",
    x"062EBE6E",
    x"062E7A39",
    x"062E361E",
    x"062DF21E",
    x"062DAE39",
    x"062D6A6E",
    x"062D26BE",
    x"062CE328",
    x"062C9FAD",
    x"062C5C4B",
    x"062C1904",
    x"062BD5D8",
    x"062B92C5",
    x"062B4FCD",
    x"062B0CEF",
    x"062ACA2B",
    x"062A8781",
    x"062A44F1",
    x"062A027B",
    x"0629C01F",
    x"06297DDD",
    x"06293BB5",
    x"0628F9A6",
    x"0628B7B2",
    x"062875D7",
    x"06283416",
    x"0627F26E",
    x"0627B0E0",
    x"06276F6C",
    x"06272E11",
    x"0626ECD0",
    x"0626ABA8",
    x"06266A9A",
    x"062629A5",
    x"0625E8C9",
    x"0625A807",
    x"0625675E",
    x"062526CE",
    x"0624E658",
    x"0624A5FA",
    x"062465B6",
    x"0624258B",
    x"0623E579",
    x"0623A57F",
    x"0623659F",
    x"062325D8",
    x"0622E62A",
    x"0622A694",
    x"06226718",
    x"062227B4",
    x"0621E869",
    x"0621A936",
    x"06216A1C",
    x"06212B1B",
    x"0620EC33",
    x"0620AD63",
    x"06206EAB",
    x"0620300C",
    x"061FF186",
    x"061FB317",
    x"061F74C2",
    x"061F3684",
    x"061EF85F",
    x"061EBA52",
    x"061E7C5E",
    x"061E3E81",
    x"061E00BD",
    x"061DC310",
    x"061D857C",
    x"061D4800",
    x"061D0A9C",
    x"061CCD50",
    x"061C901C",
    x"061C52FF",
    x"061C15FB",
    x"061BD90E",
    x"061B9C39",
    x"061B5F7C",
    x"061B22D7",
    x"061AE649",
    x"061AA9D3",
    x"061A6D74",
    x"061A312D",
    x"0619F4FE",
    x"0619B8E6",
    x"06197CE5",
    x"061940FC",
    x"0619052A",
    x"0618C970",
    x"06188DCD",
    x"06185241",
    x"061816CD",
    x"0617DB6F",
    x"0617A029",
    x"061764FA",
    x"061729E2",
    x"0616EEE2",
    x"0616B3F8",
    x"06167925",
    x"06163E69",
    x"061603C4",
    x"0615C936",
    x"06158EBF",
    x"0615545F",
    x"06151A15",
    x"0614DFE2",
    x"0614A5C6",
    x"06146BC1",
    x"061431D2",
    x"0613F7FA",
    x"0613BE38",
    x"0613848D",
    x"06134AF9",
    x"0613117B",
    x"0612D813",
    x"06129EC2",
    x"06126587",
    x"06122C62",
    x"0611F354",
    x"0611BA5C",
    x"0611817B",
    x"061148AF",
    x"06110FFA",
    x"0610D75B",
    x"06109ED2",
    x"0610665F",
    x"06102E02",
    x"060FF5BB",
    x"060FBD8A",
    x"060F856F",
    x"060F4D69",
    x"060F157A",
    x"060EDDA1",
    x"060EA5DD",
    x"060E6E2F",
    x"060E3697",
    x"060DFF14",
    x"060DC7A8",
    x"060D9050",
    x"060D590F",
    x"060D21E3",
    x"060CEACC",
    x"060CB3CB",
    x"060C7CE0",
    x"060C460A",
    x"060C0F49",
    x"060BD89E",
    x"060BA208",
    x"060B6B87",
    x"060B351C",
    x"060AFEC6",
    x"060AC885",
    x"060A9259",
    x"060A5C42",
    x"060A2641",
    x"0609F055",
    x"0609BA7D",
    x"060984BB",
    x"06094F0D",
    x"06091975",
    x"0608E3F2",
    x"0608AE83",
    x"06087929",
    x"060843E4",
    x"06080EB4",
    x"0607D999",
    x"0607A492",
    x"06076FA0",
    x"06073AC3",
    x"060705FA",
    x"0606D146",
    x"06069CA7",
    x"0606681C",
    x"060633A5",
    x"0605FF43",
    x"0605CAF6",
    x"060596BD",
    x"06056298",
    x"06052E88",
    x"0604FA8C",
    x"0604C6A4",
    x"060492D1",
    x"06045F11",
    x"06042B66",
    x"0603F7CF",
    x"0603C44D",
    x"060390DE",
    x"06035D84",
    x"06032A3D",
    x"0602F70B",
    x"0602C3EC",
    x"060290E1",
    x"06025DEB",
    x"06022B08",
    x"0601F839",
    x"0601C57E",
    x"060192D7",
    x"06016043",
    x"06012DC4",
    x"0600FB58",
    x"0600C8FF",
    x"060096BB",
    x"0600648A",
    x"0600326C",
    x"06000062",
    x"05FF9CD8",
    x"05FF3912",
    x"05FED573",
    x"05FE71FB",
    x"05FE0EAA",
    x"05FDAB80",
    x"05FD487C",
    x"05FCE59F",
    x"05FC82E8",
    x"05FC2059",
    x"05FBBDEF",
    x"05FB5BAC",
    x"05FAF990",
    x"05FA9799",
    x"05FA35C9",
    x"05F9D41F",
    x"05F9729B",
    x"05F9113E",
    x"05F8B006",
    x"05F84EF4",
    x"05F7EE08",
    x"05F78D42",
    x"05F72CA2",
    x"05F6CC27",
    x"05F66BD2",
    x"05F60BA3",
    x"05F5AB99",
    x"05F54BB5",
    x"05F4EBF6",
    x"05F48C5C",
    x"05F42CE8",
    x"05F3CD99",
    x"05F36E70",
    x"05F30F6B",
    x"05F2B08C",
    x"05F251D1",
    x"05F1F33C",
    x"05F194CB",
    x"05F1367F",
    x"05F0D859",
    x"05F07A56",
    x"05F01C79",
    x"05EFBEC0",
    x"05EF612C",
    x"05EF03BC",
    x"05EEA671",
    x"05EE494A",
    x"05EDEC48",
    x"05ED8F69",
    x"05ED32B0",
    x"05ECD61A",
    x"05EC79A8",
    x"05EC1D5B",
    x"05EBC131",
    x"05EB652C",
    x"05EB094A",
    x"05EAAD8D",
    x"05EA51F3",
    x"05E9F67D",
    x"05E99B2A",
    x"05E93FFB",
    x"05E8E4F0",
    x"05E88A08",
    x"05E82F44",
    x"05E7D4A3",
    x"05E77A26",
    x"05E71FCC",
    x"05E6C595",
    x"05E66B82",
    x"05E61191",
    x"05E5B7C4",
    x"05E55E1A",
    x"05E50492",
    x"05E4AB2E",
    x"05E451ED",
    x"05E3F8CE",
    x"05E39FD2",
    x"05E346F9",
    x"05E2EE43",
    x"05E295AF",
    x"05E23D3E",
    x"05E1E4EF",
    x"05E18CC3",
    x"05E134B9",
    x"05E0DCD2",
    x"05E0850D",
    x"05E02D6A",
    x"05DFD5E9",
    x"05DF7E8B",
    x"05DF274E",
    x"05DED034",
    x"05DE793C",
    x"05DE2265",
    x"05DDCBB1",
    x"05DD751E",
    x"05DD1EAD",
    x"05DCC85E",
    x"05DC7231",
    x"05DC1C25",
    x"05DBC63B",
    x"05DB7072",
    x"05DB1ACB",
    x"05DAC545",
    x"05DA6FE1",
    x"05DA1A9E",
    x"05D9C57C",
    x"05D9707B",
    x"05D91B9C",
    x"05D8C6DE",
    x"05D87241",
    x"05D81DC4",
    x"05D7C969",
    x"05D7752F",
    x"05D72116",
    x"05D6CD1D",
    x"05D67945",
    x"05D6258E",
    x"05D5D1F8",
    x"05D57E82",
    x"05D52B2D",
    x"05D4D7F9",
    x"05D484E4",
    x"05D431F1",
    x"05D3DF1D",
    x"05D38C6A",
    x"05D339D8",
    x"05D2E765",
    x"05D29513",
    x"05D242E1",
    x"05D1F0CF",
    x"05D19EDD",
    x"05D14D0B",
    x"05D0FB58",
    x"05D0A9C6",
    x"05D05854",
    x"05D00701",
    x"05CFB5CE",
    x"05CF64BB",
    x"05CF13C8",
    x"05CEC2F4",
    x"05CE723F",
    x"05CE21AA",
    x"05CDD135",
    x"05CD80DF",
    x"05CD30A8",
    x"05CCE091",
    x"05CC9099",
    x"05CC40C0",
    x"05CBF106",
    x"05CBA16C",
    x"05CB51F0",
    x"05CB0294",
    x"05CAB356",
    x"05CA6437",
    x"05CA1538",
    x"05C9C657",
    x"05C97795",
    x"05C928F1",
    x"05C8DA6D",
    x"05C88C07",
    x"05C83DBF",
    x"05C7EF96",
    x"05C7A18C",
    x"05C753A0",
    x"05C705D3",
    x"05C6B824",
    x"05C66A93",
    x"05C61D20",
    x"05C5CFCC",
    x"05C58296",
    x"05C5357E",
    x"05C4E884",
    x"05C49BA8",
    x"05C44EEB",
    x"05C4024B",
    x"05C3B5C9",
    x"05C36965",
    x"05C31D1E",
    x"05C2D0F6",
    x"05C284EB",
    x"05C238FE",
    x"05C1ED2F",
    x"05C1A17D",
    x"05C155E8",
    x"05C10A72",
    x"05C0BF18",
    x"05C073DC",
    x"05C028BE",
    x"05BFDDBD",
    x"05BF92D9",
    x"05BF4812",
    x"05BEFD68",
    x"05BEB2DC",
    x"05BE686C",
    x"05BE1E1A",
    x"05BDD3E5",
    x"05BD89CD",
    x"05BD3FD1",
    x"05BCF5F3",
    x"05BCAC31",
    x"05BC628C",
    x"05BC1904",
    x"05BBCF99",
    x"05BB864A",
    x"05BB3D18",
    x"05BAF402",
    x"05BAAB09",
    x"05BA622D",
    x"05BA196C",
    x"05B9D0C9",
    x"05B98841",
    x"05B93FD6",
    x"05B8F787",
    x"05B8AF55",
    x"05B8673E",
    x"05B81F44",
    x"05B7D766",
    x"05B78FA4",
    x"05B747FE",
    x"05B70074",
    x"05B6B905",
    x"05B671B3",
    x"05B62A7C",
    x"05B5E362",
    x"05B59C63",
    x"05B55580",
    x"05B50EB8",
    x"05B4C80C",
    x"05B4817C",
    x"05B43B07",
    x"05B3F4AE",
    x"05B3AE70",
    x"05B3684D",
    x"05B32246",
    x"05B2DC5B",
    x"05B2968A",
    x"05B250D5",
    x"05B20B3B",
    x"05B1C5BC",
    x"05B18058",
    x"05B13B10",
    x"05B0F5E2",
    x"05B0B0D0",
    x"05B06BD8",
    x"05B026FB",
    x"05AFE23A",
    x"05AF9D93",
    x"05AF5907",
    x"05AF1495",
    x"05AED03E",
    x"05AE8C02",
    x"05AE47E1",
    x"05AE03DA",
    x"05ADBFEE",
    x"05AD7C1C",
    x"05AD3865",
    x"05ACF4C8",
    x"05ACB146",
    x"05AC6DDE",
    x"05AC2A90",
    x"05ABE75C",
    x"05ABA443",
    x"05AB6144",
    x"05AB1E5F",
    x"05AADB94",
    x"05AA98E4",
    x"05AA564D",
    x"05AA13D0",
    x"05A9D16D",
    x"05A98F25",
    x"05A94CF6",
    x"05A90AE0",
    x"05A8C8E5",
    x"05A88703",
    x"05A8453C",
    x"05A8038D",
    x"05A7C1F9",
    x"05A7807E",
    x"05A73F1C",
    x"05A6FDD4",
    x"05A6BCA6",
    x"05A67B91",
    x"05A63A96",
    x"05A5F9B3",
    x"05A5B8EA",
    x"05A5783B",
    x"05A537A4",
    x"05A4F727",
    x"05A4B6C3",
    x"05A47679",
    x"05A43647",
    x"05A3F62E",
    x"05A3B62E",
    x"05A37648",
    x"05A3367A",
    x"05A2F6C5",
    x"05A2B729",
    x"05A277A6",
    x"05A2383C",
    x"05A1F8EA",
    x"05A1B9B1",
    x"05A17A91",
    x"05A13B8A",
    x"05A0FC9B",
    x"05A0BDC4",
    x"05A07F06",
    x"05A04061",
    x"05A001D4",
    x"059FC35F",
    x"059F8503",
    x"059F46C0",
    x"059F0894",
    x"059ECA81",
    x"059E8C86",
    x"059E4EA3",
    x"059E10D8",
    x"059DD326",
    x"059D958B",
    x"059D5809",
    x"059D1A9F",
    x"059CDD4C",
    x"059CA012",
    x"059C62EF",
    x"059C25E4",
    x"059BE8F2",
    x"059BAC16",
    x"059B6F53",
    x"059B32A7",
    x"059AF613",
    x"059AB997",
    x"059A7D32",
    x"059A40E5",
    x"059A04B0",
    x"0599C892",
    x"05998C8B",
    x"0599509C",
    x"059914C4",
    x"0598D904",
    x"05989D5B",
    x"059861C9",
    x"0598264E",
    x"0597EAEB",
    x"0597AF9F",
    x"0597746A",
    x"0597394C",
    x"0596FE45",
    x"0596C355",
    x"0596887C",
    x"05964DBA",
    x"0596130F",
    x"0595D87B",
    x"05959DFE",
    x"05956398",
    x"05952948",
    x"0594EF10",
    x"0594B4EE",
    x"05947AE2",
    x"059440EE",
    x"05940710",
    x"0593CD48",
    x"05939397",
    x"059359FD",
    x"05932079",
    x"0592E70B",
    x"0592ADB4",
    x"05927474",
    x"05923B49",
    x"05920235",
    x"0591C938",
    x"05919050",
    x"0591577F",
    x"05911EC4",
    x"0590E61F",
    x"0590AD90",
    x"05907517",
    x"05903CB5",
    x"05900468",
    x"058FCC31",
    x"058F9410",
    x"058F5C05",
    x"058F2410",
    x"058EEC31",
    x"058EB468",
    x"058E7CB4",
    x"058E4516",
    x"058E0D8E",
    x"058DD61C",
    x"058D9EBF",
    x"058D6778",
    x"058D3046",
    x"058CF92A",
    x"058CC223",
    x"058C8B32",
    x"058C5457",
    x"058C1D90",
    x"058BE6E0",
    x"058BB044",
    x"058B79BE",
    x"058B434D",
    x"058B0CF1",
    x"058AD6AB",
    x"058AA07A",
    x"058A6A5D",
    x"058A3456",
    x"0589FE65",
    x"0589C888",
    x"058992C0",
    x"05895D0D",
    x"0589276F",
    x"0588F1E6",
    x"0588BC72",
    x"05888713",
    x"058851C9",
    x"05881C93",
    x"0587E772",
    x"0587B266",
    x"05877D6F",
    x"0587488C",
    x"058713BE",
    x"0586DF05",
    x"0586AA60",
    x"058675D0",
    x"05864154",
    x"05860CED",
    x"0585D89A",
    x"0585A45B",
    x"05857031",
    x"05853C1C",
    x"0585081A",
    x"0584D42D",
    x"0584A055",
    x"05846C90",
    x"058438E0",
    x"05840544",
    x"0583D1BC",
    x"05839E48",
    x"05836AE8",
    x"0583379C",
    x"05830465",
    x"0582D141",
    x"05829E31",
    x"05826B35",
    x"0582384D",
    x"05820579",
    x"0581D2B9",
    x"0581A00D",
    x"05816D74",
    x"05813AEF",
    x"0581087E",
    x"0580D620",
    x"0580A3D7",
    x"058071A0",
    x"05803F7E",
    x"05800D6F",
    x"057FB6E7",
    x"057F5317",
    x"057EEF6E",
    x"057E8BEC",
    x"057E2890",
    x"057DC55C",
    x"057D624E",
    x"057CFF67",
    x"057C9CA7",
    x"057C3A0D",
    x"057BD799",
    x"057B754C",
    x"057B1326",
    x"057AB125",
    x"057A4F4B",
    x"0579ED97",
    x"05798C0A",
    x"05792AA2",
    x"0578C960",
    x"05786845",
    x"0578074F",
    x"0577A67F",
    x"057745D5",
    x"0576E550",
    x"057684F2",
    x"057624B8",
    x"0575C4A5",
    x"057564B7",
    x"057504EE",
    x"0574A54B",
    x"057445CD",
    x"0573E674",
    x"05738741",
    x"05732833",
    x"0572C94A",
    x"05726A85",
    x"05720BE6",
    x"0571AD6C",
    x"05714F17",
    x"0570F0E6",
    x"057092DB",
    x"057034F4",
    x"056FD731",
    x"056F7993",
    x"056F1C1A",
    x"056EBEC5",
    x"056E6195",
    x"056E0489",
    x"056DA7A2",
    x"056D4ADE",
    x"056CEE3F",
    x"056C91C4",
    x"056C356D",
    x"056BD93A",
    x"056B7D2B",
    x"056B2140",
    x"056AC579",
    x"056A69D6",
    x"056A0E57",
    x"0569B2FB",
    x"056957C3",
    x"0568FCAE",
    x"0568A1BD",
    x"056846F0",
    x"0567EC46",
    x"056791BF",
    x"0567375C",
    x"0566DD1C",
    x"056682FF",
    x"05662906",
    x"0565CF2F",
    x"0565757C",
    x"05651BEB",
    x"0564C27E",
    x"05646934",
    x"0564100C",
    x"0563B707",
    x"05635E25",
    x"05630565",
    x"0562ACC9",
    x"0562544E",
    x"0561FBF7",
    x"0561A3C2",
    x"05614BAF",
    x"0560F3BE",
    x"05609BF0",
    x"05604445",
    x"055FECBB",
    x"055F9554",
    x"055F3E0E",
    x"055EE6EB",
    x"055E8FEA",
    x"055E390B",
    x"055DE24D",
    x"055D8BB2",
    x"055D3538",
    x"055CDEE0",
    x"055C88AA",
    x"055C3295",
    x"055BDCA2",
    x"055B86D1",
    x"055B3121",
    x"055ADB93",
    x"055A8626",
    x"055A30DA",
    x"0559DBAF",
    x"055986A6",
    x"055931BE",
    x"0558DCF7",
    x"05588852",
    x"055833CD",
    x"0557DF69",
    x"05578B26",
    x"05573704",
    x"0556E303",
    x"05568F23",
    x"05563B63",
    x"0555E7C5",
    x"05559446",
    x"055540E9",
    x"0554EDAC",
    x"05549A8F",
    x"05544793",
    x"0553F4B7",
    x"0553A1FC",
    x"05534F60",
    x"0552FCE6",
    x"0552AA8B",
    x"05525850",
    x"05520636",
    x"0551B43B",
    x"05516261",
    x"055110A7",
    x"0550BF0C",
    x"05506D91",
    x"05501C36",
    x"054FCAFB",
    x"054F79E0",
    x"054F28E4",
    x"054ED808",
    x"054E874B",
    x"054E36AE",
    x"054DE631",
    x"054D95D2",
    x"054D4593",
    x"054CF574",
    x"054CA574",
    x"054C5593",
    x"054C05D1",
    x"054BB62E",
    x"054B66AA",
    x"054B1746",
    x"054AC800",
    x"054A78DA",
    x"054A29D2",
    x"0549DAE9",
    x"05498C1F",
    x"05493D73",
    x"0548EEE7",
    x"0548A079",
    x"05485229",
    x"054803F9",
    x"0547B5E6",
    x"054767F2",
    x"05471A1D",
    x"0546CC66",
    x"05467ECD",
    x"05463153",
    x"0545E3F7",
    x"054596B9",
    x"05454999",
    x"0544FC97",
    x"0544AFB4",
    x"054462EE",
    x"05441646",
    x"0543C9BD",
    x"05437D51",
    x"05433103",
    x"0542E4D2",
    x"054298C0",
    x"05424CCB",
    x"054200F4",
    x"0541B53A",
    x"0541699E",
    x"05411E20",
    x"0540D2BF",
    x"0540877B",
    x"05403C55",
    x"053FF14C",
    x"053FA660",
    x"053F5B92",
    x"053F10E1",
    x"053EC64D",
    x"053E7BD6",
    x"053E317C",
    x"053DE73F",
    x"053D9D1F",
    x"053D531C",
    x"053D0936",
    x"053CBF6D",
    x"053C75C1",
    x"053C2C31",
    x"053BE2BE",
    x"053B9968",
    x"053B502E",
    x"053B0711",
    x"053ABE11",
    x"053A752D",
    x"053A2C65",
    x"0539E3BA",
    x"05399B2B",
    x"053952B9",
    x"05390A63",
    x"0538C229",
    x"05387A0B",
    x"05383209",
    x"0537EA24",
    x"0537A25B",
    x"05375AAD",
    x"0537131C",
    x"0536CBA6",
    x"0536844D",
    x"05363D0F",
    x"0535F5ED",
    x"0535AEE7",
    x"053567FC",
    x"0535212D",
    x"0534DA7A",
    x"053493E3",
    x"05344D67",
    x"05340706",
    x"0533C0C1",
    x"05337A98",
    x"05333489",
    x"0532EE97",
    x"0532A8BF",
    x"05326303",
    x"05321D62",
    x"0531D7DC",
    x"05319271",
    x"05314D21",
    x"053107ED",
    x"0530C2D3",
    x"05307DD4",
    x"053038F1",
    x"052FF428",
    x"052FAF7A",
    x"052F6AE7",
    x"052F266F",
    x"052EE211",
    x"052E9DCE",
    x"052E59A6",
    x"052E1598",
    x"052DD1A5",
    x"052D8DCC",
    x"052D4A0E",
    x"052D066A",
    x"052CC2E1",
    x"052C7F72",
    x"052C3C1D",
    x"052BF8E3",
    x"052BB5C3",
    x"052B72BD",
    x"052B2FD1",
    x"052AED00",
    x"052AAA48",
    x"052A67AA",
    x"052A2527",
    x"0529E2BD",
    x"0529A06E",
    x"05295E38",
    x"05291C1C",
    x"0528DA1A",
    x"05289832",
    x"05285663",
    x"052814AE",
    x"0527D313",
    x"05279191",
    x"05275029",
    x"05270EDB",
    x"0526CDA6",
    x"05268C8A",
    x"05264B88",
    x"05260A9F",
    x"0525C9D0",
    x"05258919",
    x"0525487C",
    x"052507F9",
    x"0524C78E",
    x"0524873D",
    x"05244705",
    x"052406E5",
    x"0523C6DF",
    x"052386F2",
    x"0523471E",
    x"05230762",
    x"0522C7C0",
    x"05228836",
    x"052248C5",
    x"0522096D",
    x"0521CA2E",
    x"05218B07",
    x"05214BF9",
    x"05210D04",
    x"0520CE27",
    x"05208F63",
    x"052050B7",
    x"05201224",
    x"051FD3A9",
    x"051F9547",
    x"051F56FC",
    x"051F18CB",
    x"051EDAB1",
    x"051E9CB0",
    x"051E5EC7",
    x"051E20F6",
    x"051DE33D",
    x"051DA59C",
    x"051D6813",
    x"051D2AA3",
    x"051CED4A",
    x"051CB009",
    x"051C72E1",
    x"051C35D0",
    x"051BF8D7",
    x"051BBBF5",
    x"051B7F2C",
    x"051B427A",
    x"051B05E0",
    x"051AC95D",
    x"051A8CF2",
    x"051A509F",
    x"051A1463",
    x"0519D83F",
    x"05199C32",
    x"0519603D",
    x"0519245F",
    x"0518E899",
    x"0518ACEA",
    x"05187152",
    x"051835D1",
    x"0517FA68",
    x"0517BF15",
    x"051783DA",
    x"051748B6",
    x"05170DA9",
    x"0516D2B4",
    x"051697D5",
    x"05165D0D",
    x"0516225C",
    x"0515E7C2",
    x"0515AD3F",
    x"051572D3",
    x"0515387D",
    x"0514FE3F",
    x"0514C417",
    x"05148A05",
    x"0514500B",
    x"05141627",
    x"0513DC5A",
    x"0513A2A3",
    x"05136903",
    x"05132F79",
    x"0512F605",
    x"0512BCA9",
    x"05128362",
    x"05124A32",
    x"05121118",
    x"0511D814",
    x"05119F27",
    x"05116650",
    x"05112D8F",
    x"0510F4E5",
    x"0510BC50",
    x"051083D1",
    x"05104B69",
    x"05101316",
    x"050FDADA",
    x"050FA2B3",
    x"050F6AA3",
    x"050F32A8",
    x"050EFAC3",
    x"050EC2F4",
    x"050E8B3B",
    x"050E5397",
    x"050E1C0A",
    x"050DE492",
    x"050DAD2F",
    x"050D75E2",
    x"050D3EAB",
    x"050D0789",
    x"050CD07D",
    x"050C9986",
    x"050C62A5",
    x"050C2BD9",
    x"050BF523",
    x"050BBE82",
    x"050B87F6",
    x"050B5180",
    x"050B1B1E",
    x"050AE4D2",
    x"050AAE9C",
    x"050A787A",
    x"050A426D",
    x"050A0C76",
    x"0509D694",
    x"0509A0C6",
    x"05096B0E",
    x"0509356B",
    x"0508FFDC",
    x"0508CA63",
    x"050894FE",
    x"05085FAE",
    x"05082A73",
    x"0507F54D",
    x"0507C03C",
    x"05078B3F",
    x"05075657",
    x"05072184",
    x"0506ECC5",
    x"0506B81B",
    x"05068385",
    x"05064F04",
    x"05061A97",
    x"0505E63F",
    x"0505B1FB",
    x"05057DCC",
    x"050549B1",
    x"050515AA",
    x"0504E1B8",
    x"0504ADDA",
    x"05047A10",
    x"0504465B",
    x"050412B9",
    x"0503DF2C",
    x"0503ABB3",
    x"0503784E",
    x"050344FD",
    x"050311C0",
    x"0502DE97",
    x"0502AB82",
    x"05027881",
    x"05024594",
    x"050212BB",
    x"0501DFF5",
    x"0501AD44",
    x"05017AA6",
    x"0501481C",
    x"050115A6",
    x"0500E343",
    x"0500B0F4",
    x"05007EB9",
    x"05004C91",
    x"05001A7D",
    x"04FFD0F9",
    x"04FF6D1E",
    x"04FF096B",
    x"04FEA5DF",
    x"04FE427A",
    x"04FDDF3B",
    x"04FD7C23",
    x"04FD1932",
    x"04FCB668",
    x"04FC53C4",
    x"04FBF146",
    x"04FB8EEF",
    x"04FB2CBE",
    x"04FACAB4",
    x"04FA68D0",
    x"04FA0712",
    x"04F9A57B",
    x"04F94409",
    x"04F8E2BD",
    x"04F88198",
    x"04F82098",
    x"04F7BFBE",
    x"04F75F0A",
    x"04F6FE7C",
    x"04F69E13",
    x"04F63DD0",
    x"04F5DDB3",
    x"04F57DBB",
    x"04F51DE9",
    x"04F4BE3C",
    x"04F45EB4",
    x"04F3FF52",
    x"04F3A015",
    x"04F340FD",
    x"04F2E20A",
    x"04F2833C",
    x"04F22493",
    x"04F1C610",
    x"04F167B1",
    x"04F10977",
    x"04F0AB61",
    x"04F04D71",
    x"04EFEFA5",
    x"04EF91FD",
    x"04EF347B",
    x"04EED71C",
    x"04EE79E3",
    x"04EE1CCD",
    x"04EDBFDC",
    x"04ED630F",
    x"04ED0667",
    x"04ECA9E2",
    x"04EC4D82",
    x"04EBF146",
    x"04EB952D",
    x"04EB3939",
    x"04EADD69",
    x"04EA81BC",
    x"04EA2633",
    x"04E9CACE",
    x"04E96F8D",
    x"04E9146F",
    x"04E8B975",
    x"04E85E9E",
    x"04E803EB",
    x"04E7A95B",
    x"04E74EEF",
    x"04E6F4A5",
    x"04E69A7F",
    x"04E6407D",
    x"04E5E69D",
    x"04E58CE0",
    x"04E53347",
    x"04E4D9D0",
    x"04E4807D",
    x"04E4274C",
    x"04E3CE3E",
    x"04E37553",
    x"04E31C8A",
    x"04E2C3E5",
    x"04E26B61",
    x"04E21301",
    x"04E1BAC2",
    x"04E162A7",
    x"04E10AAD",
    x"04E0B2D6",
    x"04E05B22",
    x"04E0038F",
    x"04DFAC1F",
    x"04DF54D1",
    x"04DEFDA5",
    x"04DEA69A",
    x"04DE4FB2",
    x"04DDF8EC",
    x"04DDA248",
    x"04DD4BC5",
    x"04DCF565",
    x"04DC9F26",
    x"04DC4908",
    x"04DBF30D",
    x"04DB9D32",
    x"04DB477A",
    x"04DAF1E3",
    x"04DA9C6D",
    x"04DA4718",
    x"04D9F1E5",
    x"04D99CD3",
    x"04D947E3",
    x"04D8F313",
    x"04D89E65",
    x"04D849D7",
    x"04D7F56B",
    x"04D7A120",
    x"04D74CF5",
    x"04D6F8EC",
    x"04D6A503",
    x"04D6513B",
    x"04D5FD93",
    x"04D5AA0C",
    x"04D556A6",
    x"04D50361",
    x"04D4B03C",
    x"04D45D37",
    x"04D40A53",
    x"04D3B78F",
    x"04D364EB",
    x"04D31268",
    x"04D2C005",
    x"04D26DC2",
    x"04D21B9F",
    x"04D1C99C",
    x"04D177BA",
    x"04D125F7",
    x"04D0D454",
    x"04D082D1",
    x"04D0316E",
    x"04CFE02A",
    x"04CF8F07",
    x"04CF3E03",
    x"04CEED1E",
    x"04CE9C59",
    x"04CE4BB4",
    x"04CDFB2E",
    x"04CDAAC8",
    x"04CD5A81",
    x"04CD0A59",
    x"04CCBA51",
    x"04CC6A68",
    x"04CC1A9E",
    x"04CBCAF3",
    x"04CB7B67",
    x"04CB2BFA",
    x"04CADCAD",
    x"04CA8D7E",
    x"04CA3E6E",
    x"04C9EF7D",
    x"04C9A0AB",
    x"04C951F8",
    x"04C90363",
    x"04C8B4ED",
    x"04C86696",
    x"04C8185D",
    x"04C7CA42",
    x"04C77C47",
    x"04C72E69",
    x"04C6E0AA",
    x"04C6930A",
    x"04C64588",
    x"04C5F823",
    x"04C5AADE",
    x"04C55DB6",
    x"04C510AC",
    x"04C4C3C1",
    x"04C476F3",
    x"04C42A44",
    x"04C3DDB2",
    x"04C3913F",
    x"04C344E9",
    x"04C2F8B1",
    x"04C2AC97",
    x"04C2609A",
    x"04C214BB",
    x"04C1C8FA",
    x"04C17D56",
    x"04C131D0",
    x"04C0E667",
    x"04C09B1C",
    x"04C04FEE",
    x"04C004DD",
    x"04BFB9EA",
    x"04BF6F14",
    x"04BF245B",
    x"04BED9C0",
    x"04BE8F41",
    x"04BE44E0",
    x"04BDFA9B",
    x"04BDB074",
    x"04BD666A",
    x"04BD1C7C",
    x"04BCD2AB",
    x"04BC88F7",
    x"04BC3F60",
    x"04BBF5E6",
    x"04BBAC88",
    x"04BB6347",
    x"04BB1A23",
    x"04BAD11B",
    x"04BA882F",
    x"04BA3F60",
    x"04B9F6AE",
    x"04B9AE18",
    x"04B9659E",
    x"04B91D40",
    x"04B8D4FF",
    x"04B88CDA",
    x"04B844D1",
    x"04B7FCE4",
    x"04B7B513",
    x"04B76D5E",
    x"04B725C6",
    x"04B6DE49",
    x"04B696E8",
    x"04B64FA3",
    x"04B6087A",
    x"04B5C16C",
    x"04B57A7B",
    x"04B533A5",
    x"04B4ECEA",
    x"04B4A64C",
    x"04B45FC8",
    x"04B41961",
    x"04B3D315",
    x"04B38CE4",
    x"04B346CE",
    x"04B300D4",
    x"04B2BAF6",
    x"04B27532",
    x"04B22F8A",
    x"04B1E9FD",
    x"04B1A48B",
    x"04B15F35",
    x"04B119F9",
    x"04B0D4D8",
    x"04B08FD3",
    x"04B04AE8",
    x"04B00618",
    x"04AFC163",
    x"04AF7CC9",
    x"04AF384A",
    x"04AEF3E5",
    x"04AEAF9B",
    x"04AE6B6C",
    x"04AE2757",
    x"04ADE35D",
    x"04AD9F7E",
    x"04AD5BB9",
    x"04AD180E",
    x"04ACD47E",
    x"04AC9108",
    x"04AC4DAC",
    x"04AC0A6B",
    x"04ABC744",
    x"04AB8438",
    x"04AB4145",
    x"04AAFE6C",
    x"04AABBAE",
    x"04AA790A",
    x"04AA3680",
    x"04A9F40F",
    x"04A9B1B9",
    x"04A96F7C",
    x"04A92D5A",
    x"04A8EB51",
    x"04A8A962",
    x"04A8678D",
    x"04A825D1",
    x"04A7E42F",
    x"04A7A2A7",
    x"04A76138",
    x"04A71FE3",
    x"04A6DEA7",
    x"04A69D85",
    x"04A65C7C",
    x"04A61B8D",
    x"04A5DAB6",
    x"04A599FA",
    x"04A55956",
    x"04A518CC",
    x"04A4D85B",
    x"04A49803",
    x"04A457C4",
    x"04A4179E",
    x"04A3D792",
    x"04A3979E",
    x"04A357C3",
    x"04A31801",
    x"04A2D858",
    x"04A298C8",
    x"04A25951",
    x"04A219F2",
    x"04A1DAAD",
    x"04A19B80",
    x"04A15C6B",
    x"04A11D6F",
    x"04A0DE8C",
    x"04A09FC1",
    x"04A0610F",
    x"04A02276",
    x"049FE3F4",
    x"049FA58C",
    x"049F673B",
    x"049F2903",
    x"049EEAE3",
    x"049EACDB",
    x"049E6EEC",
    x"049E3115",
    x"049DF356",
    x"049DB5AF",
    x"049D7820",
    x"049D3AA9",
    x"049CFD4A",
    x"049CC003",
    x"049C82D4",
    x"049C45BD",
    x"049C08BD",
    x"049BCBD6",
    x"049B8F06",
    x"049B524E",
    x"049B15AE",
    x"049AD925",
    x"049A9CB4",
    x"049A605B",
    x"049A2419",
    x"0499E7EE",
    x"0499ABDC",
    x"04996FE0",
    x"049933FC",
    x"0498F82F",
    x"0498BC7A",
    x"049880DC",
    x"04984556",
    x"049809E6",
    x"0497CE8E",
    x"0497934D",
    x"04975823",
    x"04971D10",
    x"0496E214",
    x"0496A72F",
    x"04966C61",
    x"049631AA",
    x"0495F70B",
    x"0495BC81",
    x"0495820F",
    x"049547B4",
    x"04950D6F",
    x"0494D341",
    x"0494992A",
    x"04945F2A",
    x"04942540",
    x"0493EB6D",
    x"0493B1B0",
    x"0493780A",
    x"04933E7A",
    x"04930501",
    x"0492CB9E",
    x"04929252",
    x"0492591C",
    x"04921FFC",
    x"0491E6F3",
    x"0491AE00",
    x"04917523",
    x"04913C5C",
    x"049103AC",
    x"0490CB11",
    x"0490928D",
    x"04905A1F",
    x"049021C7",
    x"048FE984",
    x"048FB158",
    x"048F7942",
    x"048F4141",
    x"048F0957",
    x"048ED182",
    x"048E99C3",
    x"048E621A",
    x"048E2A87",
    x"048DF309",
    x"048DBBA1",
    x"048D844E",
    x"048D4D11",
    x"048D15EA",
    x"048CDED8",
    x"048CA7DC",
    x"048C70F5",
    x"048C3A24",
    x"048C0368",
    x"048BCCC1",
    x"048B9630",
    x"048B5FB4",
    x"048B294D",
    x"048AF2FB",
    x"048ABCBF",
    x"048A8698",
    x"048A5086",
    x"048A1A89",
    x"0489E4A1",
    x"0489AECE",
    x"04897911",
    x"04894368",
    x"04890DD4",
    x"0488D855",
    x"0488A2EB",
    x"04886D96",
    x"04883855",
    x"0488032A",
    x"0487CE13",
    x"04879911",
    x"04876423",
    x"04872F4A",
    x"0486FA86",
    x"0486C5D7",
    x"0486913C",
    x"04865CB5",
    x"04862843",
    x"0485F3E6",
    x"0485BF9D",
    x"04858B68",
    x"04855748",
    x"0485233C",
    x"0484EF44",
    x"0484BB61",
    x"04848792",
    x"048453D7",
    x"04842030",
    x"0483EC9E",
    x"0483B91F",
    x"048385B5",
    x"0483525F",
    x"04831F1D",
    x"0482EBEF",
    x"0482B8D4",
    x"048285CE",
    x"048252DC",
    x"04821FFD",
    x"0481ED33",
    x"0481BA7C",
    x"048187D9",
    x"0481554A",
    x"048122CF",
    x"0480F067",
    x"0480BE13",
    x"04808BD2",
    x"048059A5",
    x"0480278C",
    x"047FEB0D",
    x"047F8729",
    x"047F236B",
    x"047EBFD5",
    x"047E5C66",
    x"047DF91D",
    x"047D95FB",
    x"047D3300",
    x"047CD02B",
    x"047C6D7D",
    x"047C0AF6",
    x"047BA894",
    x"047B465A",
    x"047AE445",
    x"047A8257",
    x"047A2090",
    x"0479BEEE",
    x"04795D72",
    x"0478FC1D",
    x"04789AED",
    x"047839E4",
    x"0477D900",
    x"04777842",
    x"047717AA",
    x"0476B738",
    x"047656EB",
    x"0475F6C4",
    x"047596C2",
    x"047536E6",
    x"0474D72F",
    x"0474779E",
    x"04741832",
    x"0473B8EB",
    x"047359C9",
    x"0472FACD",
    x"04729BF5",
    x"04723D43",
    x"0471DEB6",
    x"0471804D",
    x"04712209",
    x"0470C3EA",
    x"047065F0",
    x"0470081B",
    x"046FAA6A",
    x"046F4CDE",
    x"046EEF76",
    x"046E9233",
    x"046E3514",
    x"046DD819",
    x"046D7B43",
    x"046D1E91",
    x"046CC203",
    x"046C6599",
    x"046C0953",
    x"046BAD32",
    x"046B5134",
    x"046AF55A",
    x"046A99A4",
    x"046A3E12",
    x"0469E2A4",
    x"04698759",
    x"04692C32",
    x"0468D12F",
    x"0468764F",
    x"04681B92",
    x"0467C0F9",
    x"04676683",
    x"04670C31",
    x"0466B202",
    x"046657F6",
    x"0465FE0D",
    x"0465A447",
    x"04654AA5",
    x"0464F125",
    x"046497C8",
    x"04643E8F",
    x"0463E578",
    x"04638C83",
    x"046333B2",
    x"0462DB03",
    x"04628277",
    x"04622A0D",
    x"0461D1C6",
    x"046179A1",
    x"0461219F",
    x"0460C9BF",
    x"04607201",
    x"04601A66",
    x"045FC2EC",
    x"045F6B95",
    x"045F1460",
    x"045EBD4D",
    x"045E665C",
    x"045E0F8D",
    x"045DB8E0",
    x"045D6255",
    x"045D0BEB",
    x"045CB5A4",
    x"045C5F7E",
    x"045C0979",
    x"045BB396",
    x"045B5DD5",
    x"045B0835",
    x"045AB2B6",
    x"045A5D59",
    x"045A081D",
    x"0459B303",
    x"04595E09",
    x"04590931",
    x"0458B47A",
    x"04585FE4",
    x"04580B6F",
    x"0457B71B",
    x"045762E8",
    x"04570ED6",
    x"0456BAE5",
    x"04566714",
    x"04561364",
    x"0455BFD5",
    x"04556C66",
    x"04551918",
    x"0454C5EB",
    x"045472DE",
    x"04541FF1",
    x"0453CD25",
    x"04537A79",
    x"045327ED",
    x"0452D581",
    x"04528336",
    x"0452310B",
    x"0451DF00",
    x"04518D15",
    x"04513B49",
    x"0450E99E",
    x"04509813",
    x"045046A7",
    x"044FF55C",
    x"044FA430",
    x"044F5323",
    x"044F0237",
    x"044EB16A",
    x"044E60BC",
    x"044E102E",
    x"044DBFBF",
    x"044D6F70",
    x"044D1F40",
    x"044CCF30",
    x"044C7F3F",
    x"044C2F6C",
    x"044BDFB9",
    x"044B9026",
    x"044B40B1",
    x"044AF15B",
    x"044AA224",
    x"044A530C",
    x"044A0413",
    x"0449B539",
    x"0449667E",
    x"044917E1",
    x"0448C963",
    x"04487B04",
    x"04482CC3",
    x"0447DEA1",
    x"0447909D",
    x"044742B8",
    x"0446F4F1",
    x"0446A748",
    x"044659BE",
    x"04460C52",
    x"0445BF05",
    x"044571D5",
    x"044524C4",
    x"0444D7D0",
    x"04448AFB",
    x"04443E44",
    x"0443F1AA",
    x"0443A52F",
    x"044358D1",
    x"04430C91",
    x"0442C06F",
    x"0442746B",
    x"04422884",
    x"0441DCBB",
    x"04419110",
    x"04414582",
    x"0440FA12",
    x"0440AEBF",
    x"04406389",
    x"04401871",
    x"043FCD76",
    x"043F8298",
    x"043F37D8",
    x"043EED35",
    x"043EA2AF",
    x"043E5846",
    x"043E0DFA",
    x"043DC3CB",
    x"043D79B9",
    x"043D2FC4",
    x"043CE5EB",
    x"043C9C30",
    x"043C5291",
    x"043C090F",
    x"043BBFAA",
    x"043B7662",
    x"043B2D36",
    x"043AE426",
    x"043A9B33",
    x"043A525D",
    x"043A09A3",
    x"0439C106",
    x"04397884",
    x"0439301F",
    x"0438E7D7",
    x"04389FAA",
    x"0438579A",
    x"04380FA6",
    x"0437C7CE",
    x"04378012",
    x"04373872",
    x"0436F0EE",
    x"0436A985",
    x"04366239",
    x"04361B09",
    x"0435D3F4",
    x"04358CFB",
    x"0435461E",
    x"0434FF5C",
    x"0434B8B6",
    x"0434722C",
    x"04342BBD",
    x"0433E56A",
    x"04339F32",
    x"04335915",
    x"04331314",
    x"0432CD2E",
    x"04328764",
    x"043241B5",
    x"0431FC21",
    x"0431B6A8",
    x"0431714A",
    x"04312C07",
    x"0430E6DF",
    x"0430A1D3",
    x"04305CE1",
    x"0430180A",
    x"042FD34E",
    x"042F8EAD",
    x"042F4A27",
    x"042F05BB",
    x"042EC16A",
    x"042E7D34",
    x"042E3918",
    x"042DF517",
    x"042DB131",
    x"042D6D65",
    x"042D29B3",
    x"042CE61C",
    x"042CA2A0",
    x"042C5F3D",
    x"042C1BF5",
    x"042BD8C7",
    x"042B95B4",
    x"042B52BA",
    x"042B0FDB",
    x"042ACD16",
    x"042A8A6B",
    x"042A47DA",
    x"042A0563",
    x"0429C306",
    x"042980C2",
    x"04293E99",
    x"0428FC8A",
    x"0428BA94",
    x"042878B8",
    x"042836F5",
    x"0427F54D",
    x"0427B3BE",
    x"04277248",
    x"042730ED",
    x"0426EFAA",
    x"0426AE81",
    x"04266D72",
    x"04262C7C",
    x"0425EB9F",
    x"0425AADC",
    x"04256A32",
    x"042529A1",
    x"0424E929",
    x"0424A8CB",
    x"04246885",
    x"04242859",
    x"0423E846",
    x"0423A84B",
    x"0423686A",
    x"042328A2",
    x"0422E8F2",
    x"0422A95C",
    x"042269DE",
    x"04222A79",
    x"0421EB2D",
    x"0421ABF9",
    x"04216CDE",
    x"04212DDC",
    x"0420EEF3",
    x"0420B022",
    x"04207169",
    x"042032C9",
    x"041FF441",
    x"041FB5D2",
    x"041F777B",
    x"041F393D",
    x"041EFB17",
    x"041EBD09",
    x"041E7F13",
    x"041E4135",
    x"041E0370",
    x"041DC5C3",
    x"041D882D",
    x"041D4AB0",
    x"041D0D4B",
    x"041CCFFE",
    x"041C92C9",
    x"041C55AB",
    x"041C18A6",
    x"041BDBB8",
    x"041B9EE2",
    x"041B6224",
    x"041B257D",
    x"041AE8EE",
    x"041AAC77",
    x"041A7018",
    x"041A33D0",
    x"0419F79F",
    x"0419BB86",
    x"04197F85",
    x"0419439B",
    x"041907C8",
    x"0418CC0C",
    x"04189068",
    x"041854DC",
    x"04181966",
    x"0417DE08",
    x"0417A2C1",
    x"04176791",
    x"04172C78",
    x"0416F176",
    x"0416B68B",
    x"04167BB7",
    x"041640FA",
    x"04160654",
    x"0415CBC5",
    x"0415914D",
    x"041556EC",
    x"04151CA1",
    x"0414E26E",
    x"0414A850",
    x"04146E4A",
    x"0414345A",
    x"0413FA81",
    x"0413C0BF",
    x"04138713",
    x"04134D7D",
    x"041313FE",
    x"0412DA95",
    x"0412A143",
    x"04126807",
    x"04122EE2",
    x"0411F5D3",
    x"0411BCDA",
    x"041183F7",
    x"04114B2B",
    x"04111274",
    x"0410D9D4",
    x"0410A14A",
    x"041068D6",
    x"04103078",
    x"040FF830",
    x"040FBFFE",
    x"040F87E2",
    x"040F4FDC",
    x"040F17EC",
    x"040EE012",
    x"040EA84D",
    x"040E709E",
    x"040E3905",
    x"040E0181",
    x"040DCA14",
    x"040D92BC",
    x"040D5B79",
    x"040D244C",
    x"040CED35",
    x"040CB633",
    x"040C7F46",
    x"040C486F",
    x"040C11AE",
    x"040BDB02",
    x"040BA46B",
    x"040B6DE9",
    x"040B377D",
    x"040B0126",
    x"040ACAE4",
    x"040A94B7",
    x"040A5EA0",
    x"040A289D",
    x"0409F2B0",
    x"0409BCD8",
    x"04098714",
    x"04095166",
    x"04091BCD",
    x"0408E648",
    x"0408B0D9",
    x"04087B7E",
    x"04084638",
    x"04081107",
    x"0407DBEB",
    x"0407A6E4",
    x"040771F1",
    x"04073D12",
    x"04070849",
    x"0406D394",
    x"04069EF4",
    x"04066A68",
    x"040635F1",
    x"0406018E",
    x"0405CD3F",
    x"04059905",
    x"040564E0",
    x"040530CE",
    x"0404FCD2",
    x"0404C8E9",
    x"04049515",
    x"04046154",
    x"04042DA9",
    x"0403FA11",
    x"0403C68D",
    x"0403931E",
    x"04035FC2",
    x"04032C7B",
    x"0402F947",
    x"0402C628",
    x"0402931D",
    x"04026025",
    x"04022D42",
    x"0401FA72",
    x"0401C7B6",
    x"0401950E",
    x"04016279",
    x"04012FF9",
    x"0400FD8C",
    x"0400CB33",
    x"040098ED",
    x"040066BB",
    x"0400349D",
    x"04000292",
    x"03FFA136",
    x"03FF3D6E",
    x"03FED9CE",
    x"03FE7654",
    x"03FE1301",
    x"03FDAFD5",
    x"03FD4CD0",
    x"03FCE9F1",
    x"03FC8739",
    x"03FC24A8",
    x"03FBC23C",
    x"03FB5FF8",
    x"03FAFDD9",
    x"03FA9BE1",
    x"03FA3A10",
    x"03F9D864",
    x"03F976DF",
    x"03F9157F",
    x"03F8B446",
    x"03F85332",
    x"03F7F245",
    x"03F7917D",
    x"03F730DB",
    x"03F6D05F",
    x"03F67008",
    x"03F60FD7",
    x"03F5AFCC",
    x"03F54FE6",
    x"03F4F025",
    x"03F4908A",
    x"03F43114",
    x"03F3D1C4",
    x"03F37299",
    x"03F31392",
    x"03F2B4B1",
    x"03F255F5",
    x"03F1F75E",
    x"03F198EC",
    x"03F13A9F",
    x"03F0DC76",
    x"03F07E72",
    x"03F02093",
    x"03EFC2D9",
    x"03EF6543",
    x"03EF07D2",
    x"03EEAA85",
    x"03EE4D5D",
    x"03EDF058",
    x"03ED9379",
    x"03ED36BD",
    x"03ECDA26",
    x"03EC7DB3",
    x"03EC2164",
    x"03EBC539",
    x"03EB6932",
    x"03EB0D4F",
    x"03EAB18F",
    x"03EA55F4",
    x"03E9FA7C",
    x"03E99F28",
    x"03E943F8",
    x"03E8E8EB",
    x"03E88E02",
    x"03E8333C",
    x"03E7D89A",
    x"03E77E1B",
    x"03E723BF",
    x"03E6C987",
    x"03E66F72",
    x"03E61580",
    x"03E5BBB1",
    x"03E56205",
    x"03E5087C",
    x"03E4AF16",
    x"03E455D3",
    x"03E3FCB3",
    x"03E3A3B6",
    x"03E34ADB",
    x"03E2F224",
    x"03E2998E",
    x"03E2411C",
    x"03E1E8CB",
    x"03E1909E",
    x"03E13892",
    x"03E0E0A9",
    x"03E088E3",
    x"03E0313E",
    x"03DFD9BC",
    x"03DF825C",
    x"03DF2B1E",
    x"03DED403",
    x"03DE7D09",
    x"03DE2631",
    x"03DDCF7B",
    x"03DD78E7",
    x"03DD2274",
    x"03DCCC24",
    x"03DC75F5",
    x"03DC1FE8",
    x"03DBC9FC",
    x"03DB7432",
    x"03DB1E89",
    x"03DAC902",
    x"03DA739C",
    x"03DA1E58",
    x"03D9C934",
    x"03D97432",
    x"03D91F52",
    x"03D8CA92",
    x"03D875F3",
    x"03D82176",
    x"03D7CD19",
    x"03D778DE",
    x"03D724C3",
    x"03D6D0C9",
    x"03D67CF0",
    x"03D62937",
    x"03D5D59F",
    x"03D58228",
    x"03D52ED2",
    x"03D4DB9C",
    x"03D48886",
    x"03D43591",
    x"03D3E2BC",
    x"03D39008",
    x"03D33D74",
    x"03D2EB00",
    x"03D298AC",
    x"03D24679",
    x"03D1F465",
    x"03D1A272",
    x"03D1509E",
    x"03D0FEEB",
    x"03D0AD57",
    x"03D05BE3",
    x"03D00A8F",
    x"03CFB95B",
    x"03CF6846",
    x"03CF1751",
    x"03CEC67C",
    x"03CE75C6",
    x"03CE2530",
    x"03CDD4B9",
    x"03CD8462",
    x"03CD342A",
    x"03CCE411",
    x"03CC9418",
    x"03CC443D",
    x"03CBF482",
    x"03CBA4E6",
    x"03CB5569",
    x"03CB060C",
    x"03CAB6CD",
    x"03CA67AD",
    x"03CA18AC",
    x"03C9C9CA",
    x"03C97B06",
    x"03C92C61",
    x"03C8DDDB",
    x"03C88F74",
    x"03C8412B",
    x"03C7F301",
    x"03C7A4F5",
    x"03C75708",
    x"03C70939",
    x"03C6BB89",
    x"03C66DF7",
    x"03C62083",
    x"03C5D32D",
    x"03C585F6",
    x"03C538DD",
    x"03C4EBE2",
    x"03C49F05",
    x"03C45245",
    x"03C405A4",
    x"03C3B921",
    x"03C36CBC",
    x"03C32074",
    x"03C2D44A",
    x"03C2883E",
    x"03C23C50",
    x"03C1F07F",
    x"03C1A4CC",
    x"03C15936",
    x"03C10DBE",
    x"03C0C263",
    x"03C07726",
    x"03C02C06",
    x"03BFE104",
    x"03BF961F",
    x"03BF4B57",
    x"03BF00AC",
    x"03BEB61E",
    x"03BE6BAD",
    x"03BE215A",
    x"03BDD723",
    x"03BD8D0A",
    x"03BD430D",
    x"03BCF92D",
    x"03BCAF6A",
    x"03BC65C4",
    x"03BC1C3B",
    x"03BBD2CE",
    x"03BB897E",
    x"03BB404B",
    x"03BAF734",
    x"03BAAE3A",
    x"03BA655C",
    x"03BA1C9A",
    x"03B9D3F6",
    x"03B98B6D",
    x"03B94301",
    x"03B8FAB1",
    x"03B8B27D",
    x"03B86A65",
    x"03B8226A",
    x"03B7DA8A",
    x"03B792C7",
    x"03B74B1F",
    x"03B70394",
    x"03B6BC25",
    x"03B674D1",
    x"03B62D99",
    x"03B5E67D",
    x"03B59F7D",
    x"03B55899",
    x"03B511D0",
    x"03B4CB23",
    x"03B48491",
    x"03B43E1B",
    x"03B3F7C1",
    x"03B3B182",
    x"03B36B5E",
    x"03B32556",
    x"03B2DF69",
    x"03B29997",
    x"03B253E1",
    x"03B20E46",
    x"03B1C8C6",
    x"03B18361",
    x"03B13E17",
    x"03B0F8E8",
    x"03B0B3D5",
    x"03B06EDC",
    x"03B029FE",
    x"03AFE53B",
    x"03AFA093",
    x"03AF5C06",
    x"03AF1793",
    x"03AED33B",
    x"03AE8EFE",
    x"03AE4ADB",
    x"03AE06D3",
    x"03ADC2E6",
    x"03AD7F13",
    x"03AD3B5B",
    x"03ACF7BD",
    x"03ACB439",
    x"03AC70D0",
    x"03AC2D81",
    x"03ABEA4C",
    x"03ABA732",
    x"03AB6432",
    x"03AB214C",
    x"03AADE80",
    x"03AA9BCE",
    x"03AA5936",
    x"03AA16B8",
    x"03A9D454",
    x"03A9920A",
    x"03A94FDA",
    x"03A90DC4",
    x"03A8CBC7",
    x"03A889E5",
    x"03A8481C",
    x"03A8066C",
    x"03A7C4D7",
    x"03A7835B",
    x"03A741F8",
    x"03A700AF",
    x"03A6BF7F",
    x"03A67E69",
    x"03A63D6D",
    x"03A5FC89",
    x"03A5BBBF",
    x"03A57B0F",
    x"03A53A77",
    x"03A4F9F9",
    x"03A4B994",
    x"03A47948",
    x"03A43915",
    x"03A3F8FB",
    x"03A3B8FB",
    x"03A37913",
    x"03A33944",
    x"03A2F98E",
    x"03A2B9F1",
    x"03A27A6D",
    x"03A23B01",
    x"03A1FBAF",
    x"03A1BC75",
    x"03A17D53",
    x"03A13E4B",
    x"03A0FF5B",
    x"03A0C083",
    x"03A081C4",
    x"03A0431E",
    x"03A00490",
    x"039FC61A",
    x"039F87BD",
    x"039F4978",
    x"039F0B4C",
    x"039ECD37",
    x"039E8F3B",
    x"039E5158",
    x"039E138C",
    x"039DD5D8",
    x"039D983D",
    x"039D5AB9",
    x"039D1D4E",
    x"039CDFFA",
    x"039CA2BF",
    x"039C659B",
    x"039C288F",
    x"039BEB9C",
    x"039BAEBF",
    x"039B71FB",
    x"039B354E",
    x"039AF8B9",
    x"039ABC3C",
    x"039A7FD6",
    x"039A4388",
    x"039A0752",
    x"0399CB32",
    x"03998F2B",
    x"0399533B",
    x"03991762",
    x"0398DBA0",
    x"03989FF6",
    x"03986463",
    x"039828E8",
    x"0397ED83",
    x"0397B236",
    x"03977700",
    x"03973BE1",
    x"039700D9",
    x"0396C5E8",
    x"03968B0F",
    x"0396504C",
    x"039615A0",
    x"0395DB0B",
    x"0395A08D",
    x"03956625",
    x"03952BD5",
    x"0394F19B",
    x"0394B778",
    x"03947D6C",
    x"03944376",
    x"03940997",
    x"0393CFCF",
    x"0393961D",
    x"03935C81",
    x"039322FD",
    x"0392E98E",
    x"0392B036",
    x"039276F4",
    x"03923DC9",
    x"039204B4",
    x"0391CBB5",
    x"039192CD",
    x"039159FB",
    x"0391213F",
    x"0390E899",
    x"0390B009",
    x"0390778F",
    x"03903F2C",
    x"039006DE",
    x"038FCEA6",
    x"038F9684",
    x"038F5E79",
    x"038F2683",
    x"038EEEA2",
    x"038EB6D8",
    x"038E7F24",
    x"038E4785",
    x"038E0FFC",
    x"038DD888",
    x"038DA12B",
    x"038D69E2",
    x"038D32B0",
    x"038CFB93",
    x"038CC48B",
    x"038C8D99",
    x"038C56BD",
    x"038C1FF5",
    x"038BE944",
    x"038BB2A7",
    x"038B7C20",
    x"038B45AE",
    x"038B0F52",
    x"038AD90A",
    x"038AA2D8",
    x"038A6CBB",
    x"038A36B3",
    x"038A00C0",
    x"0389CAE2",
    x"0389951A",
    x"03895F66",
    x"038929C7",
    x"0388F43D",
    x"0388BEC8",
    x"03888968",
    x"0388541D",
    x"03881EE7",
    x"0387E9C5",
    x"0387B4B8",
    x"03877FC0",
    x"03874ADC",
    x"0387160D",
    x"0386E153",
    x"0386ACAD",
    x"0386781C",
    x"0386439F",
    x"03860F37",
    x"0385DAE3",
    x"0385A6A4",
    x"03857279",
    x"03853E63",
    x"03850A60",
    x"0384D672",
    x"0384A299",
    x"03846ED3",
    x"03843B22",
    x"03840785",
    x"0383D3FC",
    x"0383A088",
    x"03836D27",
    x"038339DA",
    x"038306A2",
    x"0382D37D",
    x"0382A06D",
    x"03826D70",
    x"03823A87",
    x"038207B2",
    x"0381D4F1",
    x"0381A244",
    x"03816FAA",
    x"03813D24",
    x"03810AB2",
    x"0380D854",
    x"0380A609",
    x"038073D2",
    x"038041AF",
    x"03800F9F",
    x"037FBB45",
    x"037F5774",
    x"037EF3C9",
    x"037E9045",
    x"037E2CE8",
    x"037DC9B2",
    x"037D66A3",
    x"037D03BA",
    x"037CA0F8",
    x"037C3E5C",
    x"037BDBE7",
    x"037B7998",
    x"037B1770",
    x"037AB56E",
    x"037A5392",
    x"0379F1DD",
    x"0379904D",
    x"03792EE4",
    x"0378CDA1",
    x"03786C83",
    x"03780B8C",
    x"0377AABA",
    x"03774A0E",
    x"0376E988",
    x"03768928",
    x"037628ED",
    x"0375C8D8",
    x"037568E8",
    x"0375091E",
    x"0374A979",
    x"037449FA",
    x"0373EA9F",
    x"03738B6A",
    x"03732C5A",
    x"0372CD70",
    x"03726EAA",
    x"03721009",
    x"0371B18D",
    x"03715336",
    x"0370F504",
    x"037096F7",
    x"0370390E",
    x"036FDB4A",
    x"036F7DAB",
    x"036F2030",
    x"036EC2DA",
    x"036E65A8",
    x"036E089A",
    x"036DABB1",
    x"036D4EEC",
    x"036CF24C",
    x"036C95CF",
    x"036C3976",
    x"036BDD42",
    x"036B8132",
    x"036B2545",
    x"036AC97C",
    x"036A6DD8",
    x"036A1257",
    x"0369B6F9",
    x"03695BC0",
    x"036900AA",
    x"0368A5B7",
    x"03684AE8",
    x"0367F03D",
    x"036795B4",
    x"03673B50",
    x"0366E10E",
    x"036686F0",
    x"03662CF5",
    x"0365D31D",
    x"03657968",
    x"03651FD6",
    x"0364C667",
    x"03646D1B",
    x"036413F2",
    x"0363BAEB",
    x"03636207",
    x"03630947",
    x"0362B0A8",
    x"0362582D",
    x"0361FFD3",
    x"0361A79D",
    x"03614F88",
    x"0360F796",
    x"03609FC7",
    x"0360481A",
    x"035FF08F",
    x"035F9926",
    x"035F41DF",
    x"035EEABA",
    x"035E93B8",
    x"035E3CD7",
    x"035DE618",
    x"035D8F7B",
    x"035D3900",
    x"035CE2A6",
    x"035C8C6F",
    x"035C3659",
    x"035BE064",
    x"035B8A91",
    x"035B34E0",
    x"035ADF50",
    x"035A89E2",
    x"035A3494",
    x"0359DF68",
    x"03598A5E",
    x"03593574",
    x"0358E0AC",
    x"03588C05",
    x"0358377F",
    x"0357E319",
    x"03578ED5",
    x"03573AB2",
    x"0356E6AF",
    x"035692CE",
    x"03563F0D",
    x"0355EB6C",
    x"035597ED",
    x"0355448E",
    x"0354F14F",
    x"03549E31",
    x"03544B33",
    x"0353F856",
    x"0353A599",
    x"035352FD",
    x"03530081",
    x"0352AE24",
    x"03525BE9",
    x"035209CD",
    x"0351B7D1",
    x"035165F5",
    x"03511439",
    x"0350C29D",
    x"03507121",
    x"03501FC5",
    x"034FCE88",
    x"034F7D6B",
    x"034F2C6E",
    x"034EDB91",
    x"034E8AD3",
    x"034E3A34",
    x"034DE9B5",
    x"034D9956",
    x"034D4915",
    x"034CF8F5",
    x"034CA8F3",
    x"034C5911",
    x"034C094D",
    x"034BB9A9",
    x"034B6A24",
    x"034B1ABE",
    x"034ACB77",
    x"034A7C4F",
    x"034A2D46",
    x"0349DE5C",
    x"03498F90",
    x"034940E4",
    x"0348F256",
    x"0348A3E6",
    x"03485596",
    x"03480764",
    x"0347B950",
    x"03476B5B",
    x"03471D84",
    x"0346CFCC",
    x"03468232",
    x"034634B6",
    x"0345E758",
    x"03459A19",
    x"03454CF8",
    x"0344FFF5",
    x"0344B310",
    x"03446649",
    x"034419A0",
    x"0343CD15",
    x"034380A8",
    x"03433459",
    x"0342E827",
    x"03429C13",
    x"0342501D",
    x"03420445",
    x"0341B88A",
    x"03416CEC",
    x"0341216D",
    x"0340D60A",
    x"03408AC5",
    x"03403F9E",
    x"033FF494",
    x"033FA9A7",
    x"033F5ED7",
    x"033F1425",
    x"033EC98F",
    x"033E7F17",
    x"033E34BC",
    x"033DEA7E",
    x"033DA05D",
    x"033D5659",
    x"033D0C71",
    x"033CC2A7",
    x"033C78F9",
    x"033C2F68",
    x"033BE5F4",
    x"033B9C9D",
    x"033B5362",
    x"033B0A44",
    x"033AC142",
    x"033A785D",
    x"033A2F94",
    x"0339E6E7",
    x"03399E57",
    x"033955E4",
    x"03390D8C",
    x"0338C551",
    x"03387D32",
    x"0338352F",
    x"0337ED49",
    x"0337A57E",
    x"03375DCF",
    x"0337163D",
    x"0336CEC6",
    x"0336876B",
    x"0336402C",
    x"0335F909",
    x"0335B201",
    x"03356B16",
    x"03352446",
    x"0334DD91",
    x"033496F9",
    x"0334507B",
    x"03340A1A",
    x"0333C3D4",
    x"03337DA9",
    x"03333799",
    x"0332F1A5",
    x"0332ABCD",
    x"0332660F",
    x"0332206D",
    x"0331DAE6",
    x"0331957A",
    x"03315029",
    x"03310AF3",
    x"0330C5D8",
    x"033080D9",
    x"03303BF4",
    x"032FF72A",
    x"032FB27B",
    x"032F6DE6",
    x"032F296D",
    x"032EE50E",
    x"032EA0CA",
    x"032E5CA0",
    x"032E1891",
    x"032DD49D",
    x"032D90C3",
    x"032D4D04",
    x"032D095F",
    x"032CC5D5",
    x"032C8265",
    x"032C3F0F",
    x"032BFBD3",
    x"032BB8B2",
    x"032B75AB",
    x"032B32BE",
    x"032AEFEB",
    x"032AAD33",
    x"032A6A94",
    x"032A280F",
    x"0329E5A5",
    x"0329A354",
    x"0329611D",
    x"03291F00",
    x"0328DCFD",
    x"03289B13",
    x"03285944",
    x"0328178E",
    x"0327D5F1",
    x"0327946E",
    x"03275305",
    x"032711B6",
    x"0326D07F",
    x"03268F63",
    x"03264E5F",
    x"03260D75",
    x"0325CCA5",
    x"03258BEE",
    x"03254B50",
    x"03250ACB",
    x"0324CA5F",
    x"03248A0D",
    x"032449D3",
    x"032409B3",
    x"0323C9AC",
    x"032389BD",
    x"032349E8",
    x"03230A2C",
    x"0322CA88",
    x"03228AFD",
    x"03224B8B",
    x"03220C32",
    x"0321CCF2",
    x"03218DCA",
    x"03214EBB",
    x"03210FC5",
    x"0320D0E7",
    x"03209221",
    x"03205375",
    x"032014E0",
    x"031FD664",
    x"031F9801",
    x"031F59B6",
    x"031F1B83",
    x"031EDD68",
    x"031E9F66",
    x"031E617B",
    x"031E23A9",
    x"031DE5F0",
    x"031DA84E",
    x"031D6AC4",
    x"031D2D52",
    x"031CEFF9",
    x"031CB2B7",
    x"031C758D",
    x"031C387B",
    x"031BFB81",
    x"031BBE9F",
    x"031B81D4",
    x"031B4521",
    x"031B0886",
    x"031ACC02",
    x"031A8F97",
    x"031A5342",
    x"031A1705",
    x"0319DAE0",
    x"03199ED2",
    x"031962DC",
    x"031926FD",
    x"0318EB36",
    x"0318AF85",
    x"031873ED",
    x"0318386B",
    x"0317FD00",
    x"0317C1AD",
    x"03178671",
    x"03174B4C",
    x"0317103E",
    x"0316D547",
    x"03169A68",
    x"03165F9F",
    x"031624ED",
    x"0315EA52",
    x"0315AFCE",
    x"03157561",
    x"03153B0A",
    x"031500CA",
    x"0314C6A2",
    x"03148C8F",
    x"03145294",
    x"031418AF",
    x"0313DEE0",
    x"0313A529",
    x"03136B87",
    x"031331FD",
    x"0312F888",
    x"0312BF2A",
    x"031285E3",
    x"03124CB2",
    x"03121397",
    x"0311DA93",
    x"0311A1A4",
    x"031168CC",
    x"0311300A",
    x"0310F75F",
    x"0310BEC9",
    x"0310864A",
    x"03104DE0",
    x"0310158D",
    x"030FDD4F",
    x"030FA528",
    x"030F6D16",
    x"030F351B",
    x"030EFD35",
    x"030EC565",
    x"030E8DAB",
    x"030E5606",
    x"030E1E77",
    x"030DE6FE",
    x"030DAF9B",
    x"030D784D",
    x"030D4115",
    x"030D09F2",
    x"030CD2E5",
    x"030C9BED",
    x"030C650B",
    x"030C2E3F",
    x"030BF787",
    x"030BC0E5",
    x"030B8A58",
    x"030B53E1",
    x"030B1D7F",
    x"030AE732",
    x"030AB0FA",
    x"030A7AD8",
    x"030A44CA",
    x"030A0ED2",
    x"0309D8EF",
    x"0309A320",
    x"03096D67",
    x"030937C3",
    x"03090234",
    x"0308CCB9",
    x"03089754",
    x"03086203",
    x"03082CC7",
    x"0307F7A0",
    x"0307C28E",
    x"03078D90",
    x"030758A7",
    x"030723D3",
    x"0306EF13",
    x"0306BA68",
    x"030685D1",
    x"0306514F",
    x"03061CE2",
    x"0305E889",
    x"0305B444",
    x"03058014",
    x"03054BF8",
    x"030517F1",
    x"0304E3FD",
    x"0304B01E",
    x"03047C54",
    x"0304489D",
    x"030414FB",
    x"0303E16D",
    x"0303ADF3",
    x"03037A8D",
    x"0303473B",
    x"030313FD",
    x"0302E0D4",
    x"0302ADBE",
    x"03027ABC",
    x"030247CE",
    x"030214F4",
    x"0301E22D",
    x"0301AF7B",
    x"03017CDC",
    x"03014A51",
    x"030117DA",
    x"0300E577",
    x"0300B327",
    x"030080EB",
    x"03004EC2",
    x"03001CAD",
    x"02FFD558",
    x"02FF717C",
    x"02FF0DC7",
    x"02FEAA39",
    x"02FE46D2",
    x"02FDE392",
    x"02FD8078",
    x"02FD1D85",
    x"02FCBAB9",
    x"02FC5813",
    x"02FBF594",
    x"02FB933C",
    x"02FB3109",
    x"02FACEFD",
    x"02FA6D18",
    x"02FA0B58",
    x"02F9A9BF",
    x"02F9484B",
    x"02F8E6FE",
    x"02F885D7",
    x"02F824D6",
    x"02F7C3FA",
    x"02F76344",
    x"02F702B5",
    x"02F6A24A",
    x"02F64206",
    x"02F5E1E7",
    x"02F581ED",
    x"02F52219",
    x"02F4C26B",
    x"02F462E1",
    x"02F4037D",
    x"02F3A43F",
    x"02F34525",
    x"02F2E630",
    x"02F28761",
    x"02F228B7",
    x"02F1CA31",
    x"02F16BD1",
    x"02F10D95",
    x"02F0AF7E",
    x"02F0518C",
    x"02EFF3BE",
    x"02EF9615",
    x"02EF3891",
    x"02EEDB31",
    x"02EE7DF6",
    x"02EE20DF",
    x"02EDC3EC",
    x"02ED671E",
    x"02ED0A74",
    x"02ECADEE",
    x"02EC518C",
    x"02EBF54E",
    x"02EB9934",
    x"02EB3D3E",
    x"02EAE16C",
    x"02EA85BE",
    x"02EA2A34",
    x"02E9CECD",
    x"02E9738A",
    x"02E9186B",
    x"02E8BD6F",
    x"02E86297",
    x"02E807E2",
    x"02E7AD51",
    x"02E752E2",
    x"02E6F898",
    x"02E69E70",
    x"02E6446C",
    x"02E5EA8B",
    x"02E590CD",
    x"02E53732",
    x"02E4DDBA",
    x"02E48464",
    x"02E42B32",
    x"02E3D223",
    x"02E37936",
    x"02E3206C",
    x"02E2C7C5",
    x"02E26F40",
    x"02E216DE",
    x"02E1BE9E",
    x"02E16681",
    x"02E10E86",
    x"02E0B6AD",
    x"02E05EF7",
    x"02E00763",
    x"02DFAFF1",
    x"02DF58A2",
    x"02DF0174",
    x"02DEAA69",
    x"02DE537F",
    x"02DDFCB7",
    x"02DDA611",
    x"02DD4F8D",
    x"02DCF92B",
    x"02DCA2EB",
    x"02DC4CCC",
    x"02DBF6CF",
    x"02DBA0F3",
    x"02DB4B39",
    x"02DAF5A0",
    x"02DAA029",
    x"02DA4AD3",
    x"02D9F59F",
    x"02D9A08B",
    x"02D94B99",
    x"02D8F6C8",
    x"02D8A218",
    x"02D84D8A",
    x"02D7F91C",
    x"02D7A4CF",
    x"02D750A3",
    x"02D6FC98",
    x"02D6A8AE",
    x"02D654E4",
    x"02D6013B",
    x"02D5ADB3",
    x"02D55A4C",
    x"02D50705",
    x"02D4B3DE",
    x"02D460D8",
    x"02D40DF2",
    x"02D3BB2D",
    x"02D36888",
    x"02D31603",
    x"02D2C39F",
    x"02D2715B",
    x"02D21F36",
    x"02D1CD32",
    x"02D17B4E",
    x"02D1298A",
    x"02D0D7E6",
    x"02D08661",
    x"02D034FD",
    x"02CFE3B8",
    x"02CF9293",
    x"02CF418D",
    x"02CEF0A7",
    x"02CE9FE1",
    x"02CE4F3B",
    x"02CDFEB3",
    x"02CDAE4C",
    x"02CD5E03",
    x"02CD0DDA",
    x"02CCBDD0",
    x"02CC6DE6",
    x"02CC1E1A",
    x"02CBCE6E",
    x"02CB7EE1",
    x"02CB2F73",
    x"02CAE024",
    x"02CA90F4",
    x"02CA41E3",
    x"02C9F2F0",
    x"02C9A41D",
    x"02C95568",
    x"02C906D2",
    x"02C8B85B",
    x"02C86A02",
    x"02C81BC8",
    x"02C7CDAC",
    x"02C77FAF",
    x"02C731D1",
    x"02C6E410",
    x"02C6966F",
    x"02C648EB",
    x"02C5FB86",
    x"02C5AE3E",
    x"02C56115",
    x"02C5140B",
    x"02C4C71E",
    x"02C47A4F",
    x"02C42D9E",
    x"02C3E10B",
    x"02C39496",
    x"02C3483F",
    x"02C2FC06",
    x"02C2AFEA",
    x"02C263EC",
    x"02C2180C",
    x"02C1CC4A",
    x"02C180A5",
    x"02C1351D",
    x"02C0E9B3",
    x"02C09E67",
    x"02C05337",
    x"02C00825",
    x"02BFBD31",
    x"02BF725A",
    x"02BF27A0",
    x"02BEDD03",
    x"02BE9283",
    x"02BE4820",
    x"02BDFDDB",
    x"02BDB3B2",
    x"02BD69A6",
    x"02BD1FB7",
    x"02BCD5E5",
    x"02BC8C30",
    x"02BC4298",
    x"02BBF91C",
    x"02BBAFBD",
    x"02BB667B",
    x"02BB1D55",
    x"02BAD44C",
    x"02BA8B5F",
    x"02BA428F",
    x"02B9F9DB",
    x"02B9B144",
    x"02B968C9",
    x"02B9206A",
    x"02B8D827",
    x"02B89001",
    x"02B847F7",
    x"02B80009",
    x"02B7B837",
    x"02B77081",
    x"02B728E7",
    x"02B6E169",
    x"02B69A07",
    x"02B652C1",
    x"02B60B96",
    x"02B5C487",
    x"02B57D95",
    x"02B536BD",
    x"02B4F002",
    x"02B4A962",
    x"02B462DD",
    x"02B41C75",
    x"02B3D627",
    x"02B38FF5",
    x"02B349DF",
    x"02B303E4",
    x"02B2BE04",
    x"02B2783F",
    x"02B23296",
    x"02B1ED08",
    x"02B1A795",
    x"02B1623D",
    x"02B11D00",
    x"02B0D7DE",
    x"02B092D7",
    x"02B04DEB",
    x"02B0091A",
    x"02AFC464",
    x"02AF7FC9",
    x"02AF3B48",
    x"02AEF6E2",
    x"02AEB297",
    x"02AE6E67",
    x"02AE2A51",
    x"02ADE656",
    x"02ADA275",
    x"02AD5EAF",
    x"02AD1B03",
    x"02ACD772",
    x"02AC93FB",
    x"02AC509E",
    x"02AC0D5C",
    x"02ABCA34",
    x"02AB8726",
    x"02AB4432",
    x"02AB0159",
    x"02AABE99",
    x"02AA7BF4",
    x"02AA3968",
    x"02A9F6F7",
    x"02A9B49F",
    x"02A97262",
    x"02A9303E",
    x"02A8EE34",
    x"02A8AC44",
    x"02A86A6D",
    x"02A828B1",
    x"02A7E70E",
    x"02A7A584",
    x"02A76414",
    x"02A722BE",
    x"02A6E181",
    x"02A6A05E",
    x"02A65F54",
    x"02A61E63",
    x"02A5DD8C",
    x"02A59CCE",
    x"02A55C29",
    x"02A51B9E",
    x"02A4DB2C",
    x"02A49AD3",
    x"02A45A93",
    x"02A41A6C",
    x"02A3DA5E",
    x"02A39A69",
    x"02A35A8E",
    x"02A31ACB",
    x"02A2DB21",
    x"02A29B90",
    x"02A25C17",
    x"02A21CB8",
    x"02A1DD71",
    x"02A19E43",
    x"02A15F2D",
    x"02A12030",
    x"02A0E14C",
    x"02A0A280",
    x"02A063CD",
    x"02A02532",
    x"029FE6B0",
    x"029FA846",
    x"029F69F4",
    x"029F2BBB",
    x"029EED9A",
    x"029EAF91",
    x"029E71A1",
    x"029E33C9",
    x"029DF609",
    x"029DB860",
    x"029D7AD0",
    x"029D3D59",
    x"029CFFF9",
    x"029CC2B1",
    x"029C8580",
    x"029C4868",
    x"029C0B68",
    x"029BCE7F",
    x"029B91AF",
    x"029B54F5",
    x"029B1854",
    x"029ADBCA",
    x"029A9F58",
    x"029A62FE",
    x"029A26BB",
    x"0299EA90",
    x"0299AE7C",
    x"0299727F",
    x"0299369A",
    x"0298FACD",
    x"0298BF16",
    x"02988377",
    x"029847F0",
    x"02980C7F",
    x"0297D126",
    x"029795E4",
    x"02975AB9",
    x"02971FA5",
    x"0296E4A8",
    x"0296A9C2",
    x"02966EF3",
    x"0296343C",
    x"0295F99B",
    x"0295BF11",
    x"0295849D",
    x"02954A41",
    x"02950FFB",
    x"0294D5CC",
    x"02949BB4",
    x"029461B3",
    x"029427C8",
    x"0293EDF4",
    x"0293B436",
    x"02937A8F",
    x"029340FE",
    x"02930784",
    x"0292CE20",
    x"029294D3",
    x"02925B9C",
    x"0292227B",
    x"0291E971",
    x"0291B07D",
    x"0291779F",
    x"02913ED8",
    x"02910626",
    x"0290CD8B",
    x"02909506",
    x"02905C96",
    x"0290243D",
    x"028FEBFA",
    x"028FB3CD",
    x"028F7BB6",
    x"028F43B4",
    x"028F0BC9",
    x"028ED3F3",
    x"028E9C33",
    x"028E6489",
    x"028E2CF4",
    x"028DF576",
    x"028DBE0D",
    x"028D86B9",
    x"028D4F7B",
    x"028D1853",
    x"028CE140",
    x"028CAA43",
    x"028C735B",
    x"028C3C89",
    x"028C05CC",
    x"028BCF25",
    x"028B9892",
    x"028B6215",
    x"028B2BAE",
    x"028AF55B",
    x"028ABF1E",
    x"028A88F6",
    x"028A52E3",
    x"028A1CE5",
    x"0289E6FC",
    x"0289B129",
    x"02897B6A",
    x"028945C0",
    x"0289102B",
    x"0288DAAC",
    x"0288A541",
    x"02886FEA",
    x"02883AA9",
    x"0288057D",
    x"0287D065",
    x"02879B62",
    x"02876673",
    x"0287319A",
    x"0286FCD5",
    x"0286C824",
    x"02869388",
    x"02865F01",
    x"02862A8E",
    x"0285F630",
    x"0285C1E6",
    x"02858DB0",
    x"0285598F",
    x"02852582",
    x"0284F18A",
    x"0284BDA5",
    x"028489D6",
    x"0284561A",
    x"02842272",
    x"0283EEDF",
    x"0283BB60",
    x"028387F4",
    x"0283549D",
    x"0283215A",
    x"0282EE2B",
    x"0282BB10",
    x"02828809",
    x"02825516",
    x"02822237",
    x"0281EF6B",
    x"0281BCB4",
    x"02818A10",
    x"02815780",
    x"02812503",
    x"0280F29B",
    x"0280C046",
    x"02808E05",
    x"02805BD7",
    x"028029BD",
    x"027FEF6D",
    x"027F8B87",
    x"027F27C8",
    x"027EC430",
    x"027E60BE",
    x"027DFD74",
    x"027D9A50",
    x"027D3753",
    x"027CD47D",
    x"027C71CD",
    x"027C0F44",
    x"027BACE1",
    x"027B4AA5",
    x"027AE88F",
    x"027A869F",
    x"027A24D6",
    x"0279C333",
    x"027961B5",
    x"0279005E",
    x"02789F2D",
    x"02783E22",
    x"0277DD3C",
    x"02777C7D",
    x"02771BE3",
    x"0276BB6F",
    x"02765B21",
    x"0275FAF8",
    x"02759AF5",
    x"02753B17",
    x"0274DB5E",
    x"02747BCB",
    x"02741C5E",
    x"0273BD15",
    x"02735DF2",
    x"0272FEF4",
    x"0272A01B",
    x"02724167",
    x"0271E2D8",
    x"0271846E",
    x"02712628",
    x"0270C808",
    x"02706A0C",
    x"02700C35",
    x"026FAE82",
    x"026F50F4",
    x"026EF38B",
    x"026E9646",
    x"026E3926",
    x"026DDC2A",
    x"026D7F52",
    x"026D229E",
    x"026CC60F",
    x"026C69A3",
    x"026C0D5C",
    x"026BB139",
    x"026B553A",
    x"026AF95E",
    x"026A9DA7",
    x"026A4213",
    x"0269E6A3",
    x"02698B57",
    x"0269302E",
    x"0268D529",
    x"02687A48",
    x"02681F8A",
    x"0267C4EF",
    x"02676A78",
    x"02671024",
    x"0266B5F3",
    x"02665BE6",
    x"026601FB",
    x"0265A834",
    x"02654E90",
    x"0264F50F",
    x"02649BB0",
    x"02644275",
    x"0263E95C",
    x"02639067",
    x"02633794",
    x"0262DEE3",
    x"02628656",
    x"02622DEA",
    x"0261D5A2",
    x"02617D7B",
    x"02612578",
    x"0260CD96",
    x"026075D7",
    x"02601E3A",
    x"025FC6BF",
    x"025F6F67",
    x"025F1830",
    x"025EC11C",
    x"025E6A29",
    x"025E1359",
    x"025DBCAA",
    x"025D661D",
    x"025D0FB2",
    x"025CB969",
    x"025C6342",
    x"025C0D3C",
    x"025BB757",
    x"025B6194",
    x"025B0BF3",
    x"025AB673",
    x"025A6114",
    x"025A0BD7",
    x"0259B6BB",
    x"025961C0",
    x"02590CE7",
    x"0258B82E",
    x"02586397",
    x"02580F20",
    x"0257BACB",
    x"02576696",
    x"02571283",
    x"0256BE90",
    x"02566ABE",
    x"0256170D",
    x"0255C37C",
    x"0255700C",
    x"02551CBC",
    x"0254C98D",
    x"0254767F",
    x"02542391",
    x"0253D0C3",
    x"02537E16",
    x"02532B89",
    x"0252D91C",
    x"025286CF",
    x"025234A2",
    x"0251E296",
    x"025190A9",
    x"02513EDD",
    x"0250ED30",
    x"02509BA3",
    x"02504A37",
    x"024FF8E9",
    x"024FA7BC",
    x"024F56AE",
    x"024F05C0",
    x"024EB4F2",
    x"024E6443",
    x"024E13B4",
    x"024DC344",
    x"024D72F3",
    x"024D22C2",
    x"024CD2B0",
    x"024C82BD",
    x"024C32EA",
    x"024BE335",
    x"024B93A0",
    x"024B442A",
    x"024AF4D3",
    x"024AA59B",
    x"024A5681",
    x"024A0787",
    x"0249B8AC",
    x"024969EF",
    x"02491B51",
    x"0248CCD1",
    x"02487E71",
    x"0248302F",
    x"0247E20B",
    x"02479406",
    x"0247461F",
    x"0246F857",
    x"0246AAAD",
    x"02465D22",
    x"02460FB5",
    x"0245C266",
    x"02457535",
    x"02452822",
    x"0244DB2D",
    x"02448E57",
    x"0244419E",
    x"0243F504",
    x"0243A887",
    x"02435C28",
    x"02430FE7",
    x"0242C3C3",
    x"024277BE",
    x"02422BD6",
    x"0241E00C",
    x"0241945F",
    x"024148D0",
    x"0240FD5E",
    x"0240B20A",
    x"024066D3",
    x"02401BB9",
    x"023FD0BD",
    x"023F85DE",
    x"023F3B1C",
    x"023EF078",
    x"023EA5F1",
    x"023E5B86",
    x"023E1139",
    x"023DC709",
    x"023D7CF6",
    x"023D32FF",
    x"023CE926",
    x"023C9F69",
    x"023C55C9",
    x"023C0C46",
    x"023BC2E0",
    x"023B7996",
    x"023B3069",
    x"023AE758",
    x"023A9E64",
    x"023A558C",
    x"023A0CD1",
    x"0239C432",
    x"02397BB0",
    x"0239334A",
    x"0238EB00",
    x"0238A2D2",
    x"02385AC0",
    x"023812CB",
    x"0237CAF2",
    x"02378334",
    x"02373B93",
    x"0236F40E",
    x"0236ACA4",
    x"02366557",
    x"02361E25",
    x"0235D70F",
    x"02359015",
    x"02354937",
    x"02350274",
    x"0234BBCD",
    x"02347541",
    x"02342ED1",
    x"0233E87D",
    x"0233A244",
    x"02335C26",
    x"02331624",
    x"0232D03D",
    x"02328A71",
    x"023244C0",
    x"0231FF2B",
    x"0231B9B1",
    x"02317452",
    x"02312F0E",
    x"0230E9E5",
    x"0230A4D7",
    x"02305FE5",
    x"02301B0D",
    x"022FD64F",
    x"022F91AD",
    x"022F4D26",
    x"022F08B9",
    x"022EC467",
    x"022E802F",
    x"022E3C13",
    x"022DF810",
    x"022DB429",
    x"022D705C",
    x"022D2CA9",
    x"022CE911",
    x"022CA593",
    x"022C622F",
    x"022C1EE6",
    x"022BDBB7",
    x"022B98A3",
    x"022B55A8",
    x"022B12C8",
    x"022AD001",
    x"022A8D55",
    x"022A4AC3",
    x"022A084B",
    x"0229C5EC",
    x"022983A8",
    x"0229417D",
    x"0228FF6D",
    x"0228BD76",
    x"02287B99",
    x"022839D5",
    x"0227F82C",
    x"0227B69B",
    x"02277525",
    x"022733C8",
    x"0226F284",
    x"0226B15A",
    x"0226704A",
    x"02262F53",
    x"0225EE75",
    x"0225ADB0",
    x"02256D05",
    x"02252C73",
    x"0224EBFA",
    x"0224AB9B",
    x"02246B54",
    x"02242B27",
    x"0223EB13",
    x"0223AB17",
    x"02236B35",
    x"02232B6C",
    x"0222EBBB",
    x"0222AC23",
    x"02226CA5",
    x"02222D3E",
    x"0221EDF1",
    x"0221AEBD",
    x"02216FA1",
    x"0221309D",
    x"0220F1B3",
    x"0220B2E1",
    x"02207427",
    x"02203586",
    x"021FF6FD",
    x"021FB88D",
    x"021F7A35",
    x"021F3BF5",
    x"021EFDCE",
    x"021EBFBF",
    x"021E81C8",
    x"021E43EA",
    x"021E0623",
    x"021DC875",
    x"021D8ADF",
    x"021D4D60",
    x"021D0FFA",
    x"021CD2AC",
    x"021C9575",
    x"021C5857",
    x"021C1B50",
    x"021BDE62",
    x"021BA18B",
    x"021B64CB",
    x"021B2824",
    x"021AEB94",
    x"021AAF1C",
    x"021A72BB",
    x"021A3672",
    x"0219FA41",
    x"0219BE27",
    x"02198224",
    x"02194639",
    x"02190A65",
    x"0218CEA9",
    x"02189304",
    x"02185776",
    x"02181BFF",
    x"0217E0A0",
    x"0217A558",
    x"02176A27",
    x"02172F0D",
    x"0216F40A",
    x"0216B91E",
    x"02167E4A",
    x"0216438C",
    x"021608E5",
    x"0215CE55",
    x"021593DC",
    x"02155979",
    x"02151F2E",
    x"0214E4F9",
    x"0214AADB",
    x"021470D3",
    x"021436E3",
    x"0213FD08",
    x"0213C345",
    x"02138998",
    x"02135001",
    x"02131681",
    x"0212DD18",
    x"0212A3C5",
    x"02126A88",
    x"02123161",
    x"0211F851",
    x"0211BF57",
    x"02118674",
    x"02114DA6",
    x"021114EF",
    x"0210DC4E",
    x"0210A3C3",
    x"02106B4E",
    x"021032EF",
    x"020FFAA6",
    x"020FC273",
    x"020F8A56",
    x"020F524F",
    x"020F1A5E",
    x"020EE283",
    x"020EAABD",
    x"020E730D",
    x"020E3B73",
    x"020E03EF",
    x"020DCC80",
    x"020D9527",
    x"020D5DE3",
    x"020D26B6",
    x"020CEF9D",
    x"020CB89A",
    x"020C81AD",
    x"020C4AD5",
    x"020C1413",
    x"020BDD65",
    x"020BA6CE",
    x"020B704B",
    x"020B39DE",
    x"020B0386",
    x"020ACD43",
    x"020A9715",
    x"020A60FD",
    x"020A2AFA",
    x"0209F50B",
    x"0209BF32",
    x"0209896E",
    x"020953BF",
    x"02091E25",
    x"0208E89F",
    x"0208B32F",
    x"02087DD3",
    x"0208488D",
    x"0208135B",
    x"0207DE3D",
    x"0207A935",
    x"02077441",
    x"02073F62",
    x"02070A98",
    x"0206D5E2",
    x"0206A141",
    x"02066CB4",
    x"0206383C",
    x"020603D8",
    x"0205CF89",
    x"02059B4E",
    x"02056727",
    x"02053315",
    x"0204FF17",
    x"0204CB2E",
    x"02049759",
    x"02046398",
    x"02042FEB",
    x"0203FC52",
    x"0203C8CE",
    x"0203955D",
    x"02036201",
    x"02032EB9",
    x"0202FB84",
    x"0202C864",
    x"02029558",
    x"02026260",
    x"02022F7B",
    x"0201FCAA",
    x"0201C9EE",
    x"02019745",
    x"020164AF",
    x"0201322E",
    x"0200FFC0",
    x"0200CD66",
    x"02009B20",
    x"020068ED",
    x"020036CE",
    x"020004C2",
    x"01FFA594",
    x"01FF41CB",
    x"01FEDE29",
    x"01FE7AAD",
    x"01FE1759",
    x"01FDB42B",
    x"01FD5124",
    x"01FCEE44",
    x"01FC8B8A",
    x"01FC28F7",
    x"01FBC68A",
    x"01FB6443",
    x"01FB0223",
    x"01FAA02A",
    x"01FA3E56",
    x"01F9DCA9",
    x"01F97B22",
    x"01F919C1",
    x"01F8B886",
    x"01F85771",
    x"01F7F681",
    x"01F795B8",
    x"01F73514",
    x"01F6D497",
    x"01F6743E",
    x"01F6140C",
    x"01F5B3FF",
    x"01F55417",
    x"01F4F455",
    x"01F494B8",
    x"01F43541",
    x"01F3D5EF",
    x"01F376C2",
    x"01F317BA",
    x"01F2B8D7",
    x"01F25A19",
    x"01F1FB81",
    x"01F19D0D",
    x"01F13EBE",
    x"01F0E094",
    x"01F0828E",
    x"01F024AE",
    x"01EFC6F2",
    x"01EF695A",
    x"01EF0BE7",
    x"01EEAE99",
    x"01EE516F",
    x"01EDF469",
    x"01ED9788",
    x"01ED3ACB",
    x"01ECDE32",
    x"01EC81BD",
    x"01EC256D",
    x"01EBC940",
    x"01EB6D37",
    x"01EB1153",
    x"01EAB592",
    x"01EA59F5",
    x"01E9FE7C",
    x"01E9A326",
    x"01E947F4",
    x"01E8ECE6",
    x"01E891FB",
    x"01E83734",
    x"01E7DC90",
    x"01E7820F",
    x"01E727B2",
    x"01E6CD78",
    x"01E67362",
    x"01E6196E",
    x"01E5BF9E",
    x"01E565F1",
    x"01E50C66",
    x"01E4B2FF",
    x"01E459BA",
    x"01E40099",
    x"01E3A79A",
    x"01E34EBE",
    x"01E2F604",
    x"01E29D6E",
    x"01E244F9",
    x"01E1ECA8",
    x"01E19478",
    x"01E13C6C",
    x"01E0E481",
    x"01E08CB9",
    x"01E03513",
    x"01DFDD90",
    x"01DF862E",
    x"01DF2EEF",
    x"01DED7D1",
    x"01DE80D6",
    x"01DE29FD",
    x"01DDD345",
    x"01DD7CB0",
    x"01DD263C",
    x"01DCCFEA",
    x"01DC79B9",
    x"01DC23AB",
    x"01DBCDBE",
    x"01DB77F2",
    x"01DB2248",
    x"01DACCBF",
    x"01DA7758",
    x"01DA2212",
    x"01D9CCED",
    x"01D977EA",
    x"01D92308",
    x"01D8CE46",
    x"01D879A6",
    x"01D82527",
    x"01D7D0C9",
    x"01D77C8C",
    x"01D72870",
    x"01D6D475",
    x"01D6809A",
    x"01D62CE0",
    x"01D5D947",
    x"01D585CE",
    x"01D53276",
    x"01D4DF3F",
    x"01D48C28",
    x"01D43931",
    x"01D3E65B",
    x"01D393A5",
    x"01D34110",
    x"01D2EE9B",
    x"01D29C45",
    x"01D24A10",
    x"01D1F7FC",
    x"01D1A607",
    x"01D15432",
    x"01D1027D",
    x"01D0B0E8",
    x"01D05F73",
    x"01D00E1D",
    x"01CFBCE8",
    x"01CF6BD2",
    x"01CF1ADB",
    x"01CECA05",
    x"01CE794E",
    x"01CE28B6",
    x"01CDD83E",
    x"01CD87E5",
    x"01CD37AC",
    x"01CCE791",
    x"01CC9797",
    x"01CC47BB",
    x"01CBF7FF",
    x"01CBA861",
    x"01CB58E3",
    x"01CB0984",
    x"01CABA44",
    x"01CA6B22",
    x"01CA1C20",
    x"01C9CD3C",
    x"01C97E77",
    x"01C92FD1",
    x"01C8E14A",
    x"01C892E1",
    x"01C84497",
    x"01C7F66C",
    x"01C7A85F",
    x"01C75A70",
    x"01C70CA0",
    x"01C6BEEE",
    x"01C6715B",
    x"01C623E6",
    x"01C5D68F",
    x"01C58956",
    x"01C53C3C",
    x"01C4EF3F",
    x"01C4A261",
    x"01C455A0",
    x"01C408FE",
    x"01C3BC79",
    x"01C37012",
    x"01C323CA",
    x"01C2D79F",
    x"01C28B91",
    x"01C23FA1",
    x"01C1F3CF",
    x"01C1A81B",
    x"01C15C84",
    x"01C1110B",
    x"01C0C5AF",
    x"01C07A70",
    x"01C02F4F",
    x"01BFE44B",
    x"01BF9965",
    x"01BF4E9B",
    x"01BF03EF",
    x"01BEB960",
    x"01BE6EEE",
    x"01BE249A",
    x"01BDDA62",
    x"01BD9047",
    x"01BD4649",
    x"01BCFC68",
    x"01BCB2A4",
    x"01BC68FD",
    x"01BC1F72",
    x"01BBD604",
    x"01BB8CB3",
    x"01BB437E",
    x"01BAFA66",
    x"01BAB16A",
    x"01BA688B",
    x"01BA1FC9",
    x"01B9D722",
    x"01B98E99",
    x"01B9462B",
    x"01B8FDDA",
    x"01B8B5A5",
    x"01B86D8C",
    x"01B8258F",
    x"01B7DDAE",
    x"01B795EA",
    x"01B74E41",
    x"01B706B5",
    x"01B6BF44",
    x"01B677EF",
    x"01B630B6",
    x"01B5E999",
    x"01B5A298",
    x"01B55BB2",
    x"01B514E8",
    x"01B4CE3A",
    x"01B487A7",
    x"01B44130",
    x"01B3FAD4",
    x"01B3B494",
    x"01B36E6F",
    x"01B32866",
    x"01B2E277",
    x"01B29CA5",
    x"01B256ED",
    x"01B21151",
    x"01B1CBD0",
    x"01B18669",
    x"01B1411F",
    x"01B0FBEF",
    x"01B0B6DA",
    x"01B071E0",
    x"01B02D01",
    x"01AFE83D",
    x"01AFA393",
    x"01AF5F05",
    x"01AF1A91",
    x"01AED638",
    x"01AE91FA",
    x"01AE4DD6",
    x"01AE09CD",
    x"01ADC5DE",
    x"01AD820A",
    x"01AD3E51",
    x"01ACFAB2",
    x"01ACB72D",
    x"01AC73C2",
    x"01AC3072",
    x"01ABED3D",
    x"01ABAA21",
    x"01AB6720",
    x"01AB2438",
    x"01AAE16B",
    x"01AA9EB8",
    x"01AA5C1F",
    x"01AA19A0",
    x"01A9D73B",
    x"01A994F0",
    x"01A952BF",
    x"01A910A7",
    x"01A8CEAA",
    x"01A88CC6",
    x"01A84AFC",
    x"01A8094B",
    x"01A7C7B5",
    x"01A78637",
    x"01A744D4",
    x"01A7038A",
    x"01A6C259",
    x"01A68142",
    x"01A64044",
    x"01A5FF60",
    x"01A5BE94",
    x"01A57DE3",
    x"01A53D4A",
    x"01A4FCCB",
    x"01A4BC65",
    x"01A47C18",
    x"01A43BE4",
    x"01A3FBC9",
    x"01A3BBC7",
    x"01A37BDE",
    x"01A33C0E",
    x"01A2FC57",
    x"01A2BCB9",
    x"01A27D34",
    x"01A23DC7",
    x"01A1FE73",
    x"01A1BF38",
    x"01A18016",
    x"01A1410C",
    x"01A1021B",
    x"01A0C343",
    x"01A08483",
    x"01A045DB",
    x"01A0074C",
    x"019FC8D5",
    x"019F8A77",
    x"019F4C31",
    x"019F0E04",
    x"019ECFEE",
    x"019E91F1",
    x"019E540C",
    x"019E163F",
    x"019DD88B",
    x"019D9AEE",
    x"019D5D6A",
    x"019D1FFD",
    x"019CE2A9",
    x"019CA56C",
    x"019C6847",
    x"019C2B3B",
    x"019BEE46",
    x"019BB168",
    x"019B74A3",
    x"019B37F5",
    x"019AFB5F",
    x"019ABEE1",
    x"019A827A",
    x"019A462B",
    x"019A09F3",
    x"0199CDD3",
    x"019991CB",
    x"019955D9",
    x"019919FF",
    x"0198DE3D",
    x"0198A292",
    x"019866FE",
    x"01982B81",
    x"0197F01C",
    x"0197B4CE",
    x"01977997",
    x"01973E77",
    x"0197036E",
    x"0196C87C",
    x"01968DA1",
    x"019652DD",
    x"01961830",
    x"0195DD9A",
    x"0195A31B",
    x"019568B3",
    x"01952E62",
    x"0194F427",
    x"0194BA03",
    x"01947FF5",
    x"019445FF",
    x"01940C1F",
    x"0193D255",
    x"019398A2",
    x"01935F06",
    x"01932580",
    x"0192EC11",
    x"0192B2B8",
    x"01927975",
    x"01924049",
    x"01920733",
    x"0191CE33",
    x"0191954A",
    x"01915C77",
    x"019123BA",
    x"0190EB13",
    x"0190B282",
    x"01907A07",
    x"019041A3",
    x"01900954",
    x"018FD11B",
    x"018F98F9",
    x"018F60EC",
    x"018F28F5",
    x"018EF114",
    x"018EB948",
    x"018E8193",
    x"018E49F3",
    x"018E1269",
    x"018DDAF5",
    x"018DA396",
    x"018D6C4D",
    x"018D3519",
    x"018CFDFB",
    x"018CC6F3",
    x"018C9000",
    x"018C5923",
    x"018C225A",
    x"018BEBA8",
    x"018BB50A",
    x"018B7E82",
    x"018B480F",
    x"018B11B2",
    x"018ADB6A",
    x"018AA536",
    x"018A6F19",
    x"018A3910",
    x"018A031C",
    x"0189CD3D",
    x"01899774",
    x"018961BF",
    x"01892C1F",
    x"0188F694",
    x"0188C11F",
    x"01888BBE",
    x"01885671",
    x"0188213A",
    x"0187EC17",
    x"0187B70A",
    x"01878210",
    x"01874D2C",
    x"0187185C",
    x"0186E3A1",
    x"0186AEFA",
    x"01867A68",
    x"018645EB",
    x"01861182",
    x"0185DD2D",
    x"0185A8ED",
    x"018574C1",
    x"018540AA",
    x"01850CA6",
    x"0184D8B8",
    x"0184A4DD",
    x"01847117",
    x"01843D65",
    x"018409C7",
    x"0183D63D",
    x"0183A2C7",
    x"01836F66",
    x"01833C18",
    x"018308DF",
    x"0182D5B9",
    x"0182A2A8",
    x"01826FAA",
    x"01823CC1",
    x"018209EB",
    x"0181D729",
    x"0181A47B",
    x"018171E0",
    x"01813F5A",
    x"01810CE7",
    x"0180DA88",
    x"0180A83C",
    x"01807604",
    x"018043E0",
    x"018011CF",
    x"017FBFA4",
    x"017F5BD1",
    x"017EF824",
    x"017E949F",
    x"017E3140",
    x"017DCE08",
    x"017D6AF7",
    x"017D080D",
    x"017CA549",
    x"017C42AC",
    x"017BE035",
    x"017B7DE4",
    x"017B1BBA",
    x"017AB9B7",
    x"017A57D9",
    x"0179F622",
    x"01799491",
    x"01793326",
    x"0178D1E1",
    x"017870C2",
    x"01780FC9",
    x"0177AEF6",
    x"01774E48",
    x"0176EDC1",
    x"01768D5F",
    x"01762D22",
    x"0175CD0B",
    x"01756D1A",
    x"01750D4E",
    x"0174ADA7",
    x"01744E26",
    x"0173EECA",
    x"01738F94",
    x"01733082",
    x"0172D196",
    x"017272CE",
    x"0172142C",
    x"0171B5AF",
    x"01715756",
    x"0170F922",
    x"01709B13",
    x"01703D29",
    x"016FDF64",
    x"016F81C3",
    x"016F2446",
    x"016EC6EE",
    x"016E69BB",
    x"016E0CAC",
    x"016DAFC1",
    x"016D52FA",
    x"016CF658",
    x"016C99DA",
    x"016C3D80",
    x"016BE14A",
    x"016B8538",
    x"016B294A",
    x"016ACD80",
    x"016A71D9",
    x"016A1657",
    x"0169BAF8",
    x"01695FBD",
    x"016904A5",
    x"0168A9B1",
    x"01684EE0",
    x"0167F433",
    x"016799AA",
    x"01673F43",
    x"0166E500",
    x"01668AE0",
    x"016630E4",
    x"0165D70A",
    x"01657D54",
    x"016523C0",
    x"0164CA50",
    x"01647102",
    x"016417D7",
    x"0163BECF",
    x"016365EA",
    x"01630D28",
    x"0162B488",
    x"01625C0B",
    x"016203B0",
    x"0161AB78",
    x"01615362",
    x"0160FB6F",
    x"0160A39E",
    x"01604BEF",
    x"015FF462",
    x"015F9CF8",
    x"015F45B0",
    x"015EEE89",
    x"015E9785",
    x"015E40A3",
    x"015DE9E3",
    x"015D9344",
    x"015D3CC8",
    x"015CE66D",
    x"015C9034",
    x"015C3A1C",
    x"015BE426",
    x"015B8E52",
    x"015B389F",
    x"015AE30E",
    x"015A8D9E",
    x"015A384F",
    x"0159E322",
    x"01598E15",
    x"0159392B",
    x"0158E461",
    x"01588FB8",
    x"01583B30",
    x"0157E6CA",
    x"01579284",
    x"01573E5F",
    x"0156EA5B",
    x"01569678",
    x"015642B6",
    x"0155EF14",
    x"01559B93",
    x"01554833",
    x"0154F4F3",
    x"0154A1D3",
    x"01544ED4",
    x"0153FBF6",
    x"0153A937",
    x"01535699",
    x"0153041C",
    x"0152B1BE",
    x"01525F81",
    x"01520D63",
    x"0151BB66",
    x"01516989",
    x"015117CC",
    x"0150C62E",
    x"015074B1",
    x"01502353",
    x"014FD215",
    x"014F80F7",
    x"014F2FF9",
    x"014EDF1A",
    x"014E8E5A",
    x"014E3DBA",
    x"014DED3A",
    x"014D9CD9",
    x"014D4C97",
    x"014CFC75",
    x"014CAC72",
    x"014C5C8E",
    x"014C0CCA",
    x"014BBD24",
    x"014B6D9E",
    x"014B1E37",
    x"014ACEEF",
    x"014A7FC5",
    x"014A30BB",
    x"0149E1CF",
    x"01499302",
    x"01494454",
    x"0148F5C5",
    x"0148A754",
    x"01485902",
    x"01480ACF",
    x"0147BCBA",
    x"01476EC3",
    x"014720EB",
    x"0146D331",
    x"01468596",
    x"01463819",
    x"0145EABA",
    x"01459D7A",
    x"01455057",
    x"01450353",
    x"0144B66D",
    x"014469A4",
    x"01441CFA",
    x"0143D06E",
    x"014383FF",
    x"014337AF",
    x"0142EB7C",
    x"01429F67",
    x"0142536F",
    x"01420795",
    x"0141BBD9",
    x"0141703B",
    x"014124B9",
    x"0140D956",
    x"01408E10",
    x"014042E7",
    x"013FF7DB",
    x"013FACED",
    x"013F621C",
    x"013F1769",
    x"013ECCD2",
    x"013E8259",
    x"013E37FC",
    x"013DEDBD",
    x"013DA39A",
    x"013D5995",
    x"013D0FAC",
    x"013CC5E1",
    x"013C7C32",
    x"013C32A0",
    x"013BE92A",
    x"013B9FD1",
    x"013B5695",
    x"013B0D76",
    x"013AC473",
    x"013A7B8C",
    x"013A32C2",
    x"0139EA15",
    x"0139A183",
    x"0139590E",
    x"013910B6",
    x"0138C879",
    x"01388059",
    x"01383855",
    x"0137F06D",
    x"0137A8A1",
    x"013760F1",
    x"0137195E",
    x"0136D1E6",
    x"01368A8A",
    x"01364349",
    x"0135FC25",
    x"0135B51C",
    x"01356E2F",
    x"0135275E",
    x"0134E0A9",
    x"01349A0F",
    x"01345390",
    x"01340D2D",
    x"0133C6E6",
    x"013380BA",
    x"01333AA9",
    x"0132F4B4",
    x"0132AEDA",
    x"0132691C",
    x"01322378",
    x"0131DDF0",
    x"01319883",
    x"01315331",
    x"01310DFA",
    x"0130C8DE",
    x"013083DD",
    x"01303EF7",
    x"012FFA2C",
    x"012FB57B",
    x"012F70E6",
    x"012F2C6B",
    x"012EE80B",
    x"012EA3C6",
    x"012E5F9B",
    x"012E1B8B",
    x"012DD796",
    x"012D93BB",
    x"012D4FFA",
    x"012D0C54",
    x"012CC8C8",
    x"012C8557",
    x"012C4200",
    x"012BFEC4",
    x"012BBBA1",
    x"012B7899",
    x"012B35AB",
    x"012AF2D7",
    x"012AB01D",
    x"012A6D7D",
    x"012A2AF8",
    x"0129E88C",
    x"0129A63A",
    x"01296402",
    x"012921E4",
    x"0128DFE0",
    x"01289DF5",
    x"01285C24",
    x"01281A6D",
    x"0127D8CF",
    x"0127974C",
    x"012755E1",
    x"01271490",
    x"0126D359",
    x"0126923B",
    x"01265137",
    x"0126104C",
    x"0125CF7A",
    x"01258EC2",
    x"01254E23",
    x"01250D9D",
    x"0124CD30",
    x"01248CDC",
    x"01244CA2",
    x"01240C80",
    x"0123CC78",
    x"01238C89",
    x"01234CB2",
    x"01230CF5",
    x"0122CD50",
    x"01228DC4",
    x"01224E51",
    x"01220EF7",
    x"0121CFB6",
    x"0121908D",
    x"0121517D",
    x"01211285",
    x"0120D3A6",
    x"012094E0",
    x"01205632",
    x"0120179D",
    x"011FD920",
    x"011F9ABB",
    x"011F5C6F",
    x"011F1E3B",
    x"011EE01F",
    x"011EA21C",
    x"011E6430",
    x"011E265D",
    x"011DE8A2",
    x"011DAB00",
    x"011D6D75",
    x"011D3002",
    x"011CF2A7",
    x"011CB564",
    x"011C7839",
    x"011C3B26",
    x"011BFE2B",
    x"011BC148",
    x"011B847C",
    x"011B47C8",
    x"011B0B2C",
    x"011ACEA8",
    x"011A923B",
    x"011A55E5",
    x"011A19A8",
    x"0119DD81",
    x"0119A173",
    x"0119657B",
    x"0119299B",
    x"0118EDD3",
    x"0118B221",
    x"01187687",
    x"01183B05",
    x"0117FF99",
    x"0117C445",
    x"01178908",
    x"01174DE2",
    x"011712D3",
    x"0116D7DB",
    x"01169CFB",
    x"01166231",
    x"0116277E",
    x"0115ECE2",
    x"0115B25D",
    x"011577EE",
    x"01153D97",
    x"01150356",
    x"0114C92C",
    x"01148F19",
    x"0114551D",
    x"01141B37",
    x"0113E167",
    x"0113A7AF",
    x"01136E0C",
    x"01133481",
    x"0112FB0B",
    x"0112C1AC",
    x"01128864",
    x"01124F32",
    x"01121616",
    x"0111DD11",
    x"0111A421",
    x"01116B48",
    x"01113286",
    x"0110F9D9",
    x"0110C142",
    x"011088C2",
    x"01105057",
    x"01101803",
    x"010FDFC5",
    x"010FA79C",
    x"010F6F8A",
    x"010F378D",
    x"010EFFA6",
    x"010EC7D5",
    x"010E901A",
    x"010E5875",
    x"010E20E5",
    x"010DE96B",
    x"010DB207",
    x"010D7AB8",
    x"010D437F",
    x"010D0C5B",
    x"010CD54D",
    x"010C9E55",
    x"010C6771",
    x"010C30A4",
    x"010BF9EB",
    x"010BC348",
    x"010B8CBB",
    x"010B5643",
    x"010B1FDF",
    x"010AE992",
    x"010AB359",
    x"010A7D35",
    x"010A4727",
    x"010A112E",
    x"0109DB4A",
    x"0109A57B",
    x"01096FC0",
    x"01093A1B",
    x"0109048B",
    x"0108CF10",
    x"010899A9",
    x"01086458",
    x"01082F1B",
    x"0107F9F3",
    x"0107C4E0",
    x"01078FE1",
    x"01075AF7",
    x"01072622",
    x"0106F161",
    x"0106BCB5",
    x"0106881E",
    x"0106539B",
    x"01061F2D",
    x"0105EAD3",
    x"0105B68D",
    x"0105825C",
    x"01054E3F",
    x"01051A37",
    x"0104E643",
    x"0104B263",
    x"01047E97",
    x"01044AE0",
    x"0104173D",
    x"0103E3AE",
    x"0103B033",
    x"01037CCC",
    x"01034979",
    x"0103163B",
    x"0102E310",
    x"0102AFF9",
    x"01027CF7",
    x"01024A08",
    x"0102172D",
    x"0101E466",
    x"0101B1B2",
    x"01017F13",
    x"01014C87",
    x"01011A0F",
    x"0100E7AB",
    x"0100B55A",
    x"0100831D",
    x"010050F4",
    x"01001EDE",
    x"00FFD9B7",
    x"00FF75D9",
    x"00FF1223",
    x"00FEAE93",
    x"00FE4B2A",
    x"00FDE7E8",
    x"00FD84CD",
    x"00FD21D9",
    x"00FCBF0B",
    x"00FC5C63",
    x"00FBF9E3",
    x"00FB9788",
    x"00FB3554",
    x"00FAD346",
    x"00FA715F",
    x"00FA0F9E",
    x"00F9AE03",
    x"00F94C8E",
    x"00F8EB3F",
    x"00F88A16",
    x"00F82913",
    x"00F7C836",
    x"00F7677F",
    x"00F706ED",
    x"00F6A681",
    x"00F6463B",
    x"00F5E61A",
    x"00F5861F",
    x"00F5264A",
    x"00F4C699",
    x"00F4670E",
    x"00F407A9",
    x"00F3A868",
    x"00F3494D",
    x"00F2EA57",
    x"00F28B86",
    x"00F22CDA",
    x"00F1CE53",
    x"00F16FF1",
    x"00F111B4",
    x"00F0B39B",
    x"00F055A7",
    x"00EFF7D8",
    x"00EF9A2E",
    x"00EF3CA8",
    x"00EEDF46",
    x"00EE8209",
    x"00EE24F1",
    x"00EDC7FC",
    x"00ED6B2C",
    x"00ED0E81",
    x"00ECB1F9",
    x"00EC5595",
    x"00EBF956",
    x"00EB9D3B",
    x"00EB4143",
    x"00EAE570",
    x"00EA89C0",
    x"00EA2E34",
    x"00E9D2CC",
    x"00E97787",
    x"00E91C66",
    x"00E8C169",
    x"00E8668F",
    x"00E80BD9",
    x"00E7B146",
    x"00E756D6",
    x"00E6FC8A",
    x"00E6A261",
    x"00E6485B",
    x"00E5EE79",
    x"00E594B9",
    x"00E53B1C",
    x"00E4E1A3",
    x"00E4884C",
    x"00E42F18",
    x"00E3D607",
    x"00E37D19",
    x"00E3244E",
    x"00E2CBA5",
    x"00E2731E",
    x"00E21ABB",
    x"00E1C279",
    x"00E16A5B",
    x"00E1125E",
    x"00E0BA84",
    x"00E062CD",
    x"00E00B37",
    x"00DFB3C4",
    x"00DF5C73",
    x"00DF0544",
    x"00DEAE37",
    x"00DE574C",
    x"00DE0082",
    x"00DDA9DB",
    x"00DD5356",
    x"00DCFCF2",
    x"00DCA6B0",
    x"00DC5090",
    x"00DBFA91",
    x"00DBA4B4",
    x"00DB4EF8",
    x"00DAF95E",
    x"00DAA3E6",
    x"00DA4E8E",
    x"00D9F958",
    x"00D9A443",
    x"00D94F50",
    x"00D8FA7D",
    x"00D8A5CC",
    x"00D8513C",
    x"00D7FCCD",
    x"00D7A87E",
    x"00D75451",
    x"00D70044",
    x"00D6AC59",
    x"00D6588E",
    x"00D604E4",
    x"00D5B15A",
    x"00D55DF1",
    x"00D50AA9",
    x"00D4B781",
    x"00D46479",
    x"00D41192",
    x"00D3BECB",
    x"00D36C25",
    x"00D3199F",
    x"00D2C739",
    x"00D274F3",
    x"00D222CE",
    x"00D1D0C8",
    x"00D17EE2",
    x"00D12D1D",
    x"00D0DB77",
    x"00D089F1",
    x"00D0388B",
    x"00CFE745",
    x"00CF961F",
    x"00CF4518",
    x"00CEF431",
    x"00CEA369",
    x"00CE52C1",
    x"00CE0238",
    x"00CDB1CF",
    x"00CD6186",
    x"00CD115B",
    x"00CCC150",
    x"00CC7164",
    x"00CC2197",
    x"00CBD1EA",
    x"00CB825B",
    x"00CB32EC",
    x"00CAE39C",
    x"00CA946A",
    x"00CA4558",
    x"00C9F664",
    x"00C9A78F",
    x"00C958D9",
    x"00C90A42",
    x"00C8BBC9",
    x"00C86D6F",
    x"00C81F33",
    x"00C7D117",
    x"00C78318",
    x"00C73538",
    x"00C6E777",
    x"00C699D3",
    x"00C64C4E",
    x"00C5FEE8",
    x"00C5B19F",
    x"00C56475",
    x"00C51769",
    x"00C4CA7B",
    x"00C47DAA",
    x"00C430F8",
    x"00C3E464",
    x"00C397EE",
    x"00C34B95",
    x"00C2FF5B",
    x"00C2B33E",
    x"00C2673F",
    x"00C21B5D",
    x"00C1CF99",
    x"00C183F3",
    x"00C1386A",
    x"00C0ECFF",
    x"00C0A1B1",
    x"00C05681",
    x"00C00B6E",
    x"00BFC078",
    x"00BF759F",
    x"00BF2AE4",
    x"00BEE046",
    x"00BE95C5",
    x"00BE4B61",
    x"00BE011A",
    x"00BDB6F0",
    x"00BD6CE3",
    x"00BD22F3",
    x"00BCD91F",
    x"00BC8F69",
    x"00BC45CF",
    x"00BBFC52",
    x"00BBB2F2",
    x"00BB69AF",
    x"00BB2088",
    x"00BAD77D",
    x"00BA8E8F",
    x"00BA45BE",
    x"00B9FD09",
    x"00B9B470",
    x"00B96BF4",
    x"00B92394",
    x"00B8DB50",
    x"00B89328",
    x"00B84B1D",
    x"00B8032E",
    x"00B7BB5B",
    x"00B773A3",
    x"00B72C08",
    x"00B6E489",
    x"00B69D26",
    x"00B655DE",
    x"00B60EB3",
    x"00B5C7A3",
    x"00B580AF",
    x"00B539D6",
    x"00B4F319",
    x"00B4AC78",
    x"00B465F3",
    x"00B41F89",
    x"00B3D93A",
    x"00B39307",
    x"00B34CEF",
    x"00B306F3",
    x"00B2C112",
    x"00B27B4C",
    x"00B235A1",
    x"00B1F012",
    x"00B1AA9E",
    x"00B16545",
    x"00B12007",
    x"00B0DAE4",
    x"00B095DC",
    x"00B050EE",
    x"00B00C1C",
    x"00AFC765",
    x"00AF82C9",
    x"00AF3E47",
    x"00AEF9E0",
    x"00AEB594",
    x"00AE7162",
    x"00AE2D4B",
    x"00ADE94F",
    x"00ADA56D",
    x"00AD61A5",
    x"00AD1DF8",
    x"00ACDA66",
    x"00AC96EE",
    x"00AC5390",
    x"00AC104C",
    x"00ABCD23",
    x"00AB8A14",
    x"00AB471F",
    x"00AB0445",
    x"00AAC184",
    x"00AA7EDD",
    x"00AA3C51",
    x"00A9F9DE",
    x"00A9B786",
    x"00A97547",
    x"00A93322",
    x"00A8F117",
    x"00A8AF26",
    x"00A86D4E",
    x"00A82B90",
    x"00A7E9EC",
    x"00A7A861",
    x"00A766F0",
    x"00A72599",
    x"00A6E45B",
    x"00A6A337",
    x"00A6622C",
    x"00A6213A",
    x"00A5E062",
    x"00A59FA3",
    x"00A55EFD",
    x"00A51E70",
    x"00A4DDFD",
    x"00A49DA3",
    x"00A45D62",
    x"00A41D3A",
    x"00A3DD2B",
    x"00A39D35",
    x"00A35D58",
    x"00A31D94",
    x"00A2DDE9",
    x"00A29E57",
    x"00A25EDD",
    x"00A21F7D",
    x"00A1E035",
    x"00A1A106",
    x"00A161EF",
    x"00A122F1",
    x"00A0E40C",
    x"00A0A53F",
    x"00A0668B",
    x"00A027EF",
    x"009FE96B",
    x"009FAB00",
    x"009F6CAE",
    x"009F2E73",
    x"009EF051",
    x"009EB248",
    x"009E7456",
    x"009E367D",
    x"009DF8BC",
    x"009DBB12",
    x"009D7D81",
    x"009D4008",
    x"009D02A7",
    x"009CC55E",
    x"009C882D",
    x"009C4B14",
    x"009C0E12",
    x"009BD129",
    x"009B9457",
    x"009B579D",
    x"009B1AFB",
    x"009ADE70",
    x"009AA1FD",
    x"009A65A1",
    x"009A295D",
    x"0099ED31",
    x"0099B11C",
    x"0099751F",
    x"00993939",
    x"0098FD6A",
    x"0098C1B3",
    x"00988613",
    x"00984A8A",
    x"00980F18",
    x"0097D3BE",
    x"0097987B",
    x"00975D4F",
    x"0097223A",
    x"0096E73C",
    x"0096AC55",
    x"00967185",
    x"009636CD",
    x"0095FC2B",
    x"0095C1A0",
    x"0095872B",
    x"00954CCE",
    x"00951287",
    x"0094D858",
    x"00949E3E",
    x"0094643C",
    x"00942A50",
    x"0093F07B",
    x"0093B6BC",
    x"00937D14",
    x"00934382",
    x"00930A07",
    x"0092D0A3",
    x"00929754",
    x"00925E1C",
    x"009224FB",
    x"0091EBEF",
    x"0091B2FA",
    x"00917A1C",
    x"00914153",
    x"009108A1",
    x"0090D004",
    x"0090977E",
    x"00905F0E",
    x"009026B4",
    x"008FEE70",
    x"008FB641",
    x"008F7E29",
    x"008F4627",
    x"008F0E3A",
    x"008ED664",
    x"008E9EA3",
    x"008E66F8",
    x"008E2F62",
    x"008DF7E3",
    x"008DC079",
    x"008D8924",
    x"008D51E6",
    x"008D1ABC",
    x"008CE3A9",
    x"008CACAB",
    x"008C75C2",
    x"008C3EEF",
    x"008C0831",
    x"008BD188",
    x"008B9AF5",
    x"008B6477",
    x"008B2E0E",
    x"008AF7BB",
    x"008AC17D",
    x"008A8B54",
    x"008A5540",
    x"008A1F41",
    x"0089E958",
    x"0089B383",
    x"00897DC3",
    x"00894819",
    x"00891283",
    x"0088DD02",
    x"0088A796",
    x"0088723F",
    x"00883CFD",
    x"008807D0",
    x"0087D2B7",
    x"00879DB3",
    x"008768C4",
    x"008733E9",
    x"0086FF23",
    x"0086CA72",
    x"008695D5",
    x"0086614D",
    x"00862CD9",
    x"0085F87A",
    x"0085C42F",
    x"00858FF8",
    x"00855BD6",
    x"008527C9",
    x"0084F3CF",
    x"0084BFEA",
    x"00848C19",
    x"0084585D",
    x"008424B4",
    x"0083F120",
    x"0083BDA0",
    x"00838A34",
    x"008356DC",
    x"00832398",
    x"0082F068",
    x"0082BD4C",
    x"00828A44",
    x"00825750",
    x"00822470",
    x"0081F1A4",
    x"0081BEEB",
    x"00818C47",
    x"008159B6",
    x"00812738",
    x"0080F4CF",
    x"0080C279",
    x"00809037",
    x"00805E08",
    x"00802BEE",
    x"007FF9E6",
    x"007FC7F2",
    x"007F9612",
    x"007F6445",
    x"007F328C",
    x"007F00E6",
    x"007ECF53",
    x"007E9DD4",
    x"007E6C68",
    x"007E3B0F",
    x"007E09C9",
    x"007DD897",
    x"007DA778",
    x"007D766C",
    x"007D4574",
    x"007D148E",
    x"007CE3BC",
    x"007CB2FC",
    x"007C8250",
    x"007C51B6",
    x"007C2130",
    x"007BF0BC",
    x"007BC05C",
    x"007B900E",
    x"007B5FD3",
    x"007B2FAB",
    x"007AFF96",
    x"007ACF94",
    x"007A9FA4",
    x"007A6FC7",
    x"007A3FFC",
    x"007A1045",
    x"0079E0A0",
    x"0079B10D",
    x"0079818D",
    x"00795220",
    x"007922C5",
    x"0078F37D",
    x"0078C447",
    x"00789524",
    x"00786613",
    x"00783714",
    x"00780827",
    x"0077D94D",
    x"0077AA86",
    x"00777BD0",
    x"00774D2D",
    x"00771E9C",
    x"0076F01D",
    x"0076C1B0",
    x"00769356",
    x"0076650D",
    x"007636D7",
    x"007608B2",
    x"0075DAA0",
    x"0075ACA0",
    x"00757EB1",
    x"007550D5",
    x"0075230A",
    x"0074F551",
    x"0074C7AA",
    x"00749A15",
    x"00746C92",
    x"00743F20",
    x"007411C1",
    x"0073E472",
    x"0073B736",
    x"00738A0B",
    x"00735CF2",
    x"00732FEB",
    x"007302F5",
    x"0072D610",
    x"0072A93E",
    x"00727C7C",
    x"00724FCC",
    x"0072232E",
    x"0071F6A1",
    x"0071CA25",
    x"00719DBB",
    x"00717162",
    x"0071451A",
    x"007118E4",
    x"0070ECBF",
    x"0070C0AB",
    x"007094A8",
    x"007068B7",
    x"00703CD6",
    x"00701107",
    x"006FE549",
    x"006FB99C",
    x"006F8E00",
    x"006F6275",
    x"006F36FB",
    x"006F0B92",
    x"006EE03A",
    x"006EB4F3",
    x"006E89BD",
    x"006E5E97",
    x"006E3383",
    x"006E087F",
    x"006DDD8C",
    x"006DB2AA",
    x"006D87D9",
    x"006D5D18",
    x"006D3268",
    x"006D07C9",
    x"006CDD3A",
    x"006CB2BC",
    x"006C884E",
    x"006C5DF1",
    x"006C33A5",
    x"006C0969",
    x"006BDF3D",
    x"006BB522",
    x"006B8B18",
    x"006B611E",
    x"006B3734",
    x"006B0D5B",
    x"006AE392",
    x"006AB9D9",
    x"006A9030",
    x"006A6698",
    x"006A3D10",
    x"006A1398",
    x"0069EA31",
    x"0069C0D9",
    x"00699792",
    x"00696E5B",
    x"00694534",
    x"00691C1D",
    x"0068F316",
    x"0068CA1F",
    x"0068A138",
    x"00687861",
    x"00684F9A",
    x"006826E3",
    x"0067FE3C",
    x"0067D5A4",
    x"0067AD1D",
    x"006784A5",
    x"00675C3D",
    x"006733E5",
    x"00670B9D",
    x"0066E364",
    x"0066BB3B",
    x"00669322",
    x"00666B18",
    x"0066431E",
    x"00661B33",
    x"0065F359",
    x"0065CB8D",
    x"0065A3D2",
    x"00657C25",
    x"00655489",
    x"00652CFB",
    x"0065057D",
    x"0064DE0F",
    x"0064B6B0",
    x"00648F60",
    x"00646820",
    x"006440EF",
    x"006419CD",
    x"0063F2BB",
    x"0063CBB8",
    x"0063A4C4",
    x"00637DDF",
    x"00635709",
    x"00633043",
    x"0063098C",
    x"0062E2E3",
    x"0062BC4A",
    x"006295C0",
    x"00626F45",
    x"006248D9",
    x"0062227C",
    x"0061FC2E",
    x"0061D5EF",
    x"0061AFBF",
    x"0061899E",
    x"0061638C",
    x"00613D88",
    x"00611794",
    x"0060F1AE",
    x"0060CBD7",
    x"0060A60F",
    x"00608055",
    x"00605AAA",
    x"0060350E",
    x"00600F81",
    x"005FEA02",
    x"005FC492",
    x"005F9F31",
    x"005F79DE",
    x"005F5499",
    x"005F2F64",
    x"005F0A3C",
    x"005EE524",
    x"005EC019",
    x"005E9B1D",
    x"005E7630",
    x"005E5151",
    x"005E2C81",
    x"005E07BE",
    x"005DE30A",
    x"005DBE65",
    x"005D99CE",
    x"005D7545",
    x"005D50CA",
    x"005D2C5E",
    x"005D07FF",
    x"005CE3AF",
    x"005CBF6E",
    x"005C9B3A",
    x"005C7714",
    x"005C52FD",
    x"005C2EF3",
    x"005C0AF8",
    x"005BE70B",
    x"005BC32C",
    x"005B9F5A",
    x"005B7B97",
    x"005B57E2",
    x"005B343A",
    x"005B10A1",
    x"005AED15",
    x"005AC998",
    x"005AA628",
    x"005A82C6",
    x"005A5F72",
    x"005A3C2B",
    x"005A18F3",
    x"0059F5C8",
    x"0059D2AB",
    x"0059AF9B",
    x"00598C9A",
    x"005969A5",
    x"005946BF",
    x"005923E6",
    x"0059011B",
    x"0058DE5D",
    x"0058BBAD",
    x"0058990B",
    x"00587676",
    x"005853EE",
    x"00583174",
    x"00580F07",
    x"0057ECA8",
    x"0057CA57",
    x"0057A812",
    x"005785DB",
    x"005763B2",
    x"00574195",
    x"00571F86",
    x"0056FD85",
    x"0056DB90",
    x"0056B9A9",
    x"005697CF",
    x"00567603",
    x"00565443",
    x"00563291",
    x"005610EC",
    x"0055EF54",
    x"0055CDC9",
    x"0055AC4B",
    x"00558ADA",
    x"00556976",
    x"00554820",
    x"005526D6",
    x"00550599",
    x"0054E46A",
    x"0054C347",
    x"0054A231",
    x"00548128",
    x"0054602C",
    x"00543F3D",
    x"00541E5B",
    x"0053FD85",
    x"0053DCBD",
    x"0053BC01",
    x"00539B52",
    x"00537AAF",
    x"00535A1A",
    x"00533991",
    x"00531915",
    x"0052F8A5",
    x"0052D843",
    x"0052B7EC",
    x"005297A3",
    x"00527766",
    x"00525736",
    x"00523712",
    x"005216FB",
    x"0051F6F0",
    x"0051D6F2",
    x"0051B700",
    x"0051971B",
    x"00517742",
    x"00515776",
    x"005137B6",
    x"00511802",
    x"0050F85B",
    x"0050D8C0",
    x"0050B931",
    x"005099AF",
    x"00507A39",
    x"00505AD0",
    x"00503B72",
    x"00501C21",
    x"004FFCDC",
    x"004FDDA4",
    x"004FBE77",
    x"004F9F57",
    x"004F8043",
    x"004F613B",
    x"004F423F",
    x"004F234F",
    x"004F046B",
    x"004EE594",
    x"004EC6C8",
    x"004EA808",
    x"004E8955",
    x"004E6AAD",
    x"004E4C11",
    x"004E2D81",
    x"004E0EFE",
    x"004DF086",
    x"004DD21A",
    x"004DB3BA",
    x"004D9565",
    x"004D771D",
    x"004D58E0",
    x"004D3AAF",
    x"004D1C8A",
    x"004CFE71",
    x"004CE064",
    x"004CC262",
    x"004CA46C",
    x"004C8681",
    x"004C68A3",
    x"004C4AD0",
    x"004C2D08",
    x"004C0F4C",
    x"004BF19C",
    x"004BD3F8",
    x"004BB65F",
    x"004B98D1",
    x"004B7B4F",
    x"004B5DD9",
    x"004B406E",
    x"004B230F",
    x"004B05BB",
    x"004AE872",
    x"004ACB35",
    x"004AAE03",
    x"004A90DD",
    x"004A73C2",
    x"004A56B3",
    x"004A39AE",
    x"004A1CB5",
    x"0049FFC8",
    x"0049E2E6",
    x"0049C60F",
    x"0049A943",
    x"00498C82",
    x"00496FCD",
    x"00495323",
    x"00493684",
    x"004919F0",
    x"0048FD68",
    x"0048E0EA",
    x"0048C478",
    x"0048A811",
    x"00488BB5",
    x"00486F64",
    x"0048531E",
    x"004836E3",
    x"00481AB3",
    x"0047FE8E",
    x"0047E274",
    x"0047C665",
    x"0047AA61",
    x"00478E68",
    x"0047727A",
    x"00475697",
    x"00473ABE",
    x"00471EF1",
    x"0047032E",
    x"0046E776",
    x"0046CBC9",
    x"0046B027",
    x"00469490",
    x"00467903",
    x"00465D81",
    x"0046420A",
    x"0046269D",
    x"00460B3C",
    x"0045EFE5",
    x"0045D498",
    x"0045B957",
    x"00459E1F",
    x"004582F3",
    x"004567D1",
    x"00454CBA",
    x"004531AD",
    x"004516AB",
    x"0044FBB3",
    x"0044E0C6",
    x"0044C5E4",
    x"0044AB0C",
    x"0044903E",
    x"0044757B",
    x"00445AC2",
    x"00444014",
    x"00442570",
    x"00440AD7",
    x"0043F048",
    x"0043D5C3",
    x"0043BB49",
    x"0043A0D9",
    x"00438673",
    x"00436C18",
    x"004351C7",
    x"00433780",
    x"00431D43",
    x"00430311",
    x"0042E8E9",
    x"0042CECB",
    x"0042B4B7",
    x"00429AAE",
    x"004280AF",
    x"004266B9",
    x"00424CCE",
    x"004232ED",
    x"00421917",
    x"0041FF4A",
    x"0041E587",
    x"0041CBCE",
    x"0041B220",
    x"0041987B",
    x"00417EE1",
    x"00416550",
    x"00414BCA",
    x"0041324D",
    x"004118DA",
    x"0040FF72",
    x"0040E613",
    x"0040CCBE",
    x"0040B373",
    x"00409A32",
    x"004080FA",
    x"004067CD",
    x"00404EA9",
    x"0040358F",
    x"00401C7F",
    x"00400379",
    x"003FEA7D",
    x"003FD18A",
    x"003FB8A1",
    x"003F9FC2",
    x"003F86EC",
    x"003F6E20",
    x"003F555E",
    x"003F3CA6",
    x"003F23F7",
    x"003F0B51",
    x"003EF2B6",
    x"003EDA24",
    x"003EC19B",
    x"003EA91D",
    x"003E90A7",
    x"003E783C",
    x"003E5FD9",
    x"003E4781",
    x"003E2F31",
    x"003E16EC",
    x"003DFEB0",
    x"003DE67D",
    x"003DCE53",
    x"003DB634",
    x"003D9E1D",
    x"003D8610",
    x"003D6E0C",
    x"003D5612",
    x"003D3E21",
    x"003D263A",
    x"003D0E5B",
    x"003CF686",
    x"003CDEBB",
    x"003CC6F8",
    x"003CAF3F",
    x"003C978F",
    x"003C7FE9",
    x"003C684B",
    x"003C50B7",
    x"003C392C",
    x"003C21AB",
    x"003C0A32",
    x"003BF2C3",
    x"003BDB5C",
    x"003BC3FF",
    x"003BACAB",
    x"003B9560",
    x"003B7E1F",
    x"003B66E6",
    x"003B4FB6",
    x"003B3890",
    x"003B2172",
    x"003B0A5D",
    x"003AF352",
    x"003ADC4F",
    x"003AC556",
    x"003AAE65",
    x"003A977E",
    x"003A809F",
    x"003A69C9",
    x"003A52FC",
    x"003A3C38",
    x"003A257D",
    x"003A0ECB",
    x"0039F822",
    x"0039E181",
    x"0039CAE9",
    x"0039B45B",
    x"00399DD4",
    x"00398757",
    x"003970E3",
    x"00395A77",
    x"00394414",
    x"00392DBA",
    x"00391768",
    x"00390120",
    x"0038EADF",
    x"0038D4A8",
    x"0038BE79",
    x"0038A853",
    x"00389236",
    x"00387C21",
    x"00386615",
    x"00385011",
    x"00383A16",
    x"00382424",
    x"00380E3A",
    x"0037F859",
    x"0037E280",
    x"0037CCB0",
    x"0037B6E8",
    x"0037A129",
    x"00378B72",
    x"003775C4",
    x"0037601E",
    x"00374A81",
    x"003734EC",
    x"00371F5F",
    x"003709DB",
    x"0036F460",
    x"0036DEED",
    x"0036C982",
    x"0036B41F",
    x"00369EC5",
    x"00368973",
    x"0036742A",
    x"00365EE8",
    x"003649AF",
    x"0036347F",
    x"00361F56",
    x"00360A36",
    x"0035F51E",
    x"0035E00F",
    x"0035CB07",
    x"0035B608",
    x"0035A111",
    x"00358C22",
    x"0035773C",
    x"0035625D",
    x"00354D87",
    x"003538B9",
    x"003523F2",
    x"00350F34",
    x"0034FA7F",
    x"0034E5D1",
    x"0034D12B",
    x"0034BC8D",
    x"0034A7F8",
    x"0034936A",
    x"00347EE5",
    x"00346A67",
    x"003455F1",
    x"00344184",
    x"00342D1E",
    x"003418C1",
    x"0034046B",
    x"0033F01D",
    x"0033DBD7",
    x"0033C799",
    x"0033B363",
    x"00339F35",
    x"00338B0F",
    x"003376F1",
    x"003362DA",
    x"00334ECB",
    x"00333AC4",
    x"003326C5",
    x"003312CE",
    x"0032FEDF",
    x"0032EAF7",
    x"0032D717",
    x"0032C33F",
    x"0032AF6F",
    x"00329BA6",
    x"003287E5",
    x"0032742C",
    x"0032607A",
    x"00324CD0",
    x"0032392E",
    x"00322594",
    x"00321201",
    x"0031FE76",
    x"0031EAF2",
    x"0031D776",
    x"0031C402",
    x"0031B095",
    x"00319D30",
    x"003189D2",
    x"0031767C",
    x"0031632E",
    x"00314FE7",
    x"00313CA7",
    x"0031296F",
    x"0031163F",
    x"00310316",
    x"0030EFF4",
    x"0030DCDA",
    x"0030C9C8",
    x"0030B6BD",
    x"0030A3B9",
    x"003090BD",
    x"00307DC8",
    x"00306ADB",
    x"003057F4",
    x"00304516",
    x"0030323F",
    x"00301F6F",
    x"00300CA6",
    x"002FF9E5",
    x"002FE72B",
    x"002FD478",
    x"002FC1CD",
    x"002FAF29",
    x"002F9C8C",
    x"002F89F6",
    x"002F7768",
    x"002F64E1",
    x"002F5261",
    x"002F3FE9",
    x"002F2D77",
    x"002F1B0D",
    x"002F08AA",
    x"002EF64E",
    x"002EE3FA",
    x"002ED1AC",
    x"002EBF66",
    x"002EAD27",
    x"002E9AEF",
    x"002E88BE",
    x"002E7694",
    x"002E6471",
    x"002E5255",
    x"002E4041",
    x"002E2E33",
    x"002E1C2D",
    x"002E0A2D",
    x"002DF835",
    x"002DE643",
    x"002DD459",
    x"002DC275",
    x"002DB099",
    x"002D9EC3",
    x"002D8CF5",
    x"002D7B2D",
    x"002D696D",
    x"002D57B3",
    x"002D4600",
    x"002D3454",
    x"002D22AF",
    x"002D1111",
    x"002CFF7A",
    x"002CEDEA",
    x"002CDC60",
    x"002CCADD",
    x"002CB962",
    x"002CA7ED",
    x"002C967E",
    x"002C8517",
    x"002C73B6",
    x"002C625D",
    x"002C5109",
    x"002C3FBD",
    x"002C2E78",
    x"002C1D39",
    x"002C0C01",
    x"002BFAD0",
    x"002BE9A5",
    x"002BD881",
    x"002BC764",
    x"002BB64D",
    x"002BA53D",
    x"002B9434",
    x"002B8332",
    x"002B7236",
    x"002B6140",
    x"002B5052",
    x"002B3F6A",
    x"002B2E88",
    x"002B1DAD",
    x"002B0CD9",
    x"002AFC0B",
    x"002AEB44",
    x"002ADA83",
    x"002AC9C9",
    x"002AB916",
    x"002AA869",
    x"002A97C2",
    x"002A8722",
    x"002A7689",
    x"002A65F5",
    x"002A5569",
    x"002A44E3",
    x"002A3463",
    x"002A23EA",
    x"002A1377",
    x"002A030B",
    x"0029F2A5",
    x"0029E245",
    x"0029D1EC",
    x"0029C199",
    x"0029B14D",
    x"0029A107",
    x"002990C7",
    x"0029808D",
    x"0029705A",
    x"0029602E",
    x"00295007",
    x"00293FE7",
    x"00292FCD",
    x"00291FBA",
    x"00290FAD",
    x"0028FFA6",
    x"0028EFA5",
    x"0028DFAA",
    x"0028CFB6",
    x"0028BFC8",
    x"0028AFE0",
    x"00289FFF",
    x"00289023",
    x"0028804E",
    x"0028707F",
    x"002860B6",
    x"002850F3",
    x"00284137",
    x"00283180",
    x"002821D0",
    x"00281226",
    x"00280282",
    x"0027F2E4",
    x"0027E34C",
    x"0027D3BB",
    x"0027C42F",
    x"0027B4A9",
    x"0027A52A",
    x"002795B0",
    x"0027863D",
    x"002776CF",
    x"00276768",
    x"00275807",
    x"002748AB",
    x"00273956",
    x"00272A06",
    x"00271ABD",
    x"00270B79",
    x"0026FC3C",
    x"0026ED04",
    x"0026DDD3",
    x"0026CEA7",
    x"0026BF81",
    x"0026B061",
    x"0026A148",
    x"00269233",
    x"00268325",
    x"0026741D",
    x"0026651B",
    x"0026561E",
    x"00264727",
    x"00263836",
    x"0026294B",
    x"00261A66",
    x"00260B87",
    x"0025FCAD",
    x"0025EDD9",
    x"0025DF0B",
    x"0025D043",
    x"0025C181",
    x"0025B2C4",
    x"0025A40D",
    x"0025955C",
    x"002586B0",
    x"0025780B",
    x"0025696A",
    x"00255AD0",
    x"00254C3C",
    x"00253DAD",
    x"00252F23",
    x"002520A0",
    x"00251222",
    x"002503AA",
    x"0024F537",
    x"0024E6CA",
    x"0024D863",
    x"0024CA01",
    x"0024BBA5",
    x"0024AD4E",
    x"00249EFD",
    x"002490B2",
    x"0024826C",
    x"0024742C",
    x"002465F2",
    x"002457BD",
    x"0024498D",
    x"00243B63",
    x"00242D3F",
    x"00241F20",
    x"00241106",
    x"002402F3",
    x"0023F4E4",
    x"0023E6DB",
    x"0023D8D8",
    x"0023CADA",
    x"0023BCE1",
    x"0023AEEE",
    x"0023A101",
    x"00239318",
    x"00238536",
    x"00237758",
    x"00236980",
    x"00235BAE",
    x"00234DE1",
    x"00234019",
    x"00233257",
    x"0023249A",
    x"002316E2",
    x"00230930",
    x"0022FB83",
    x"0022EDDB",
    x"0022E039",
    x"0022D29C",
    x"0022C505",
    x"0022B772",
    x"0022A9E5",
    x"00229C5E",
    x"00228EDB",
    x"0022815E",
    x"002273E6",
    x"00226673",
    x"00225906",
    x"00224B9E",
    x"00223E3B",
    x"002230DD",
    x"00222385",
    x"00221631",
    x"002208E3",
    x"0021FB9B",
    x"0021EE57",
    x"0021E118",
    x"0021D3DF",
    x"0021C6AB",
    x"0021B97C",
    x"0021AC52",
    x"00219F2D",
    x"0021920E",
    x"002184F3",
    x"002177DE",
    x"00216ACD",
    x"00215DC2",
    x"002150BC",
    x"002143BB",
    x"002136BF",
    x"002129C8",
    x"00211CD7",
    x"00210FEA",
    x"00210302",
    x"0020F61F",
    x"0020E942",
    x"0020DC69",
    x"0020CF96",
    x"0020C2C7",
    x"0020B5FD",
    x"0020A939",
    x"00209C79",
    x"00208FBF",
    x"00208309",
    x"00207658",
    x"002069AC",
    x"00205D06",
    x"00205064",
    x"002043C7",
    x"0020372F",
    x"00202A9C",
    x"00201E0E",
    x"00201184",
    x"00200500",
    x"001FF880",
    x"001FEC06",
    x"001FDF90",
    x"001FD31F",
    x"001FC6B3",
    x"001FBA4C",
    x"001FADE9",
    x"001FA18C",
    x"001F9533",
    x"001F88DF",
    x"001F7C90",
    x"001F7046",
    x"001F6401",
    x"001F57C0",
    x"001F4B84",
    x"001F3F4D",
    x"001F331B",
    x"001F26ED",
    x"001F1AC4",
    x"001F0EA0",
    x"001F0281",
    x"001EF666",
    x"001EEA50",
    x"001EDE3F",
    x"001ED233",
    x"001EC62B",
    x"001EBA28",
    x"001EAE29",
    x"001EA230",
    x"001E963B",
    x"001E8A4A",
    x"001E7E5F",
    x"001E7278",
    x"001E6695",
    x"001E5AB8",
    x"001E4EDE",
    x"001E430A",
    x"001E373A",
    x"001E2B6F",
    x"001E1FA8",
    x"001E13E6",
    x"001E0829",
    x"001DFC70",
    x"001DF0BB",
    x"001DE50C",
    x"001DD960",
    x"001DCDBA",
    x"001DC218",
    x"001DB67A",
    x"001DAAE1",
    x"001D9F4D",
    x"001D93BD",
    x"001D8831",
    x"001D7CAA",
    x"001D7128",
    x"001D65AA",
    x"001D5A30",
    x"001D4EBB",
    x"001D434B",
    x"001D37DF",
    x"001D2C77",
    x"001D2114",
    x"001D15B5",
    x"001D0A5B",
    x"001CFF05",
    x"001CF3B4",
    x"001CE867",
    x"001CDD1E",
    x"001CD1DA",
    x"001CC69A",
    x"001CBB5F",
    x"001CB028",
    x"001CA4F5",
    x"001C99C7",
    x"001C8E9D",
    x"001C8378",
    x"001C7856",
    x"001C6D3A",
    x"001C6221",
    x"001C570D",
    x"001C4BFD",
    x"001C40F2",
    x"001C35EA",
    x"001C2AE7",
    x"001C1FE9",
    x"001C14EF",
    x"001C09F8",
    x"001BFF07",
    x"001BF419",
    x"001BE930",
    x"001BDE4B",
    x"001BD36A",
    x"001BC88E",
    x"001BBDB6",
    x"001BB2E2",
    x"001BA812",
    x"001B9D46",
    x"001B927F",
    x"001B87BC",
    x"001B7CFD",
    x"001B7242",
    x"001B678C",
    x"001B5CD9",
    x"001B522B",
    x"001B4781",
    x"001B3CDB",
    x"001B323A",
    x"001B279C",
    x"001B1D03",
    x"001B126D",
    x"001B07DC",
    x"001AFD4F",
    x"001AF2C6",
    x"001AE842",
    x"001ADDC1",
    x"001AD344",
    x"001AC8CC",
    x"001ABE57",
    x"001AB3E7",
    x"001AA97B",
    x"001A9F13",
    x"001A94AF",
    x"001A8A4F",
    x"001A7FF3",
    x"001A759B",
    x"001A6B47",
    x"001A60F7",
    x"001A56AB",
    x"001A4C63",
    x"001A421F",
    x"001A37DF",
    x"001A2DA4",
    x"001A236C",
    x"001A1938",
    x"001A0F08",
    x"001A04DC",
    x"0019FAB4",
    x"0019F090",
    x"0019E670",
    x"0019DC54",
    x"0019D23C",
    x"0019C828",
    x"0019BE18",
    x"0019B40C",
    x"0019AA03",
    x"00199FFF",
    x"001995FE",
    x"00198C02",
    x"00198209",
    x"00197814",
    x"00196E23",
    x"00196436",
    x"00195A4D",
    x"00195067",
    x"00194686",
    x"00193CA8",
    x"001932CF",
    x"001928F9",
    x"00191F26",
    x"00191558",
    x"00190B8E",
    x"001901C7",
    x"0018F804",
    x"0018EE45",
    x"0018E48A",
    x"0018DAD3",
    x"0018D11F",
    x"0018C770",
    x"0018BDC4",
    x"0018B41B",
    x"0018AA77",
    x"0018A0D6",
    x"00189739",
    x"00188DA0",
    x"0018840A",
    x"00187A79",
    x"001870EB",
    x"00186761",
    x"00185DDA",
    x"00185457",
    x"00184AD8",
    x"0018415D",
    x"001837E5",
    x"00182E71",
    x"00182501",
    x"00181B94",
    x"0018122B",
    x"001808C6",
    x"0017FF64",
    x"0017F606",
    x"0017ECAC",
    x"0017E356",
    x"0017DA03",
    x"0017D0B3",
    x"0017C768",
    x"0017BE1F",
    x"0017B4DB",
    x"0017AB9A",
    x"0017A25D",
    x"00179923",
    x"00178FED",
    x"001786BB",
    x"00177D8C",
    x"00177461",
    x"00176B39",
    x"00176215",
    x"001758F4",
    x"00174FD8",
    x"001746BE",
    x"00173DA8",
    x"00173496",
    x"00172B87",
    x"0017227C",
    x"00171974",
    x"00171070",
    x"0017076F",
    x"0016FE72",
    x"0016F579",
    x"0016EC82",
    x"0016E390",
    x"0016DAA1",
    x"0016D1B5",
    x"0016C8CD",
    x"0016BFE8",
    x"0016B707",
    x"0016AE29",
    x"0016A54F",
    x"00169C78",
    x"001693A5",
    x"00168AD5",
    x"00168208",
    x"0016793F",
    x"00167079",
    x"001667B7",
    x"00165EF8",
    x"0016563D",
    x"00164D85",
    x"001644D0",
    x"00163C1F",
    x"00163371",
    x"00162AC7",
    x"00162220",
    x"0016197C",
    x"001610DC",
    x"0016083F",
    x"0015FFA6",
    x"0015F70F",
    x"0015EE7D",
    x"0015E5ED",
    x"0015DD61",
    x"0015D4D8",
    x"0015CC53",
    x"0015C3D1",
    x"0015BB52",
    x"0015B2D6",
    x"0015AA5E",
    x"0015A1E9",
    x"00159978",
    x"00159109",
    x"0015889E",
    x"00158037",
    x"001577D2",
    x"00156F71",
    x"00156713",
    x"00155EB8",
    x"00155661",
    x"00154E0D",
    x"001545BC",
    x"00153D6E",
    x"00153524",
    x"00152CDD",
    x"00152499",
    x"00151C58",
    x"0015141B",
    x"00150BE1",
    x"001503AA",
    x"0014FB76",
    x"0014F345",
    x"0014EB18",
    x"0014E2ED",
    x"0014DAC6",
    x"0014D2A3",
    x"0014CA82",
    x"0014C264",
    x"0014BA4A",
    x"0014B233",
    x"0014AA1F",
    x"0014A20E",
    x"00149A00",
    x"001491F6",
    x"001489EE",
    x"001481EA",
    x"001479E9",
    x"001471EB",
    x"001469F0",
    x"001461F8",
    x"00145A03",
    x"00145211",
    x"00144A23",
    x"00144238",
    x"00143A4F",
    x"0014326A",
    x"00142A88",
    x"001422A9",
    x"00141ACD",
    x"001412F4",
    x"00140B1E",
    x"0014034B",
    x"0013FB7B",
    x"0013F3AF",
    x"0013EBE5",
    x"0013E41E",
    x"0013DC5B",
    x"0013D49A",
    x"0013CCDD",
    x"0013C522",
    x"0013BD6B",
    x"0013B5B6",
    x"0013AE05",
    x"0013A656",
    x"00139EAB",
    x"00139702",
    x"00138F5D",
    x"001387BA",
    x"0013801B",
    x"0013787E",
    x"001370E5",
    x"0013694E",
    x"001361BA",
    x"00135A2A",
    x"0013529C",
    x"00134B11",
    x"00134389",
    x"00133C04",
    x"00133482",
    x"00132D03",
    x"00132587",
    x"00131E0E",
    x"00131698",
    x"00130F24",
    x"001307B4",
    x"00130046",
    x"0012F8DC",
    x"0012F174",
    x"0012EA0F",
    x"0012E2AD",
    x"0012DB4E",
    x"0012D3F2",
    x"0012CC98",
    x"0012C542",
    x"0012BDEE",
    x"0012B69D",
    x"0012AF50",
    x"0012A804",
    x"0012A0BC",
    x"00129977",
    x"00129234",
    x"00128AF5",
    x"001283B8",
    x"00127C7E",
    x"00127547",
    x"00126E12",
    x"001266E1",
    x"00125FB2",
    x"00125886",
    x"0012515D",
    x"00124A36",
    x"00124313",
    x"00123BF2",
    x"001234D4",
    x"00122DB9",
    x"001226A0",
    x"00121F8A",
    x"00121877",
    x"00121167",
    x"00120A5A",
    x"0012034F",
    x"0011FC47",
    x"0011F542",
    x"0011EE40",
    x"0011E740",
    x"0011E043",
    x"0011D949",
    x"0011D251",
    x"0011CB5C",
    x"0011C46A",
    x"0011BD7B",
    x"0011B68E",
    x"0011AFA4",
    x"0011A8BD",
    x"0011A1D9",
    x"00119AF7",
    x"00119417",
    x"00118D3B",
    x"00118661",
    x"00117F8A",
    x"001178B5",
    x"001171E4",
    x"00116B15",
    x"00116448",
    x"00115D7E",
    x"001156B7",
    x"00114FF2",
    x"00114931",
    x"00114271",
    x"00113BB5",
    x"001134FB",
    x"00112E43",
    x"0011278E",
    x"001120DC",
    x"00111A2D",
    x"00111380",
    x"00110CD6",
    x"0011062E",
    x"0010FF89",
    x"0010F8E6",
    x"0010F246",
    x"0010EBA9",
    x"0010E50E",
    x"0010DE76",
    x"0010D7E0",
    x"0010D14D",
    x"0010CABD",
    x"0010C42F",
    x"0010BDA4",
    x"0010B71B",
    x"0010B095",
    x"0010AA11",
    x"0010A390",
    x"00109D11",
    x"00109695",
    x"0010901B",
    x"001089A4",
    x"00108330",
    x"00107CBE",
    x"0010764E",
    x"00106FE1",
    x"00106977",
    x"0010630F",
    x"00105CAA",
    x"00105647",
    x"00104FE6",
    x"00104988",
    x"0010432D",
    x"00103CD4",
    x"0010367D",
    x"00103029",
    x"001029D8",
    x"00102388",
    x"00101D3C",
    x"001016F2",
    x"001010AA",
    x"00100A65",
    x"00100422",
    x"000FFDE1",
    x"000FF7A3",
    x"000FF168",
    x"000FEB2F",
    x"000FE4F8",
    x"000FDEC4",
    x"000FD892",
    x"000FD263",
    x"000FCC36",
    x"000FC60B",
    x"000FBFE3",
    x"000FB9BD",
    x"000FB39A",
    x"000FAD79",
    x"000FA75A",
    x"000FA13E",
    x"000F9B24",
    x"000F950D",
    x"000F8EF8",
    x"000F88E5",
    x"000F82D5",
    x"000F7CC7",
    x"000F76BC",
    x"000F70B2",
    x"000F6AAC",
    x"000F64A7",
    x"000F5EA5",
    x"000F58A5",
    x"000F52A8",
    x"000F4CAD",
    x"000F46B4",
    x"000F40BD",
    x"000F3AC9",
    x"000F34D7",
    x"000F2EE8",
    x"000F28FB",
    x"000F2310",
    x"000F1D27",
    x"000F1741",
    x"000F115D",
    x"000F0B7B",
    x"000F059C",
    x"000EFFBF",
    x"000EF9E4",
    x"000EF40C",
    x"000EEE36",
    x"000EE862",
    x"000EE290",
    x"000EDCC1",
    x"000ED6F4",
    x"000ED129",
    x"000ECB60",
    x"000EC59A",
    x"000EBFD6",
    x"000EBA14",
    x"000EB455",
    x"000EAE97",
    x"000EA8DC",
    x"000EA323",
    x"000E9D6D",
    x"000E97B8",
    x"000E9206",
    x"000E8C56",
    x"000E86A8",
    x"000E80FD",
    x"000E7B54",
    x"000E75AD",
    x"000E7008",
    x"000E6A65",
    x"000E64C5",
    x"000E5F26",
    x"000E598A",
    x"000E53F0",
    x"000E4E59",
    x"000E48C3",
    x"000E4330",
    x"000E3D9F",
    x"000E3810",
    x"000E3283",
    x"000E2CF8",
    x"000E2770",
    x"000E21E9",
    x"000E1C65",
    x"000E16E3",
    x"000E1163",
    x"000E0BE6",
    x"000E066A",
    x"000E00F1",
    x"000DFB79",
    x"000DF604",
    x"000DF091",
    x"000DEB20",
    x"000DE5B2",
    x"000DE045",
    x"000DDADA",
    x"000DD572",
    x"000DD00C",
    x"000DCAA7",
    x"000DC545",
    x"000DBFE5",
    x"000DBA87",
    x"000DB52B",
    x"000DAFD2",
    x"000DAA7A",
    x"000DA525",
    x"000D9FD1",
    x"000D9A80",
    x"000D9530",
    x"000D8FE3",
    x"000D8A98",
    x"000D854F",
    x"000D8008",
    x"000D7AC3",
    x"000D7580",
    x"000D703F",
    x"000D6B00",
    x"000D65C3",
    x"000D6089",
    x"000D5B50",
    x"000D5619",
    x"000D50E5",
    x"000D4BB2",
    x"000D4682",
    x"000D4153",
    x"000D3C27",
    x"000D36FC",
    x"000D31D4",
    x"000D2CAD",
    x"000D2789",
    x"000D2266",
    x"000D1D46",
    x"000D1827",
    x"000D130B",
    x"000D0DF1",
    x"000D08D8",
    x"000D03C2",
    x"000CFEAD",
    x"000CF99B",
    x"000CF48A",
    x"000CEF7C",
    x"000CEA6F",
    x"000CE564",
    x"000CE05C",
    x"000CDB55",
    x"000CD651",
    x"000CD14E",
    x"000CCC4D",
    x"000CC74E",
    x"000CC251",
    x"000CBD56",
    x"000CB85D",
    x"000CB366",
    x"000CAE71",
    x"000CA97E",
    x"000CA48D",
    x"000C9F9D",
    x"000C9AB0",
    x"000C95C5",
    x"000C90DB",
    x"000C8BF3",
    x"000C870E",
    x"000C822A",
    x"000C7D48",
    x"000C7868",
    x"000C738A",
    x"000C6EAE",
    x"000C69D4",
    x"000C64FB",
    x"000C6025",
    x"000C5B50",
    x"000C567D",
    x"000C51AC",
    x"000C4CDD",
    x"000C4810",
    x"000C4345",
    x"000C3E7C",
    x"000C39B4",
    x"000C34EF",
    x"000C302B",
    x"000C2B69",
    x"000C26A9",
    x"000C21EB",
    x"000C1D2F",
    x"000C1874",
    x"000C13BB",
    x"000C0F05",
    x"000C0A50",
    x"000C059D",
    x"000C00EB",
    x"000BFC3C",
    x"000BF78E",
    x"000BF2E3",
    x"000BEE39",
    x"000BE990",
    x"000BE4EA",
    x"000BE046",
    x"000BDBA3",
    x"000BD702",
    x"000BD263",
    x"000BCDC6",
    x"000BC92A",
    x"000BC490",
    x"000BBFF9",
    x"000BBB62",
    x"000BB6CE",
    x"000BB23C",
    x"000BADAB",
    x"000BA91C",
    x"000BA48F",
    x"000BA003",
    x"000B9B7A",
    x"000B96F2",
    x"000B926C",
    x"000B8DE8",
    x"000B8965",
    x"000B84E4",
    x"000B8065",
    x"000B7BE8",
    x"000B776C",
    x"000B72F3",
    x"000B6E7B",
    x"000B6A04",
    x"000B6590",
    x"000B611D",
    x"000B5CAC",
    x"000B583D",
    x"000B53CF",
    x"000B4F63",
    x"000B4AF9",
    x"000B4690",
    x"000B422A",
    x"000B3DC5",
    x"000B3962",
    x"000B3500",
    x"000B30A0",
    x"000B2C42",
    x"000B27E6",
    x"000B238B",
    x"000B1F32",
    x"000B1ADA",
    x"000B1685",
    x"000B1231",
    x"000B0DDF",
    x"000B098E",
    x"000B053F",
    x"000B00F2",
    x"000AFCA6",
    x"000AF85D",
    x"000AF414",
    x"000AEFCE",
    x"000AEB89",
    x"000AE746",
    x"000AE304",
    x"000ADEC4",
    x"000ADA86",
    x"000AD64A",
    x"000AD20F",
    x"000ACDD6",
    x"000AC99E",
    x"000AC568",
    x"000AC134",
    x"000ABD01",
    x"000AB8D0",
    x"000AB4A1",
    x"000AB073",
    x"000AAC47",
    x"000AA81C",
    x"000AA3F4",
    x"000A9FCC",
    x"000A9BA7",
    x"000A9783",
    x"000A9360",
    x"000A8F40",
    x"000A8B20",
    x"000A8703",
    x"000A82E7",
    x"000A7ECD",
    x"000A7AB4",
    x"000A769D",
    x"000A7287",
    x"000A6E73",
    x"000A6A61",
    x"000A6650",
    x"000A6241",
    x"000A5E33",
    x"000A5A27",
    x"000A561D",
    x"000A5214",
    x"000A4E0D",
    x"000A4A07",
    x"000A4603",
    x"000A4200",
    x"000A3DFF",
    x"000A3A00",
    x"000A3602",
    x"000A3206",
    x"000A2E0B",
    x"000A2A12",
    x"000A261A",
    x"000A2224",
    x"000A1E30",
    x"000A1A3D",
    x"000A164B",
    x"000A125B",
    x"000A0E6D",
    x"000A0A80",
    x"000A0695",
    x"000A02AB",
    x"0009FEC2",
    x"0009FADC",
    x"0009F6F6",
    x"0009F313",
    x"0009EF31",
    x"0009EB50",
    x"0009E771",
    x"0009E393",
    x"0009DFB7",
    x"0009DBDC",
    x"0009D803",
    x"0009D42C",
    x"0009D055",
    x"0009CC81",
    x"0009C8AE",
    x"0009C4DC",
    x"0009C10C",
    x"0009BD3D",
    x"0009B970",
    x"0009B5A4",
    x"0009B1DA",
    x"0009AE11",
    x"0009AA4A",
    x"0009A684",
    x"0009A2C0",
    x"00099EFD",
    x"00099B3C",
    x"0009977C",
    x"000993BD",
    x"00099000",
    x"00098C45",
    x"0009888B",
    x"000984D2",
    x"0009811B",
    x"00097D65",
    x"000979B1",
    x"000975FE",
    x"0009724D",
    x"00096E9D",
    x"00096AEF",
    x"00096741",
    x"00096396",
    x"00095FEC",
    x"00095C43",
    x"0009589C",
    x"000954F6",
    x"00095151",
    x"00094DAE",
    x"00094A0D",
    x"0009466C",
    x"000942CE",
    x"00093F30",
    x"00093B94",
    x"000937FA",
    x"00093460",
    x"000930C9",
    x"00092D32",
    x"0009299D",
    x"0009260A",
    x"00092278",
    x"00091EE7",
    x"00091B57",
    x"000917CA",
    x"0009143D",
    x"000910B2",
    x"00090D28",
    x"0009099F",
    x"00090618",
    x"00090293",
    x"0008FF0E",
    x"0008FB8B",
    x"0008F80A",
    x"0008F48A",
    x"0008F10B",
    x"0008ED8D",
    x"0008EA11",
    x"0008E696",
    x"0008E31D",
    x"0008DFA5",
    x"0008DC2E",
    x"0008D8B9",
    x"0008D545",
    x"0008D1D2",
    x"0008CE61",
    x"0008CAF1",
    x"0008C783",
    x"0008C415",
    x"0008C0A9",
    x"0008BD3F",
    x"0008B9D5",
    x"0008B66E",
    x"0008B307",
    x"0008AFA2",
    x"0008AC3E",
    x"0008A8DB",
    x"0008A57A",
    x"0008A21A",
    x"00089EBB",
    x"00089B5E",
    x"00089802",
    x"000894A7",
    x"0008914E",
    x"00088DF6",
    x"00088A9F",
    x"00088749",
    x"000883F5",
    x"000880A2",
    x"00087D51",
    x"00087A00",
    x"000876B1",
    x"00087364",
    x"00087017",
    x"00086CCC",
    x"00086982",
    x"0008663A",
    x"000862F2",
    x"00085FAC",
    x"00085C68",
    x"00085924",
    x"000855E2",
    x"000852A1",
    x"00084F61",
    x"00084C23",
    x"000848E6",
    x"000845AA",
    x"0008426F",
    x"00083F36",
    x"00083BFE",
    x"000838C7",
    x"00083592",
    x"0008325D",
    x"00082F2A",
    x"00082BF9",
    x"000828C8",
    x"00082599",
    x"0008226B",
    x"00081F3E",
    x"00081C12",
    x"000818E8",
    x"000815BF",
    x"00081297",
    x"00080F70",
    x"00080C4B",
    x"00080927",
    x"00080604",
    x"000802E2",
    x"0007FFC1",
    x"0007FCA2",
    x"0007F984",
    x"0007F667",
    x"0007F34C",
    x"0007F031",
    x"0007ED18",
    x"0007EA00",
    x"0007E6E9",
    x"0007E3D3",
    x"0007E0BF",
    x"0007DDAC",
    x"0007DA9A",
    x"0007D789",
    x"0007D479",
    x"0007D16B",
    x"0007CE5E",
    x"0007CB52",
    x"0007C847",
    x"0007C53D",
    x"0007C235",
    x"0007BF2E",
    x"0007BC28",
    x"0007B923",
    x"0007B61F",
    x"0007B31C",
    x"0007B01B",
    x"0007AD1B",
    x"0007AA1C",
    x"0007A71E",
    x"0007A421",
    x"0007A126",
    x"00079E2B",
    x"00079B32",
    x"0007983A",
    x"00079543",
    x"0007924D",
    x"00078F59",
    x"00078C65",
    x"00078973",
    x"00078682",
    x"00078392",
    x"000780A3",
    x"00077DB6",
    x"00077AC9",
    x"000777DE",
    x"000774F3",
    x"0007720A",
    x"00076F22",
    x"00076C3B",
    x"00076956",
    x"00076671",
    x"0007638E",
    x"000760AB",
    x"00075DCA",
    x"00075AEA",
    x"0007580B",
    x"0007552D",
    x"00075251",
    x"00074F75",
    x"00074C9B",
    x"000749C1",
    x"000746E9",
    x"00074412",
    x"0007413C",
    x"00073E67",
    x"00073B93",
    x"000738C0",
    x"000735EF",
    x"0007331E",
    x"0007304F",
    x"00072D80",
    x"00072AB3",
    x"000727E7",
    x"0007251C",
    x"00072252",
    x"00071F89",
    x"00071CC1",
    x"000719FB",
    x"00071735",
    x"00071471",
    x"000711AD",
    x"00070EEB",
    x"00070C2A",
    x"00070969",
    x"000706AA",
    x"000703EC",
    x"0007012F",
    x"0006FE73",
    x"0006FBB8",
    x"0006F8FF",
    x"0006F646",
    x"0006F38E",
    x"0006F0D7",
    x"0006EE22",
    x"0006EB6D",
    x"0006E8BA",
    x"0006E608",
    x"0006E356",
    x"0006E0A6",
    x"0006DDF7",
    x"0006DB49",
    x"0006D89B",
    x"0006D5EF",
    x"0006D344",
    x"0006D09A",
    x"0006CDF1",
    x"0006CB49",
    x"0006C8A3",
    x"0006C5FD",
    x"0006C358",
    x"0006C0B4",
    x"0006BE11",
    x"0006BB70",
    x"0006B8CF",
    x"0006B62F",
    x"0006B391",
    x"0006B0F3",
    x"0006AE56",
    x"0006ABBB",
    x"0006A920",
    x"0006A687",
    x"0006A3EE",
    x"0006A157",
    x"00069EC0",
    x"00069C2B",
    x"00069996",
    x"00069703",
    x"00069470",
    x"000691DF",
    x"00068F4E",
    x"00068CBF",
    x"00068A30",
    x"000687A3",
    x"00068516",
    x"0006828B",
    x"00068000",
    x"00067D77",
    x"00067AEE",
    x"00067867",
    x"000675E0",
    x"0006735B",
    x"000670D6",
    x"00066E52",
    x"00066BD0",
    x"0006694E",
    x"000666CD",
    x"0006644E",
    x"000661CF",
    x"00065F51",
    x"00065CD5",
    x"00065A59",
    x"000657DE",
    x"00065564",
    x"000652EB",
    x"00065073",
    x"00064DFD",
    x"00064B87",
    x"00064912",
    x"0006469D",
    x"0006442A",
    x"000641B8",
    x"00063F47",
    x"00063CD7",
    x"00063A67",
    x"000637F9",
    x"0006358C",
    x"0006331F",
    x"000630B4",
    x"00062E49",
    x"00062BE0",
    x"00062977",
    x"0006270F",
    x"000624A8",
    x"00062243",
    x"00061FDE",
    x"00061D7A",
    x"00061B17",
    x"000618B5",
    x"00061653",
    x"000613F3",
    x"00061194",
    x"00060F35",
    x"00060CD8",
    x"00060A7B",
    x"00060820",
    x"000605C5",
    x"0006036B",
    x"00060112",
    x"0005FEBA",
    x"0005FC63",
    x"0005FA0D",
    x"0005F7B8",
    x"0005F564",
    x"0005F310",
    x"0005F0BE",
    x"0005EE6C",
    x"0005EC1B",
    x"0005E9CC",
    x"0005E77D",
    x"0005E52F",
    x"0005E2E2",
    x"0005E096",
    x"0005DE4A",
    x"0005DC00",
    x"0005D9B6",
    x"0005D76E",
    x"0005D526",
    x"0005D2DF",
    x"0005D099",
    x"0005CE54",
    x"0005CC10",
    x"0005C9CD",
    x"0005C78B",
    x"0005C549",
    x"0005C308",
    x"0005C0C9",
    x"0005BE8A",
    x"0005BC4C",
    x"0005BA0F",
    x"0005B7D2",
    x"0005B597",
    x"0005B35D",
    x"0005B123",
    x"0005AEEA",
    x"0005ACB2",
    x"0005AA7B",
    x"0005A845",
    x"0005A610",
    x"0005A3DB",
    x"0005A1A8",
    x"00059F75",
    x"00059D43",
    x"00059B12",
    x"000598E2",
    x"000596B3",
    x"00059484",
    x"00059257",
    x"0005902A",
    x"00058DFE",
    x"00058BD3",
    x"000589A9",
    x"00058780",
    x"00058557",
    x"0005832F",
    x"00058109",
    x"00057EE3",
    x"00057CBD",
    x"00057A99",
    x"00057876",
    x"00057653",
    x"00057431",
    x"00057210",
    x"00056FF0",
    x"00056DD1",
    x"00056BB2",
    x"00056995",
    x"00056778",
    x"0005655C",
    x"00056341",
    x"00056126",
    x"00055F0D",
    x"00055CF4",
    x"00055ADC",
    x"000558C5",
    x"000556AF",
    x"00055499",
    x"00055285",
    x"00055071",
    x"00054E5E",
    x"00054C4C",
    x"00054A3A",
    x"0005482A",
    x"0005461A",
    x"0005440B",
    x"000541FD",
    x"00053FEF",
    x"00053DE3",
    x"00053BD7",
    x"000539CC",
    x"000537C2",
    x"000535B8",
    x"000533B0",
    x"000531A8",
    x"00052FA1",
    x"00052D9B",
    x"00052B95",
    x"00052991",
    x"0005278D",
    x"0005258A",
    x"00052388",
    x"00052186",
    x"00051F85",
    x"00051D85",
    x"00051B86",
    x"00051988",
    x"0005178A",
    x"0005158E",
    x"00051392",
    x"00051196",
    x"00050F9C",
    x"00050DA2",
    x"00050BA9",
    x"000509B1",
    x"000507BA",
    x"000505C3",
    x"000503CD",
    x"000501D8",
    x"0004FFE4",
    x"0004FDF0",
    x"0004FBFD",
    x"0004FA0B",
    x"0004F81A",
    x"0004F629",
    x"0004F43A",
    x"0004F24B",
    x"0004F05C",
    x"0004EE6F",
    x"0004EC82",
    x"0004EA96",
    x"0004E8AB",
    x"0004E6C0",
    x"0004E4D6",
    x"0004E2ED",
    x"0004E105",
    x"0004DF1E",
    x"0004DD37",
    x"0004DB51",
    x"0004D96C",
    x"0004D787",
    x"0004D5A3",
    x"0004D3C0",
    x"0004D1DE",
    x"0004CFFC",
    x"0004CE1B",
    x"0004CC3B",
    x"0004CA5C",
    x"0004C87D",
    x"0004C69F",
    x"0004C4C2",
    x"0004C2E5",
    x"0004C10A",
    x"0004BF2F",
    x"0004BD54",
    x"0004BB7B",
    x"0004B9A2",
    x"0004B7CA",
    x"0004B5F2",
    x"0004B41B",
    x"0004B245",
    x"0004B070",
    x"0004AE9C",
    x"0004ACC8",
    x"0004AAF5",
    x"0004A922",
    x"0004A750",
    x"0004A57F",
    x"0004A3AF",
    x"0004A1E0",
    x"0004A011",
    x"00049E43",
    x"00049C75",
    x"00049AA8",
    x"000498DC",
    x"00049711",
    x"00049546",
    x"0004937C",
    x"000491B3",
    x"00048FEA",
    x"00048E23",
    x"00048C5B",
    x"00048A95",
    x"000488CF",
    x"0004870A",
    x"00048546",
    x"00048382",
    x"000481BF",
    x"00047FFD",
    x"00047E3B",
    x"00047C7A",
    x"00047ABA",
    x"000478FA",
    x"0004773B",
    x"0004757D",
    x"000473BF",
    x"00047202",
    x"00047046",
    x"00046E8B",
    x"00046CD0",
    x"00046B16",
    x"0004695C",
    x"000467A3",
    x"000465EB",
    x"00046434",
    x"0004627D",
    x"000460C7",
    x"00045F11",
    x"00045D5D",
    x"00045BA8",
    x"000459F5",
    x"00045842",
    x"00045690",
    x"000454DF",
    x"0004532E",
    x"0004517E",
    x"00044FCE",
    x"00044E1F",
    x"00044C71",
    x"00044AC4",
    x"00044917",
    x"0004476A",
    x"000445BF",
    x"00044414",
    x"0004426A",
    x"000440C0",
    x"00043F17",
    x"00043D6F",
    x"00043BC7",
    x"00043A20",
    x"0004387A",
    x"000436D4",
    x"0004352F",
    x"0004338A",
    x"000431E7",
    x"00043043",
    x"00042EA1",
    x"00042CFF",
    x"00042B5E",
    x"000429BD",
    x"0004281D",
    x"0004267E",
    x"000424DF",
    x"00042341",
    x"000421A3",
    x"00042007",
    x"00041E6A",
    x"00041CCF",
    x"00041B34",
    x"0004199A",
    x"00041800",
    x"00041667",
    x"000414CE",
    x"00041337",
    x"0004119F",
    x"00041009",
    x"00040E73",
    x"00040CDE",
    x"00040B49",
    x"000409B5",
    x"00040821",
    x"0004068E",
    x"000404FC",
    x"0004036B",
    x"000401D9",
    x"00040049",
    x"0003FEB9",
    x"0003FD2A",
    x"0003FB9B",
    x"0003FA0D",
    x"0003F880",
    x"0003F6F3",
    x"0003F567",
    x"0003F3DC",
    x"0003F251",
    x"0003F0C6",
    x"0003EF3D",
    x"0003EDB3",
    x"0003EC2B",
    x"0003EAA3",
    x"0003E91C",
    x"0003E795",
    x"0003E60F",
    x"0003E489",
    x"0003E304",
    x"0003E180",
    x"0003DFFC",
    x"0003DE79",
    x"0003DCF6",
    x"0003DB74",
    x"0003D9F3",
    x"0003D872",
    x"0003D6F2",
    x"0003D572",
    x"0003D3F3",
    x"0003D274",
    x"0003D0F6",
    x"0003CF79",
    x"0003CDFC",
    x"0003CC80",
    x"0003CB05",
    x"0003C98A",
    x"0003C80F",
    x"0003C695",
    x"0003C51C",
    x"0003C3A3",
    x"0003C22B",
    x"0003C0B4",
    x"0003BF3D",
    x"0003BDC6",
    x"0003BC50",
    x"0003BADB",
    x"0003B966",
    x"0003B7F2",
    x"0003B67F",
    x"0003B50C",
    x"0003B399",
    x"0003B227",
    x"0003B0B6",
    x"0003AF45",
    x"0003ADD5",
    x"0003AC65",
    x"0003AAF6",
    x"0003A988",
    x"0003A81A",
    x"0003A6AD",
    x"0003A540",
    x"0003A3D3",
    x"0003A268",
    x"0003A0FD",
    x"00039F92",
    x"00039E28",
    x"00039CBE",
    x"00039B55",
    x"000399ED",
    x"00039885",
    x"0003971E",
    x"000395B7",
    x"00039451",
    x"000392EB",
    x"00039186",
    x"00039022",
    x"00038EBE",
    x"00038D5A",
    x"00038BF7",
    x"00038A95",
    x"00038933",
    x"000387D2",
    x"00038671",
    x"00038510",
    x"000383B1",
    x"00038252",
    x"000380F3",
    x"00037F95",
    x"00037E37",
    x"00037CDA",
    x"00037B7E",
    x"00037A22",
    x"000378C6",
    x"0003776B",
    x"00037611",
    x"000374B7",
    x"0003735E",
    x"00037205",
    x"000370AD",
    x"00036F55",
    x"00036DFE",
    x"00036CA7",
    x"00036B51",
    x"000369FB",
    x"000368A6",
    x"00036751",
    x"000365FD",
    x"000364AA",
    x"00036357",
    x"00036204",
    x"000360B2",
    x"00035F61",
    x"00035E10",
    x"00035CBF",
    x"00035B6F",
    x"00035A20",
    x"000358D1",
    x"00035782",
    x"00035634",
    x"000354E7",
    x"0003539A",
    x"0003524E",
    x"00035102",
    x"00034FB6",
    x"00034E6C",
    x"00034D21",
    x"00034BD7",
    x"00034A8E",
    x"00034945",
    x"000347FD",
    x"000346B5",
    x"0003456D",
    x"00034427",
    x"000342E0",
    x"0003419A",
    x"00034055",
    x"00033F10",
    x"00033DCC",
    x"00033C88",
    x"00033B44",
    x"00033A01",
    x"000338BF",
    x"0003377D",
    x"0003363C",
    x"000334FB",
    x"000333BA",
    x"0003327A",
    x"0003313B",
    x"00032FFC",
    x"00032EBD",
    x"00032D7F",
    x"00032C42",
    x"00032B05",
    x"000329C8",
    x"0003288C",
    x"00032751",
    x"00032615",
    x"000324DB",
    x"000323A1",
    x"00032267",
    x"0003212E",
    x"00031FF5",
    x"00031EBD",
    x"00031D85",
    x"00031C4E",
    x"00031B17",
    x"000319E1",
    x"000318AB",
    x"00031775",
    x"00031640",
    x"0003150C",
    x"000313D8",
    x"000312A4",
    x"00031171",
    x"0003103F",
    x"00030F0D",
    x"00030DDB",
    x"00030CAA",
    x"00030B79",
    x"00030A49",
    x"00030919",
    x"000307EA",
    x"000306BB",
    x"0003058C",
    x"0003045F",
    x"00030331",
    x"00030204",
    x"000300D8",
    x"0002FFAB",
    x"0002FE80",
    x"0002FD55",
    x"0002FC2A",
    x"0002FB00",
    x"0002F9D6",
    x"0002F8AC",
    x"0002F783",
    x"0002F65B",
    x"0002F533",
    x"0002F40B",
    x"0002F2E4",
    x"0002F1BE",
    x"0002F097",
    x"0002EF72",
    x"0002EE4C",
    x"0002ED28",
    x"0002EC03",
    x"0002EADF",
    x"0002E9BC",
    x"0002E899",
    x"0002E776",
    x"0002E654",
    x"0002E532",
    x"0002E411",
    x"0002E2F0",
    x"0002E1CF",
    x"0002E0AF",
    x"0002DF90",
    x"0002DE71",
    x"0002DD52",
    x"0002DC34",
    x"0002DB16",
    x"0002D9F9",
    x"0002D8DC",
    x"0002D7BF",
    x"0002D6A3",
    x"0002D588",
    x"0002D46C",
    x"0002D352",
    x"0002D237",
    x"0002D11D",
    x"0002D004",
    x"0002CEEB",
    x"0002CDD2",
    x"0002CCBA",
    x"0002CBA2",
    x"0002CA8B",
    x"0002C974",
    x"0002C85E",
    x"0002C748",
    x"0002C632",
    x"0002C51D",
    x"0002C408",
    x"0002C2F4",
    x"0002C1E0",
    x"0002C0CC",
    x"0002BFB9",
    x"0002BEA6",
    x"0002BD94",
    x"0002BC82",
    x"0002BB71",
    x"0002BA60",
    x"0002B94F",
    x"0002B83F",
    x"0002B72F",
    x"0002B620",
    x"0002B511",
    x"0002B402",
    x"0002B2F4",
    x"0002B1E7",
    x"0002B0D9",
    x"0002AFCC",
    x"0002AEC0",
    x"0002ADB4",
    x"0002ACA8",
    x"0002AB9D",
    x"0002AA92",
    x"0002A988",
    x"0002A87E",
    x"0002A774",
    x"0002A66B",
    x"0002A562",
    x"0002A45A",
    x"0002A352",
    x"0002A24A",
    x"0002A143",
    x"0002A03C",
    x"00029F36",
    x"00029E30",
    x"00029D2A",
    x"00029C25",
    x"00029B20",
    x"00029A1C",
    x"00029918",
    x"00029814",
    x"00029711",
    x"0002960E",
    x"0002950C",
    x"0002940A",
    x"00029308",
    x"00029207",
    x"00029106",
    x"00029006",
    x"00028F05",
    x"00028E06",
    x"00028D07",
    x"00028C08",
    x"00028B09",
    x"00028A0B",
    x"0002890D",
    x"00028810",
    x"00028713",
    x"00028616",
    x"0002851A",
    x"0002841E",
    x"00028323",
    x"00028228",
    x"0002812D",
    x"00028033",
    x"00027F39",
    x"00027E40",
    x"00027D47",
    x"00027C4E",
    x"00027B55",
    x"00027A5D",
    x"00027966",
    x"0002786F",
    x"00027778",
    x"00027681",
    x"0002758B",
    x"00027495",
    x"000273A0",
    x"000272AB",
    x"000271B6",
    x"000270C2",
    x"00026FCE",
    x"00026EDB",
    x"00026DE8",
    x"00026CF5",
    x"00026C03",
    x"00026B11",
    x"00026A1F",
    x"0002692E",
    x"0002683D",
    x"0002674C",
    x"0002665C",
    x"0002656C",
    x"0002647D",
    x"0002638E",
    x"0002629F",
    x"000261B1",
    x"000260C3",
    x"00025FD5",
    x"00025EE8",
    x"00025DFB",
    x"00025D0F",
    x"00025C22",
    x"00025B37",
    x"00025A4B",
    x"00025960",
    x"00025875",
    x"0002578B",
    x"000256A1",
    x"000255B7",
    x"000254CE",
    x"000253E5",
    x"000252FC",
    x"00025214",
    x"0002512C",
    x"00025045",
    x"00024F5E",
    x"00024E77",
    x"00024D90",
    x"00024CAA",
    x"00024BC4",
    x"00024ADF",
    x"000249FA",
    x"00024915",
    x"00024831",
    x"0002474D",
    x"00024669",
    x"00024586",
    x"000244A3",
    x"000243C0",
    x"000242DE",
    x"000241FC",
    x"0002411A",
    x"00024039",
    x"00023F58",
    x"00023E78",
    x"00023D97",
    x"00023CB7",
    x"00023BD8",
    x"00023AF9",
    x"00023A1A",
    x"0002393B",
    x"0002385D",
    x"0002377F",
    x"000236A2",
    x"000235C5",
    x"000234E8",
    x"0002340B",
    x"0002332F",
    x"00023253",
    x"00023178",
    x"0002309D",
    x"00022FC2",
    x"00022EE7",
    x"00022E0D",
    x"00022D33",
    x"00022C5A",
    x"00022B81",
    x"00022AA8",
    x"000229CF",
    x"000228F7",
    x"0002281F",
    x"00022748",
    x"00022671",
    x"0002259A",
    x"000224C3",
    x"000223ED",
    x"00022317",
    x"00022242",
    x"0002216C",
    x"00022098",
    x"00021FC3",
    x"00021EEF",
    x"00021E1B",
    x"00021D47",
    x"00021C74",
    x"00021BA1",
    x"00021ACE",
    x"000219FC",
    x"0002192A",
    x"00021858",
    x"00021787",
    x"000216B6",
    x"000215E5",
    x"00021515",
    x"00021445",
    x"00021375",
    x"000212A6",
    x"000211D6",
    x"00021108",
    x"00021039",
    x"00020F6B",
    x"00020E9D",
    x"00020DD0",
    x"00020D02",
    x"00020C35",
    x"00020B69",
    x"00020A9C",
    x"000209D0",
    x"00020905",
    x"00020839",
    x"0002076E",
    x"000206A4",
    x"000205D9",
    x"0002050F",
    x"00020445",
    x"0002037C",
    x"000202B3",
    x"000201EA",
    x"00020121",
    x"00020059",
    x"0001FF91",
    x"0001FEC9",
    x"0001FE02",
    x"0001FD3B",
    x"0001FC74",
    x"0001FBAD",
    x"0001FAE7",
    x"0001FA21",
    x"0001F95C",
    x"0001F897",
    x"0001F7D2",
    x"0001F70D",
    x"0001F649",
    x"0001F585",
    x"0001F4C1",
    x"0001F3FD",
    x"0001F33A",
    x"0001F277",
    x"0001F1B5",
    x"0001F0F2",
    x"0001F031",
    x"0001EF6F",
    x"0001EEAD",
    x"0001EDEC",
    x"0001ED2C",
    x"0001EC6B",
    x"0001EBAB",
    x"0001EAEB",
    x"0001EA2B",
    x"0001E96C",
    x"0001E8AD",
    x"0001E7EE",
    x"0001E730",
    x"0001E672",
    x"0001E5B4",
    x"0001E4F6",
    x"0001E439",
    x"0001E37C",
    x"0001E2BF",
    x"0001E203",
    x"0001E147",
    x"0001E08B",
    x"0001DFCF",
    x"0001DF14",
    x"0001DE59",
    x"0001DD9E",
    x"0001DCE4",
    x"0001DC2A",
    x"0001DB70",
    x"0001DAB6",
    x"0001D9FD",
    x"0001D944",
    x"0001D88B",
    x"0001D7D3",
    x"0001D71B",
    x"0001D663",
    x"0001D5AB",
    x"0001D4F4",
    x"0001D43D",
    x"0001D386",
    x"0001D2CF",
    x"0001D219",
    x"0001D163",
    x"0001D0AE",
    x"0001CFF8",
    x"0001CF43",
    x"0001CE8E",
    x"0001CDDA",
    x"0001CD26",
    x"0001CC72",
    x"0001CBBE",
    x"0001CB0A",
    x"0001CA57",
    x"0001C9A4",
    x"0001C8F2",
    x"0001C83F",
    x"0001C78D",
    x"0001C6DB",
    x"0001C62A",
    x"0001C579",
    x"0001C4C8",
    x"0001C417",
    x"0001C366",
    x"0001C2B6",
    x"0001C206",
    x"0001C157",
    x"0001C0A7",
    x"0001BFF8",
    x"0001BF49",
    x"0001BE9B",
    x"0001BDEC",
    x"0001BD3E",
    x"0001BC90",
    x"0001BBE3",
    x"0001BB36",
    x"0001BA89",
    x"0001B9DC",
    x"0001B92F",
    x"0001B883",
    x"0001B7D7",
    x"0001B72C",
    x"0001B680",
    x"0001B5D5",
    x"0001B52A",
    x"0001B480",
    x"0001B3D5",
    x"0001B32B",
    x"0001B281",
    x"0001B1D8",
    x"0001B12E",
    x"0001B085",
    x"0001AFDC",
    x"0001AF34",
    x"0001AE8B",
    x"0001ADE3",
    x"0001AD3C",
    x"0001AC94",
    x"0001ABED",
    x"0001AB46",
    x"0001AA9F",
    x"0001A9F8",
    x"0001A952",
    x"0001A8AC",
    x"0001A806",
    x"0001A761",
    x"0001A6BC",
    x"0001A617",
    x"0001A572",
    x"0001A4CD",
    x"0001A429",
    x"0001A385",
    x"0001A2E1",
    x"0001A23E",
    x"0001A19B",
    x"0001A0F8",
    x"0001A055",
    x"00019FB2",
    x"00019F10",
    x"00019E6E",
    x"00019DCC",
    x"00019D2B",
    x"00019C8A",
    x"00019BE9",
    x"00019B48",
    x"00019AA7",
    x"00019A07",
    x"00019967",
    x"000198C7",
    x"00019828",
    x"00019788",
    x"000196E9",
    x"0001964A",
    x"000195AC",
    x"0001950D",
    x"0001946F",
    x"000193D1",
    x"00019334",
    x"00019296",
    x"000191F9",
    x"0001915C",
    x"000190C0",
    x"00019023",
    x"00018F87",
    x"00018EEB",
    x"00018E4F",
    x"00018DB4",
    x"00018D19",
    x"00018C7E",
    x"00018BE3",
    x"00018B48",
    x"00018AAE",
    x"00018A14",
    x"0001897A",
    x"000188E1",
    x"00018847",
    x"000187AE",
    x"00018715",
    x"0001867D",
    x"000185E4",
    x"0001854C",
    x"000184B4",
    x"0001841C",
    x"00018385",
    x"000182EE",
    x"00018257",
    x"000181C0",
    x"00018129",
    x"00018093",
    x"00017FFD",
    x"00017F67",
    x"00017ED1",
    x"00017E3C",
    x"00017DA7",
    x"00017D12",
    x"00017C7D",
    x"00017BE8",
    x"00017B54",
    x"00017AC0",
    x"00017A2C",
    x"00017999",
    x"00017905",
    x"00017872",
    x"000177DF",
    x"0001774C",
    x"000176BA",
    x"00017628",
    x"00017596",
    x"00017504",
    x"00017472",
    x"000173E1",
    x"00017350",
    x"000172BF",
    x"0001722E",
    x"0001719E",
    x"0001710D",
    x"0001707D",
    x"00016FED",
    x"00016F5E",
    x"00016ECE",
    x"00016E3F",
    x"00016DB0",
    x"00016D22",
    x"00016C93",
    x"00016C05",
    x"00016B77",
    x"00016AE9",
    x"00016A5B",
    x"000169CE",
    x"00016940",
    x"000168B3",
    x"00016827",
    x"0001679A",
    x"0001670E",
    x"00016682",
    x"000165F6",
    x"0001656A",
    x"000164DE",
    x"00016453",
    x"000163C8",
    x"0001633D",
    x"000162B3",
    x"00016228",
    x"0001619E",
    x"00016114",
    x"0001608A",
    x"00016000",
    x"00015F77",
    x"00015EEE",
    x"00015E65",
    x"00015DDC",
    x"00015D53",
    x"00015CCB",
    x"00015C43",
    x"00015BBB",
    x"00015B33",
    x"00015AAC",
    x"00015A24",
    x"0001599D",
    x"00015916",
    x"00015890",
    x"00015809",
    x"00015783",
    x"000156FD",
    x"00015677",
    x"000155F1",
    x"0001556C",
    x"000154E7",
    x"00015462",
    x"000153DD",
    x"00015358",
    x"000152D4",
    x"0001524F",
    x"000151CB",
    x"00015147",
    x"000150C4",
    x"00015040",
    x"00014FBD",
    x"00014F3A",
    x"00014EB7",
    x"00014E35",
    x"00014DB2",
    x"00014D30",
    x"00014CAE",
    x"00014C2C",
    x"00014BAA",
    x"00014B29",
    x"00014AA8",
    x"00014A27",
    x"000149A6",
    x"00014925",
    x"000148A4",
    x"00014824",
    x"000147A4",
    x"00014724",
    x"000146A5",
    x"00014625",
    x"000145A6",
    x"00014527",
    x"000144A8",
    x"00014429",
    x"000143AA",
    x"0001432C",
    x"000142AE",
    x"00014230",
    x"000141B2",
    x"00014135",
    x"000140B7",
    x"0001403A",
    x"00013FBD",
    x"00013F40",
    x"00013EC4",
    x"00013E47",
    x"00013DCB",
    x"00013D4F",
    x"00013CD3",
    x"00013C58",
    x"00013BDC",
    x"00013B61",
    x"00013AE6",
    x"00013A6B",
    x"000139F0",
    x"00013975",
    x"000138FB",
    x"00013881",
    x"00013807",
    x"0001378D",
    x"00013714",
    x"0001369A",
    x"00013621",
    x"000135A8",
    x"0001352F",
    x"000134B6",
    x"0001343E",
    x"000133C6",
    x"0001334D",
    x"000132D5",
    x"0001325E",
    x"000131E6",
    x"0001316F",
    x"000130F7",
    x"00013080",
    x"0001300A",
    x"00012F93",
    x"00012F1C",
    x"00012EA6",
    x"00012E30",
    x"00012DBA",
    x"00012D44",
    x"00012CCF",
    x"00012C59",
    x"00012BE4",
    x"00012B6F",
    x"00012AFA",
    x"00012A85",
    x"00012A11",
    x"0001299D",
    x"00012928",
    x"000128B4",
    x"00012841",
    x"000127CD",
    x"00012759",
    x"000126E6",
    x"00012673",
    x"00012600",
    x"0001258D",
    x"0001251B",
    x"000124A8",
    x"00012436",
    x"000123C4",
    x"00012352",
    x"000122E1",
    x"0001226F",
    x"000121FE",
    x"0001218C",
    x"0001211B",
    x"000120AB",
    x"0001203A",
    x"00011FC9",
    x"00011F59",
    x"00011EE9",
    x"00011E79",
    x"00011E09",
    x"00011D99",
    x"00011D2A",
    x"00011CBB",
    x"00011C4C",
    x"00011BDD",
    x"00011B6E",
    x"00011AFF",
    x"00011A91",
    x"00011A22",
    x"000119B4",
    x"00011946",
    x"000118D8",
    x"0001186B",
    x"000117FD",
    x"00011790",
    x"00011723",
    x"000116B6",
    x"00011649",
    x"000115DD",
    x"00011570",
    x"00011504",
    x"00011498",
    x"0001142C",
    x"000113C0",
    x"00011354",
    x"000112E9",
    x"0001127E",
    x"00011212",
    x"000111A7",
    x"0001113D",
    x"000110D2",
    x"00011068",
    x"00010FFD",
    x"00010F93",
    x"00010F29",
    x"00010EBF",
    x"00010E56",
    x"00010DEC",
    x"00010D83",
    x"00010D19",
    x"00010CB0",
    x"00010C48",
    x"00010BDF",
    x"00010B76",
    x"00010B0E",
    x"00010AA6",
    x"00010A3E",
    x"000109D6",
    x"0001096E",
    x"00010906",
    x"0001089F",
    x"00010838",
    x"000107D0",
    x"00010769",
    x"00010703",
    x"0001069C",
    x"00010635",
    x"000105CF",
    x"00010569",
    x"00010503",
    x"0001049D",
    x"00010437",
    x"000103D2",
    x"0001036C",
    x"00010307",
    x"000102A2",
    x"0001023D",
    x"000101D8",
    x"00010174",
    x"0001010F",
    x"000100AB",
    x"00010046",
    x"0000FFE2",
    x"0000FF7F",
    x"0000FF1B",
    x"0000FEB7",
    x"0000FE54",
    x"0000FDF1",
    x"0000FD8D",
    x"0000FD2A",
    x"0000FCC8",
    x"0000FC65",
    x"0000FC02",
    x"0000FBA0",
    x"0000FB3E",
    x"0000FADC",
    x"0000FA7A",
    x"0000FA18",
    x"0000F9B7",
    x"0000F955",
    x"0000F8F4",
    x"0000F893",
    x"0000F832",
    x"0000F7D1",
    x"0000F770",
    x"0000F70F",
    x"0000F6AF",
    x"0000F64F",
    x"0000F5EF",
    x"0000F58F",
    x"0000F52F",
    x"0000F4CF",
    x"0000F46F",
    x"0000F410",
    x"0000F3B1",
    x"0000F352",
    x"0000F2F3",
    x"0000F294",
    x"0000F235",
    x"0000F1D7",
    x"0000F178",
    x"0000F11A",
    x"0000F0BC",
    x"0000F05E",
    x"0000F000",
    x"0000EFA2",
    x"0000EF45",
    x"0000EEE7",
    x"0000EE8A",
    x"0000EE2D",
    x"0000EDD0",
    x"0000ED73",
    x"0000ED17",
    x"0000ECBA",
    x"0000EC5E",
    x"0000EC01",
    x"0000EBA5",
    x"0000EB49",
    x"0000EAED",
    x"0000EA92",
    x"0000EA36",
    x"0000E9DB",
    x"0000E980",
    x"0000E924",
    x"0000E8C9",
    x"0000E86F",
    x"0000E814",
    x"0000E7B9",
    x"0000E75F",
    x"0000E704",
    x"0000E6AA",
    x"0000E650",
    x"0000E5F6",
    x"0000E59D",
    x"0000E543",
    x"0000E4E9",
    x"0000E490",
    x"0000E437",
    x"0000E3DE",
    x"0000E385",
    x"0000E32C",
    x"0000E2D3",
    x"0000E27B",
    x"0000E222",
    x"0000E1CA",
    x"0000E172",
    x"0000E11A",
    x"0000E0C2",
    x"0000E06A",
    x"0000E013",
    x"0000DFBB",
    x"0000DF64",
    x"0000DF0D",
    x"0000DEB6",
    x"0000DE5F",
    x"0000DE08",
    x"0000DDB1",
    x"0000DD5B",
    x"0000DD04",
    x"0000DCAE",
    x"0000DC58",
    x"0000DC02",
    x"0000DBAC",
    x"0000DB56",
    x"0000DB01",
    x"0000DAAB",
    x"0000DA56",
    x"0000DA01",
    x"0000D9AC",
    x"0000D957",
    x"0000D902",
    x"0000D8AD",
    x"0000D859",
    x"0000D804",
    x"0000D7B0",
    x"0000D75C",
    x"0000D708",
    x"0000D6B4",
    x"0000D660",
    x"0000D60C",
    x"0000D5B9",
    x"0000D565",
    x"0000D512",
    x"0000D4BF",
    x"0000D46C",
    x"0000D419",
    x"0000D3C6",
    x"0000D373",
    x"0000D321",
    x"0000D2CE",
    x"0000D27C",
    x"0000D22A",
    x"0000D1D8",
    x"0000D186",
    x"0000D134",
    x"0000D0E3",
    x"0000D091",
    x"0000D040",
    x"0000CFEE",
    x"0000CF9D",
    x"0000CF4C",
    x"0000CEFB",
    x"0000CEAA",
    x"0000CE5A",
    x"0000CE09",
    x"0000CDB9",
    x"0000CD69",
    x"0000CD18",
    x"0000CCC8",
    x"0000CC78",
    x"0000CC29",
    x"0000CBD9",
    x"0000CB89",
    x"0000CB3A",
    x"0000CAEB",
    x"0000CA9B",
    x"0000CA4C",
    x"0000C9FD",
    x"0000C9AE",
    x"0000C960",
    x"0000C911",
    x"0000C8C3",
    x"0000C874",
    x"0000C826",
    x"0000C7D8",
    x"0000C78A",
    x"0000C73C",
    x"0000C6EE",
    x"0000C6A1",
    x"0000C653",
    x"0000C606",
    x"0000C5B8",
    x"0000C56B",
    x"0000C51E",
    x"0000C4D1",
    x"0000C484",
    x"0000C438",
    x"0000C3EB",
    x"0000C39F",
    x"0000C352",
    x"0000C306",
    x"0000C2BA",
    x"0000C26E",
    x"0000C222",
    x"0000C1D6",
    x"0000C18B",
    x"0000C13F",
    x"0000C0F4",
    x"0000C0A8",
    x"0000C05D",
    x"0000C012",
    x"0000BFC7",
    x"0000BF7C",
    x"0000BF31",
    x"0000BEE7",
    x"0000BE9C",
    x"0000BE52",
    x"0000BE08",
    x"0000BDBD",
    x"0000BD73",
    x"0000BD29",
    x"0000BCE0",
    x"0000BC96",
    x"0000BC4C",
    x"0000BC03",
    x"0000BBB9",
    x"0000BB70",
    x"0000BB27",
    x"0000BADE",
    x"0000BA95",
    x"0000BA4C",
    x"0000BA03",
    x"0000B9BB",
    x"0000B972",
    x"0000B92A",
    x"0000B8E2",
    x"0000B899",
    x"0000B851",
    x"0000B809",
    x"0000B7C2",
    x"0000B77A",
    x"0000B732",
    x"0000B6EB",
    x"0000B6A3",
    x"0000B65C",
    x"0000B615",
    x"0000B5CE",
    x"0000B587",
    x"0000B540",
    x"0000B4F9",
    x"0000B4B3",
    x"0000B46C",
    x"0000B426",
    x"0000B3DF",
    x"0000B399",
    x"0000B353",
    x"0000B30D",
    x"0000B2C7",
    x"0000B281",
    x"0000B23C",
    x"0000B1F6",
    x"0000B1B1",
    x"0000B16B",
    x"0000B126",
    x"0000B0E1",
    x"0000B09C",
    x"0000B057",
    x"0000B012",
    x"0000AFCD",
    x"0000AF89",
    x"0000AF44",
    x"0000AF00",
    x"0000AEBC",
    x"0000AE77",
    x"0000AE33",
    x"0000ADEF",
    x"0000ADAB",
    x"0000AD68",
    x"0000AD24",
    x"0000ACE0",
    x"0000AC9D",
    x"0000AC59",
    x"0000AC16",
    x"0000ABD3",
    x"0000AB90",
    x"0000AB4D",
    x"0000AB0A",
    x"0000AAC7",
    x"0000AA85",
    x"0000AA42",
    x"0000AA00",
    x"0000A9BD",
    x"0000A97B",
    x"0000A939",
    x"0000A8F7",
    x"0000A8B5",
    x"0000A873",
    x"0000A831",
    x"0000A7F0",
    x"0000A7AE",
    x"0000A76D",
    x"0000A72B",
    x"0000A6EA",
    x"0000A6A9",
    x"0000A668",
    x"0000A627",
    x"0000A5E6",
    x"0000A5A5",
    x"0000A565",
    x"0000A524",
    x"0000A4E4",
    x"0000A4A3",
    x"0000A463",
    x"0000A423",
    x"0000A3E3",
    x"0000A3A3",
    x"0000A363",
    x"0000A323",
    x"0000A2E3",
    x"0000A2A4",
    x"0000A264",
    x"0000A225",
    x"0000A1E6",
    x"0000A1A7",
    x"0000A167",
    x"0000A128",
    x"0000A0EA",
    x"0000A0AB",
    x"0000A06C",
    x"0000A02D",
    x"00009FEF",
    x"00009FB0",
    x"00009F72",
    x"00009F34",
    x"00009EF6",
    x"00009EB8",
    x"00009E7A",
    x"00009E3C",
    x"00009DFE",
    x"00009DC0",
    x"00009D83",
    x"00009D45",
    x"00009D08",
    x"00009CCB",
    x"00009C8E",
    x"00009C50",
    x"00009C13",
    x"00009BD6",
    x"00009B9A",
    x"00009B5D",
    x"00009B20",
    x"00009AE4",
    x"00009AA7",
    x"00009A6B",
    x"00009A2F",
    x"000099F2",
    x"000099B6",
    x"0000997A",
    x"0000993E",
    x"00009903",
    x"000098C7",
    x"0000988B",
    x"00009850",
    x"00009814",
    x"000097D9",
    x"0000979E",
    x"00009762",
    x"00009727",
    x"000096EC",
    x"000096B1",
    x"00009677",
    x"0000963C",
    x"00009601",
    x"000095C7",
    x"0000958C",
    x"00009552",
    x"00009518",
    x"000094DD",
    x"000094A3",
    x"00009469",
    x"0000942F",
    x"000093F6",
    x"000093BC",
    x"00009382",
    x"00009349",
    x"0000930F",
    x"000092D6",
    x"0000929C",
    x"00009263",
    x"0000922A",
    x"000091F1",
    x"000091B8",
    x"0000917F",
    x"00009146",
    x"0000910E",
    x"000090D5",
    x"0000909C",
    x"00009064",
    x"0000902C",
    x"00008FF3",
    x"00008FBB",
    x"00008F83",
    x"00008F4B",
    x"00008F13",
    x"00008EDB",
    x"00008EA4",
    x"00008E6C",
    x"00008E34",
    x"00008DFD",
    x"00008DC5",
    x"00008D8E",
    x"00008D57",
    x"00008D20",
    x"00008CE8",
    x"00008CB1",
    x"00008C7B",
    x"00008C44",
    x"00008C0D",
    x"00008BD6",
    x"00008BA0",
    x"00008B69",
    x"00008B33",
    x"00008AFC",
    x"00008AC6",
    x"00008A90",
    x"00008A5A",
    x"00008A24",
    x"000089EE",
    x"000089B8",
    x"00008982",
    x"0000894D",
    x"00008917",
    x"000088E2",
    x"000088AC",
    x"00008877",
    x"00008842",
    x"0000880C",
    x"000087D7",
    x"000087A2",
    x"0000876D",
    x"00008739",
    x"00008704",
    x"000086CF",
    x"0000869A",
    x"00008666",
    x"00008631",
    x"000085FD",
    x"000085C9",
    x"00008595",
    x"00008560",
    x"0000852C",
    x"000084F8",
    x"000084C4",
    x"00008491",
    x"0000845D",
    x"00008429",
    x"000083F6",
    x"000083C2",
    x"0000838F",
    x"0000835B",
    x"00008328",
    x"000082F5",
    x"000082C2",
    x"0000828F",
    x"0000825C",
    x"00008229",
    x"000081F6",
    x"000081C3",
    x"00008191",
    x"0000815E",
    x"0000812C",
    x"000080F9",
    x"000080C7",
    x"00008095",
    x"00008062",
    x"00008030",
    x"00007FFE",
    x"00007FCC",
    x"00007F9A",
    x"00007F69",
    x"00007F37",
    x"00007F05",
    x"00007ED4",
    x"00007EA2",
    x"00007E71",
    x"00007E3F",
    x"00007E0E",
    x"00007DDD",
    x"00007DAC",
    x"00007D7B",
    x"00007D4A",
    x"00007D19",
    x"00007CE8",
    x"00007CB7",
    x"00007C87",
    x"00007C56",
    x"00007C25",
    x"00007BF5",
    x"00007BC5",
    x"00007B94",
    x"00007B64",
    x"00007B34",
    x"00007B04",
    x"00007AD4",
    x"00007AA4",
    x"00007A74",
    x"00007A44",
    x"00007A14",
    x"000079E5",
    x"000079B5",
    x"00007986",
    x"00007956",
    x"00007927",
    x"000078F8",
    x"000078C8",
    x"00007899",
    x"0000786A",
    x"0000783B",
    x"0000780C",
    x"000077DD",
    x"000077AF",
    x"00007780",
    x"00007751",
    x"00007723",
    x"000076F4",
    x"000076C6",
    x"00007697",
    x"00007669",
    x"0000763B",
    x"0000760D",
    x"000075DF",
    x"000075B1",
    x"00007583",
    x"00007555",
    x"00007527",
    x"000074F9",
    x"000074CC",
    x"0000749E",
    x"00007471",
    x"00007443",
    x"00007416",
    x"000073E8",
    x"000073BB",
    x"0000738E",
    x"00007361",
    x"00007334",
    x"00007307",
    x"000072DA",
    x"000072AD",
    x"00007280",
    x"00007254",
    x"00007227",
    x"000071FB",
    x"000071CE",
    x"000071A2",
    x"00007175",
    x"00007149",
    x"0000711D",
    x"000070F1",
    x"000070C5",
    x"00007099",
    x"0000706D",
    x"00007041",
    x"00007015",
    x"00006FE9",
    x"00006FBD",
    x"00006F92",
    x"00006F66",
    x"00006F3B",
    x"00006F0F",
    x"00006EE4",
    x"00006EB9",
    x"00006E8E",
    x"00006E62",
    x"00006E37",
    x"00006E0C",
    x"00006DE1",
    x"00006DB6",
    x"00006D8C",
    x"00006D61",
    x"00006D36",
    x"00006D0C",
    x"00006CE1",
    x"00006CB6",
    x"00006C8C",
    x"00006C62",
    x"00006C37",
    x"00006C0D",
    x"00006BE3",
    x"00006BB9",
    x"00006B8F",
    x"00006B65",
    x"00006B3B",
    x"00006B11",
    x"00006AE7",
    x"00006ABD",
    x"00006A94",
    x"00006A6A",
    x"00006A41",
    x"00006A17",
    x"000069EE",
    x"000069C4",
    x"0000699B",
    x"00006972",
    x"00006949",
    x"00006920",
    x"000068F7",
    x"000068CE",
    x"000068A5",
    x"0000687C",
    x"00006853",
    x"0000682A",
    x"00006802",
    x"000067D9",
    x"000067B1",
    x"00006788",
    x"00006760",
    x"00006737",
    x"0000670F",
    x"000066E7",
    x"000066BF",
    x"00006697",
    x"0000666F",
    x"00006647",
    x"0000661F",
    x"000065F7",
    x"000065CF",
    x"000065A7",
    x"00006580",
    x"00006558",
    x"00006530",
    x"00006509",
    x"000064E2",
    x"000064BA",
    x"00006493",
    x"0000646C",
    x"00006444",
    x"0000641D",
    x"000063F6",
    x"000063CF",
    x"000063A8",
    x"00006381",
    x"0000635A",
    x"00006334",
    x"0000630D",
    x"000062E6",
    x"000062C0",
    x"00006299",
    x"00006273",
    x"0000624C",
    x"00006226",
    x"00006200",
    x"000061D9",
    x"000061B3",
    x"0000618D",
    x"00006167",
    x"00006141",
    x"0000611B",
    x"000060F5",
    x"000060CF",
    x"000060A9",
    x"00006084",
    x"0000605E",
    x"00006038",
    x"00006013",
    x"00005FED",
    x"00005FC8",
    x"00005FA2",
    x"00005F7D",
    x"00005F58",
    x"00005F33",
    x"00005F0D",
    x"00005EE8",
    x"00005EC3",
    x"00005E9E",
    x"00005E79",
    x"00005E55",
    x"00005E30",
    x"00005E0B",
    x"00005DE6",
    x"00005DC2",
    x"00005D9D",
    x"00005D78",
    x"00005D54",
    x"00005D30",
    x"00005D0B",
    x"00005CE7",
    x"00005CC3",
    x"00005C9E",
    x"00005C7A",
    x"00005C56",
    x"00005C32",
    x"00005C0E",
    x"00005BEA",
    x"00005BC6",
    x"00005BA2",
    x"00005B7F",
    x"00005B5B",
    x"00005B37",
    x"00005B14",
    x"00005AF0",
    x"00005ACD",
    x"00005AA9",
    x"00005A86",
    x"00005A63",
    x"00005A3F",
    x"00005A1C",
    x"000059F9",
    x"000059D6",
    x"000059B3",
    x"00005990",
    x"0000596D",
    x"0000594A",
    x"00005927",
    x"00005904",
    x"000058E1",
    x"000058BF",
    x"0000589C",
    x"00005879",
    x"00005857",
    x"00005834",
    x"00005812",
    x"000057F0",
    x"000057CD",
    x"000057AB",
    x"00005789",
    x"00005767",
    x"00005745",
    x"00005723",
    x"00005700",
    x"000056DF",
    x"000056BD",
    x"0000569B",
    x"00005679",
    x"00005657",
    x"00005636",
    x"00005614",
    x"000055F2",
    x"000055D1",
    x"000055AF",
    x"0000558E",
    x"0000556C",
    x"0000554B",
    x"0000552A",
    x"00005509",
    x"000054E7",
    x"000054C6",
    x"000054A5",
    x"00005484",
    x"00005463",
    x"00005442",
    x"00005421",
    x"00005400",
    x"000053E0",
    x"000053BF",
    x"0000539E",
    x"0000537E",
    x"0000535D",
    x"0000533C",
    x"0000531C",
    x"000052FB",
    x"000052DB",
    x"000052BB",
    x"0000529A",
    x"0000527A",
    x"0000525A",
    x"0000523A",
    x"0000521A",
    x"000051FA",
    x"000051DA",
    x"000051BA",
    x"0000519A",
    x"0000517A",
    x"0000515A",
    x"0000513A",
    x"0000511B",
    x"000050FB",
    x"000050DC",
    x"000050BC",
    x"0000509C",
    x"0000507D",
    x"0000505E",
    x"0000503E",
    x"0000501F",
    x"00005000",
    x"00004FE0",
    x"00004FC1",
    x"00004FA2",
    x"00004F83",
    x"00004F64",
    x"00004F45",
    x"00004F26",
    x"00004F07",
    x"00004EE8",
    x"00004EC9",
    x"00004EAB",
    x"00004E8C",
    x"00004E6D",
    x"00004E4F",
    x"00004E30",
    x"00004E12",
    x"00004DF3",
    x"00004DD5",
    x"00004DB6",
    x"00004D98",
    x"00004D7A",
    x"00004D5C",
    x"00004D3D",
    x"00004D1F",
    x"00004D01",
    x"00004CE3",
    x"00004CC5",
    x"00004CA7",
    x"00004C89",
    x"00004C6B",
    x"00004C4D",
    x"00004C30",
    x"00004C12",
    x"00004BF4",
    x"00004BD7",
    x"00004BB9",
    x"00004B9B",
    x"00004B7E",
    x"00004B60",
    x"00004B43",
    x"00004B26",
    x"00004B08",
    x"00004AEB",
    x"00004ACE",
    x"00004AB1",
    x"00004A93",
    x"00004A76",
    x"00004A59",
    x"00004A3C",
    x"00004A1F",
    x"00004A02",
    x"000049E5",
    x"000049C9",
    x"000049AC",
    x"0000498F",
    x"00004972",
    x"00004956",
    x"00004939",
    x"0000491C",
    x"00004900",
    x"000048E3",
    x"000048C7",
    x"000048AB",
    x"0000488E",
    x"00004872",
    x"00004856",
    x"00004839",
    x"0000481D",
    x"00004801",
    x"000047E5",
    x"000047C9",
    x"000047AD",
    x"00004791",
    x"00004775",
    x"00004759",
    x"0000473D",
    x"00004721",
    x"00004706",
    x"000046EA",
    x"000046CE",
    x"000046B3",
    x"00004697",
    x"0000467B",
    x"00004660",
    x"00004644",
    x"00004629",
    x"0000460E",
    x"000045F2",
    x"000045D7",
    x"000045BC",
    x"000045A1",
    x"00004585",
    x"0000456A",
    x"0000454F",
    x"00004534",
    x"00004519",
    x"000044FE",
    x"000044E3",
    x"000044C8",
    x"000044AD",
    x"00004493",
    x"00004478",
    x"0000445D",
    x"00004442",
    x"00004428",
    x"0000440D",
    x"000043F3",
    x"000043D8",
    x"000043BE",
    x"000043A3",
    x"00004389",
    x"0000436E",
    x"00004354",
    x"0000433A",
    x"00004320",
    x"00004305",
    x"000042EB",
    x"000042D1",
    x"000042B7",
    x"0000429D",
    x"00004283",
    x"00004269",
    x"0000424F",
    x"00004235",
    x"0000421B",
    x"00004202",
    x"000041E8",
    x"000041CE",
    x"000041B4",
    x"0000419B",
    x"00004181",
    x"00004168",
    x"0000414E",
    x"00004135",
    x"0000411B",
    x"00004102",
    x"000040E8",
    x"000040CF",
    x"000040B6",
    x"0000409C",
    x"00004083",
    x"0000406A",
    x"00004051",
    x"00004038",
    x"0000401F",
    x"00004006",
    x"00003FED",
    x"00003FD4",
    x"00003FBB",
    x"00003FA2",
    x"00003F89",
    x"00003F70",
    x"00003F58",
    x"00003F3F",
    x"00003F26",
    x"00003F0D",
    x"00003EF5",
    x"00003EDC",
    x"00003EC4",
    x"00003EAB",
    x"00003E93",
    x"00003E7A",
    x"00003E62",
    x"00003E4A",
    x"00003E31",
    x"00003E19",
    x"00003E01",
    x"00003DE9",
    x"00003DD0",
    x"00003DB8",
    x"00003DA0",
    x"00003D88",
    x"00003D70",
    x"00003D58",
    x"00003D40",
    x"00003D28",
    x"00003D10",
    x"00003CF9",
    x"00003CE1",
    x"00003CC9",
    x"00003CB1",
    x"00003C9A",
    x"00003C82",
    x"00003C6A",
    x"00003C53",
    x"00003C3B",
    x"00003C24",
    x"00003C0C",
    x"00003BF5",
    x"00003BDD",
    x"00003BC6",
    x"00003BAF",
    x"00003B97",
    x"00003B80",
    x"00003B69",
    x"00003B52",
    x"00003B3B",
    x"00003B23",
    x"00003B0C",
    x"00003AF5",
    x"00003ADE",
    x"00003AC7",
    x"00003AB0",
    x"00003A99",
    x"00003A83",
    x"00003A6C",
    x"00003A55",
    x"00003A3E",
    x"00003A27",
    x"00003A11",
    x"000039FA",
    x"000039E3",
    x"000039CD",
    x"000039B6",
    x"000039A0",
    x"00003989",
    x"00003973",
    x"0000395C",
    x"00003946",
    x"00003930",
    x"00003919",
    x"00003903",
    x"000038ED",
    x"000038D7",
    x"000038C0",
    x"000038AA",
    x"00003894",
    x"0000387E",
    x"00003868",
    x"00003852",
    x"0000383C",
    x"00003826",
    x"00003810",
    x"000037FA",
    x"000037E4",
    x"000037CF",
    x"000037B9",
    x"000037A3",
    x"0000378D",
    x"00003778",
    x"00003762",
    x"0000374C",
    x"00003737",
    x"00003721",
    x"0000370C",
    x"000036F6",
    x"000036E1",
    x"000036CB",
    x"000036B6",
    x"000036A1",
    x"0000368B",
    x"00003676",
    x"00003661",
    x"0000364C",
    x"00003636",
    x"00003621",
    x"0000360C",
    x"000035F7",
    x"000035E2",
    x"000035CD",
    x"000035B8",
    x"000035A3",
    x"0000358E",
    x"00003579",
    x"00003564",
    x"0000354F",
    x"0000353B",
    x"00003526",
    x"00003511",
    x"000034FC",
    x"000034E8",
    x"000034D3",
    x"000034BE",
    x"000034AA",
    x"00003495",
    x"00003481",
    x"0000346C",
    x"00003458",
    x"00003443",
    x"0000342F",
    x"0000341B",
    x"00003406",
    x"000033F2",
    x"000033DE",
    x"000033C9",
    x"000033B5",
    x"000033A1",
    x"0000338D",
    x"00003379",
    x"00003365",
    x"00003351",
    x"0000333D",
    x"00003329",
    x"00003315",
    x"00003301",
    x"000032ED",
    x"000032D9",
    x"000032C5",
    x"000032B1",
    x"0000329D",
    x"0000328A",
    x"00003276",
    x"00003262",
    x"0000324F",
    x"0000323B",
    x"00003227",
    x"00003214",
    x"00003200",
    x"000031ED",
    x"000031D9",
    x"000031C6",
    x"000031B2",
    x"0000319F",
    x"0000318C",
    x"00003178",
    x"00003165",
    x"00003152",
    x"0000313E",
    x"0000312B",
    x"00003118",
    x"00003105",
    x"000030F2",
    x"000030DF",
    x"000030CB",
    x"000030B8",
    x"000030A5",
    x"00003092",
    x"0000307F",
    x"0000306D",
    x"0000305A",
    x"00003047",
    x"00003034",
    x"00003021",
    x"0000300E",
    x"00002FFC",
    x"00002FE9",
    x"00002FD6",
    x"00002FC3",
    x"00002FB1",
    x"00002F9E",
    x"00002F8C",
    x"00002F79",
    x"00002F66",
    x"00002F54",
    x"00002F42",
    x"00002F2F",
    x"00002F1D",
    x"00002F0A",
    x"00002EF8",
    x"00002EE6",
    x"00002ED3",
    x"00002EC1",
    x"00002EAF",
    x"00002E9D",
    x"00002E8A",
    x"00002E78",
    x"00002E66",
    x"00002E54",
    x"00002E42",
    x"00002E30",
    x"00002E1E",
    x"00002E0C",
    x"00002DFA",
    x"00002DE8",
    x"00002DD6",
    x"00002DC4",
    x"00002DB2",
    x"00002DA0",
    x"00002D8F",
    x"00002D7D",
    x"00002D6B",
    x"00002D59",
    x"00002D48",
    x"00002D36",
    x"00002D24",
    x"00002D13",
    x"00002D01",
    x"00002CEF",
    x"00002CDE",
    x"00002CCC",
    x"00002CBB",
    x"00002CA9",
    x"00002C98",
    x"00002C87",
    x"00002C75",
    x"00002C64",
    x"00002C53",
    x"00002C41",
    x"00002C30",
    x"00002C1F",
    x"00002C0E",
    x"00002BFC",
    x"00002BEB",
    x"00002BDA",
    x"00002BC9",
    x"00002BB8",
    x"00002BA7",
    x"00002B96",
    x"00002B85",
    x"00002B74",
    x"00002B63",
    x"00002B52",
    x"00002B41",
    x"00002B30",
    x"00002B1F",
    x"00002B0E",
    x"00002AFE",
    x"00002AED",
    x"00002ADC",
    x"00002ACB",
    x"00002ABB",
    x"00002AAA",
    x"00002A99",
    x"00002A89",
    x"00002A78",
    x"00002A67",
    x"00002A57",
    x"00002A46",
    x"00002A36",
    x"00002A25",
    x"00002A15",
    x"00002A04",
    x"000029F4",
    x"000029E4",
    x"000029D3",
    x"000029C3",
    x"000029B3",
    x"000029A2",
    x"00002992",
    x"00002982",
    x"00002972",
    x"00002962",
    x"00002951",
    x"00002941",
    x"00002931",
    x"00002921",
    x"00002911",
    x"00002901",
    x"000028F1",
    x"000028E1",
    x"000028D1",
    x"000028C1",
    x"000028B1",
    x"000028A1",
    x"00002892",
    x"00002882",
    x"00002872",
    x"00002862",
    x"00002852",
    x"00002843",
    x"00002833",
    x"00002823",
    x"00002814",
    x"00002804",
    x"000027F4",
    x"000027E5",
    x"000027D5",
    x"000027C6",
    x"000027B6",
    x"000027A7",
    x"00002797",
    x"00002788",
    x"00002778",
    x"00002769",
    x"00002759",
    x"0000274A",
    x"0000273B",
    x"0000272B",
    x"0000271C",
    x"0000270D",
    x"000026FE",
    x"000026EE",
    x"000026DF",
    x"000026D0",
    x"000026C1",
    x"000026B2",
    x"000026A3",
    x"00002694",
    x"00002684",
    x"00002675",
    x"00002666",
    x"00002657",
    x"00002648",
    x"0000263A",
    x"0000262B",
    x"0000261C",
    x"0000260D",
    x"000025FE",
    x"000025EF",
    x"000025E0",
    x"000025D2",
    x"000025C3",
    x"000025B4",
    x"000025A5",
    x"00002597",
    x"00002588",
    x"00002579",
    x"0000256B",
    x"0000255C",
    x"0000254E",
    x"0000253F",
    x"00002530",
    x"00002522",
    x"00002513",
    x"00002505",
    x"000024F6",
    x"000024E8",
    x"000024DA",
    x"000024CB",
    x"000024BD",
    x"000024AF",
    x"000024A0",
    x"00002492",
    x"00002484",
    x"00002475",
    x"00002467",
    x"00002459",
    x"0000244B",
    x"0000243D",
    x"0000242E",
    x"00002420",
    x"00002412",
    x"00002404",
    x"000023F6",
    x"000023E8",
    x"000023DA",
    x"000023CC",
    x"000023BE",
    x"000023B0",
    x"000023A2",
    x"00002394",
    x"00002386",
    x"00002379",
    x"0000236B",
    x"0000235D",
    x"0000234F",
    x"00002341",
    x"00002334",
    x"00002326",
    x"00002318",
    x"0000230A",
    x"000022FD",
    x"000022EF",
    x"000022E1",
    x"000022D4",
    x"000022C6",
    x"000022B9",
    x"000022AB",
    x"0000229E",
    x"00002290",
    x"00002283",
    x"00002275",
    x"00002268",
    x"0000225A",
    x"0000224D",
    x"0000223F",
    x"00002232",
    x"00002225",
    x"00002217",
    x"0000220A",
    x"000021FD",
    x"000021EF",
    x"000021E2",
    x"000021D5",
    x"000021C8",
    x"000021BB",
    x"000021AD",
    x"000021A0",
    x"00002193",
    x"00002186",
    x"00002179",
    x"0000216C",
    x"0000215F",
    x"00002152",
    x"00002145",
    x"00002138",
    x"0000212B",
    x"0000211E",
    x"00002111",
    x"00002104",
    x"000020F7",
    x"000020EA",
    x"000020DE",
    x"000020D1",
    x"000020C4",
    x"000020B7",
    x"000020AA",
    x"0000209E",
    x"00002091",
    x"00002084",
    x"00002077",
    x"0000206B",
    x"0000205E",
    x"00002051",
    x"00002045",
    x"00002038",
    x"0000202C",
    x"0000201F",
    x"00002013",
    x"00002006",
    x"00001FFA",
    x"00001FED",
    x"00001FE1",
    x"00001FD4",
    x"00001FC8",
    x"00001FBB",
    x"00001FAF",
    x"00001FA3",
    x"00001F96",
    x"00001F8A",
    x"00001F7E",
    x"00001F71",
    x"00001F65",
    x"00001F59",
    x"00001F4D",
    x"00001F40",
    x"00001F34",
    x"00001F28",
    x"00001F1C",
    x"00001F10",
    x"00001F04",
    x"00001EF7",
    x"00001EEB",
    x"00001EDF",
    x"00001ED3",
    x"00001EC7",
    x"00001EBB",
    x"00001EAF",
    x"00001EA3",
    x"00001E97",
    x"00001E8B",
    x"00001E7F",
    x"00001E74",
    x"00001E68",
    x"00001E5C",
    x"00001E50",
    x"00001E44",
    x"00001E38",
    x"00001E2C",
    x"00001E21",
    x"00001E15",
    x"00001E09",
    x"00001DFD",
    x"00001DF2",
    x"00001DE6",
    x"00001DDA",
    x"00001DCF",
    x"00001DC3",
    x"00001DB7",
    x"00001DAC",
    x"00001DA0",
    x"00001D95",
    x"00001D89",
    x"00001D7E",
    x"00001D72",
    x"00001D67",
    x"00001D5B",
    x"00001D50",
    x"00001D44",
    x"00001D39",
    x"00001D2D",
    x"00001D22",
    x"00001D17",
    x"00001D0B",
    x"00001D00",
    x"00001CF5",
    x"00001CE9",
    x"00001CDE",
    x"00001CD3",
    x"00001CC8",
    x"00001CBC",
    x"00001CB1",
    x"00001CA6",
    x"00001C9B",
    x"00001C90",
    x"00001C84",
    x"00001C79",
    x"00001C6E",
    x"00001C63",
    x"00001C58",
    x"00001C4D",
    x"00001C42",
    x"00001C37",
    x"00001C2C",
    x"00001C21",
    x"00001C16",
    x"00001C0B",
    x"00001C00",
    x"00001BF5",
    x"00001BEA",
    x"00001BDF",
    x"00001BD4",
    x"00001BCA",
    x"00001BBF",
    x"00001BB4",
    x"00001BA9",
    x"00001B9E",
    x"00001B93",
    x"00001B89",
    x"00001B7E",
    x"00001B73",
    x"00001B68",
    x"00001B5E",
    x"00001B53",
    x"00001B48",
    x"00001B3E",
    x"00001B33",
    x"00001B29",
    x"00001B1E",
    x"00001B13",
    x"00001B09",
    x"00001AFE",
    x"00001AF4",
    x"00001AE9",
    x"00001ADF",
    x"00001AD4",
    x"00001ACA",
    x"00001ABF",
    x"00001AB5",
    x"00001AAA",
    x"00001AA0",
    x"00001A96",
    x"00001A8B",
    x"00001A81",
    x"00001A77",
    x"00001A6C",
    x"00001A62",
    x"00001A58",
    x"00001A4D",
    x"00001A43",
    x"00001A39",
    x"00001A2F",
    x"00001A24",
    x"00001A1A",
    x"00001A10",
    x"00001A06",
    x"000019FC",
    x"000019F1",
    x"000019E7",
    x"000019DD",
    x"000019D3",
    x"000019C9",
    x"000019BF",
    x"000019B5",
    x"000019AB",
    x"000019A1",
    x"00001997",
    x"0000198D",
    x"00001983",
    x"00001979",
    x"0000196F",
    x"00001965",
    x"0000195B",
    x"00001951",
    x"00001947",
    x"0000193E",
    x"00001934",
    x"0000192A",
    x"00001920",
    x"00001916",
    x"0000190C",
    x"00001903",
    x"000018F9",
    x"000018EF",
    x"000018E5",
    x"000018DC",
    x"000018D2",
    x"000018C8",
    x"000018BF",
    x"000018B5",
    x"000018AB",
    x"000018A2",
    x"00001898",
    x"0000188E",
    x"00001885",
    x"0000187B",
    x"00001872",
    x"00001868",
    x"0000185F",
    x"00001855",
    x"0000184C",
    x"00001842",
    x"00001839",
    x"0000182F",
    x"00001826",
    x"0000181C",
    x"00001813",
    x"0000180A",
    x"00001800",
    x"000017F7",
    x"000017ED",
    x"000017E4",
    x"000017DB",
    x"000017D2",
    x"000017C8",
    x"000017BF",
    x"000017B6",
    x"000017AC",
    x"000017A3",
    x"0000179A",
    x"00001791",
    x"00001788",
    x"0000177E",
    x"00001775",
    x"0000176C",
    x"00001763",
    x"0000175A",
    x"00001751",
    x"00001748",
    x"0000173E",
    x"00001735",
    x"0000172C",
    x"00001723",
    x"0000171A",
    x"00001711",
    x"00001708",
    x"000016FF",
    x"000016F6",
    x"000016ED",
    x"000016E4",
    x"000016DB",
    x"000016D2",
    x"000016CA",
    x"000016C1",
    x"000016B8",
    x"000016AF",
    x"000016A6",
    x"0000169D",
    x"00001694",
    x"0000168C",
    x"00001683",
    x"0000167A",
    x"00001671",
    x"00001668",
    x"00001660",
    x"00001657",
    x"0000164E",
    x"00001646",
    x"0000163D",
    x"00001634",
    x"0000162C",
    x"00001623",
    x"0000161A",
    x"00001612",
    x"00001609",
    x"00001600",
    x"000015F8",
    x"000015EF",
    x"000015E7",
    x"000015DE",
    x"000015D6",
    x"000015CD",
    x"000015C5",
    x"000015BC",
    x"000015B4",
    x"000015AB",
    x"000015A3",
    x"0000159A",
    x"00001592",
    x"00001589",
    x"00001581",
    x"00001579",
    x"00001570",
    x"00001568",
    x"0000155F",
    x"00001557",
    x"0000154F",
    x"00001546",
    x"0000153E",
    x"00001536",
    x"0000152E",
    x"00001525",
    x"0000151D",
    x"00001515",
    x"0000150D",
    x"00001504",
    x"000014FC",
    x"000014F4",
    x"000014EC",
    x"000014E4",
    x"000014DB",
    x"000014D3",
    x"000014CB",
    x"000014C3",
    x"000014BB",
    x"000014B3",
    x"000014AB",
    x"000014A3",
    x"0000149B",
    x"00001493",
    x"0000148B",
    x"00001483",
    x"0000147B",
    x"00001473",
    x"0000146B",
    x"00001463",
    x"0000145B",
    x"00001453",
    x"0000144B",
    x"00001443",
    x"0000143B",
    x"00001433",
    x"0000142B",
    x"00001423",
    x"0000141B",
    x"00001414",
    x"0000140C",
    x"00001404",
    x"000013FC",
    x"000013F4",
    x"000013ED",
    x"000013E5",
    x"000013DD",
    x"000013D5",
    x"000013CE",
    x"000013C6",
    x"000013BE",
    x"000013B6",
    x"000013AF",
    x"000013A7",
    x"0000139F",
    x"00001398",
    x"00001390",
    x"00001388",
    x"00001381",
    x"00001379",
    x"00001372",
    x"0000136A",
    x"00001362",
    x"0000135B",
    x"00001353",
    x"0000134C",
    x"00001344",
    x"0000133D",
    x"00001335",
    x"0000132E",
    x"00001326",
    x"0000131F",
    x"00001317",
    x"00001310",
    x"00001308",
    x"00001301",
    x"000012FA",
    x"000012F2",
    x"000012EB",
    x"000012E3",
    x"000012DC",
    x"000012D5",
    x"000012CD",
    x"000012C6",
    x"000012BF",
    x"000012B7",
    x"000012B0",
    x"000012A9",
    x"000012A1",
    x"0000129A",
    x"00001293",
    x"0000128C",
    x"00001284",
    x"0000127D",
    x"00001276",
    x"0000126F",
    x"00001268",
    x"00001260",
    x"00001259",
    x"00001252",
    x"0000124B",
    x"00001244",
    x"0000123D",
    x"00001235",
    x"0000122E",
    x"00001227",
    x"00001220",
    x"00001219",
    x"00001212",
    x"0000120B",
    x"00001204",
    x"000011FD",
    x"000011F6",
    x"000011EF",
    x"000011E8",
    x"000011E1",
    x"000011DA",
    x"000011D3",
    x"000011CC",
    x"000011C5",
    x"000011BE",
    x"000011B7",
    x"000011B0",
    x"000011A9",
    x"000011A2",
    x"0000119C",
    x"00001195",
    x"0000118E",
    x"00001187",
    x"00001180",
    x"00001179",
    x"00001172",
    x"0000116C",
    x"00001165",
    x"0000115E",
    x"00001157",
    x"00001151",
    x"0000114A",
    x"00001143",
    x"0000113C",
    x"00001136",
    x"0000112F",
    x"00001128",
    x"00001121",
    x"0000111B",
    x"00001114",
    x"0000110D",
    x"00001107",
    x"00001100",
    x"000010F9",
    x"000010F3",
    x"000010EC",
    x"000010E6",
    x"000010DF",
    x"000010D8",
    x"000010D2",
    x"000010CB",
    x"000010C5",
    x"000010BE",
    x"000010B8",
    x"000010B1",
    x"000010AB",
    x"000010A4",
    x"0000109E",
    x"00001097",
    x"00001091",
    x"0000108A",
    x"00001084",
    x"0000107D",
    x"00001077",
    x"00001070",
    x"0000106A",
    x"00001064",
    x"0000105D",
    x"00001057",
    x"00001050",
    x"0000104A",
    x"00001044",
    x"0000103D",
    x"00001037",
    x"00001031",
    x"0000102A",
    x"00001024",
    x"0000101E",
    x"00001017",
    x"00001011",
    x"0000100B",
    x"00001005",
    x"00000FFE",
    x"00000FF8",
    x"00000FF2",
    x"00000FEC",
    x"00000FE6",
    x"00000FDF",
    x"00000FD9",
    x"00000FD3",
    x"00000FCD",
    x"00000FC7",
    x"00000FC0",
    x"00000FBA",
    x"00000FB4",
    x"00000FAE",
    x"00000FA8",
    x"00000FA2",
    x"00000F9C",
    x"00000F96",
    x"00000F90",
    x"00000F89",
    x"00000F83",
    x"00000F7D",
    x"00000F77",
    x"00000F71",
    x"00000F6B",
    x"00000F65",
    x"00000F5F",
    x"00000F59",
    x"00000F53",
    x"00000F4D",
    x"00000F47",
    x"00000F41",
    x"00000F3B",
    x"00000F35",
    x"00000F2F",
    x"00000F29",
    x"00000F24",
    x"00000F1E",
    x"00000F18",
    x"00000F12",
    x"00000F0C",
    x"00000F06",
    x"00000F00",
    x"00000EFA",
    x"00000EF5",
    x"00000EEF",
    x"00000EE9",
    x"00000EE3",
    x"00000EDD",
    x"00000ED7",
    x"00000ED2",
    x"00000ECC",
    x"00000EC6",
    x"00000EC0",
    x"00000EBB",
    x"00000EB5",
    x"00000EAF",
    x"00000EA9",
    x"00000EA4",
    x"00000E9E",
    x"00000E98",
    x"00000E93",
    x"00000E8D",
    x"00000E87",
    x"00000E81",
    x"00000E7C",
    x"00000E76",
    x"00000E71",
    x"00000E6B",
    x"00000E65",
    x"00000E60",
    x"00000E5A",
    x"00000E54",
    x"00000E4F",
    x"00000E49",
    x"00000E44",
    x"00000E3E",
    x"00000E39",
    x"00000E33",
    x"00000E2D",
    x"00000E28",
    x"00000E22",
    x"00000E1D",
    x"00000E17",
    x"00000E12",
    x"00000E0C",
    x"00000E07",
    x"00000E01",
    x"00000DFC",
    x"00000DF6",
    x"00000DF1",
    x"00000DEC",
    x"00000DE6",
    x"00000DE1",
    x"00000DDB",
    x"00000DD6",
    x"00000DD1",
    x"00000DCB",
    x"00000DC6",
    x"00000DC0",
    x"00000DBB",
    x"00000DB6",
    x"00000DB0",
    x"00000DAB",
    x"00000DA6",
    x"00000DA0",
    x"00000D9B",
    x"00000D96",
    x"00000D90",
    x"00000D8B",
    x"00000D86",
    x"00000D80",
    x"00000D7B",
    x"00000D76",
    x"00000D71",
    x"00000D6B",
    x"00000D66",
    x"00000D61",
    x"00000D5C",
    x"00000D57",
    x"00000D51",
    x"00000D4C",
    x"00000D47",
    x"00000D42",
    x"00000D3D",
    x"00000D37",
    x"00000D32",
    x"00000D2D",
    x"00000D28",
    x"00000D23",
    x"00000D1E",
    x"00000D19",
    x"00000D13",
    x"00000D0E",
    x"00000D09",
    x"00000D04",
    x"00000CFF",
    x"00000CFA",
    x"00000CF5",
    x"00000CF0",
    x"00000CEB",
    x"00000CE6",
    x"00000CE1",
    x"00000CDC",
    x"00000CD7",
    x"00000CD2",
    x"00000CCD",
    x"00000CC8",
    x"00000CC3",
    x"00000CBE",
    x"00000CB9",
    x"00000CB4",
    x"00000CAF",
    x"00000CAA",
    x"00000CA5",
    x"00000CA0",
    x"00000C9B",
    x"00000C96",
    x"00000C91",
    x"00000C8C",
    x"00000C87",
    x"00000C83",
    x"00000C7E",
    x"00000C79",
    x"00000C74",
    x"00000C6F",
    x"00000C6A",
    x"00000C65",
    x"00000C61",
    x"00000C5C",
    x"00000C57",
    x"00000C52",
    x"00000C4D",
    x"00000C48",
    x"00000C44",
    x"00000C3F",
    x"00000C3A",
    x"00000C35",
    x"00000C31",
    x"00000C2C",
    x"00000C27",
    x"00000C22",
    x"00000C1E",
    x"00000C19",
    x"00000C14",
    x"00000C0F",
    x"00000C0B",
    x"00000C06",
    x"00000C01",
    x"00000BFD",
    x"00000BF8",
    x"00000BF3",
    x"00000BEF",
    x"00000BEA",
    x"00000BE5",
    x"00000BE1",
    x"00000BDC",
    x"00000BD7",
    x"00000BD3",
    x"00000BCE",
    x"00000BCA",
    x"00000BC5",
    x"00000BC0",
    x"00000BBC",
    x"00000BB7",
    x"00000BB3",
    x"00000BAE",
    x"00000BAA",
    x"00000BA5",
    x"00000BA0",
    x"00000B9C",
    x"00000B97",
    x"00000B93",
    x"00000B8E",
    x"00000B8A",
    x"00000B85",
    x"00000B81",
    x"00000B7C",
    x"00000B78",
    x"00000B73",
    x"00000B6F",
    x"00000B6A",
    x"00000B66",
    x"00000B62",
    x"00000B5D",
    x"00000B59",
    x"00000B54",
    x"00000B50",
    x"00000B4B",
    x"00000B47",
    x"00000B43",
    x"00000B3E",
    x"00000B3A",
    x"00000B35",
    x"00000B31",
    x"00000B2D",
    x"00000B28",
    x"00000B24",
    x"00000B20",
    x"00000B1B",
    x"00000B17",
    x"00000B13",
    x"00000B0E",
    x"00000B0A",
    x"00000B06",
    x"00000B01",
    x"00000AFD",
    x"00000AF9",
    x"00000AF4",
    x"00000AF0",
    x"00000AEC",
    x"00000AE8",
    x"00000AE3",
    x"00000ADF",
    x"00000ADB",
    x"00000AD7",
    x"00000AD2",
    x"00000ACE",
    x"00000ACA",
    x"00000AC6",
    x"00000AC2",
    x"00000ABD",
    x"00000AB9",
    x"00000AB5",
    x"00000AB1",
    x"00000AAD",
    x"00000AA8",
    x"00000AA4",
    x"00000AA0",
    x"00000A9C",
    x"00000A98",
    x"00000A94",
    x"00000A90",
    x"00000A8B",
    x"00000A87",
    x"00000A83",
    x"00000A7F",
    x"00000A7B",
    x"00000A77",
    x"00000A73",
    x"00000A6F",
    x"00000A6B",
    x"00000A67",
    x"00000A63",
    x"00000A5F",
    x"00000A5B",
    x"00000A56",
    x"00000A52",
    x"00000A4E",
    x"00000A4A",
    x"00000A46",
    x"00000A42",
    x"00000A3E",
    x"00000A3A",
    x"00000A36",
    x"00000A32",
    x"00000A2E",
    x"00000A2A",
    x"00000A26",
    x"00000A22",
    x"00000A1F",
    x"00000A1B",
    x"00000A17",
    x"00000A13",
    x"00000A0F",
    x"00000A0B",
    x"00000A07",
    x"00000A03",
    x"000009FF",
    x"000009FB",
    x"000009F7",
    x"000009F3",
    x"000009F0",
    x"000009EC",
    x"000009E8",
    x"000009E4",
    x"000009E0",
    x"000009DC",
    x"000009D8",
    x"000009D5",
    x"000009D1",
    x"000009CD",
    x"000009C9",
    x"000009C5",
    x"000009C1",
    x"000009BE",
    x"000009BA",
    x"000009B6",
    x"000009B2",
    x"000009AE",
    x"000009AB",
    x"000009A7",
    x"000009A3",
    x"0000099F",
    x"0000099C",
    x"00000998",
    x"00000994",
    x"00000990",
    x"0000098D",
    x"00000989",
    x"00000985",
    x"00000981",
    x"0000097E",
    x"0000097A",
    x"00000976",
    x"00000973",
    x"0000096F",
    x"0000096B",
    x"00000968",
    x"00000964",
    x"00000960",
    x"0000095D",
    x"00000959",
    x"00000955",
    x"00000952",
    x"0000094E",
    x"0000094A",
    x"00000947",
    x"00000943",
    x"00000940",
    x"0000093C",
    x"00000938",
    x"00000935",
    x"00000931",
    x"0000092E",
    x"0000092A",
    x"00000926",
    x"00000923",
    x"0000091F",
    x"0000091C",
    x"00000918",
    x"00000915",
    x"00000911",
    x"0000090D",
    x"0000090A",
    x"00000906",
    x"00000903",
    x"000008FF",
    x"000008FC",
    x"000008F8",
    x"000008F5",
    x"000008F1",
    x"000008EE",
    x"000008EA",
    x"000008E7",
    x"000008E3",
    x"000008E0",
    x"000008DC",
    x"000008D9",
    x"000008D6",
    x"000008D2",
    x"000008CF",
    x"000008CB",
    x"000008C8",
    x"000008C4",
    x"000008C1",
    x"000008BE",
    x"000008BA",
    x"000008B7",
    x"000008B3",
    x"000008B0",
    x"000008AD",
    x"000008A9",
    x"000008A6",
    x"000008A2",
    x"0000089F",
    x"0000089C",
    x"00000898",
    x"00000895",
    x"00000892",
    x"0000088E",
    x"0000088B",
    x"00000888",
    x"00000884",
    x"00000881",
    x"0000087E",
    x"0000087A",
    x"00000877",
    x"00000874",
    x"00000870",
    x"0000086D",
    x"0000086A",
    x"00000867",
    x"00000863",
    x"00000860",
    x"0000085D",
    x"00000859",
    x"00000856",
    x"00000853",
    x"00000850",
    x"0000084C",
    x"00000849",
    x"00000846",
    x"00000843",
    x"0000083F",
    x"0000083C",
    x"00000839",
    x"00000836",
    x"00000833",
    x"0000082F",
    x"0000082C",
    x"00000829",
    x"00000826",
    x"00000823",
    x"00000820",
    x"0000081C",
    x"00000819",
    x"00000816",
    x"00000813",
    x"00000810",
    x"0000080D",
    x"00000809",
    x"00000806",
    x"00000803",
    x"00000800",
    x"000007FD",
    x"000007FA",
    x"000007F7",
    x"000007F4",
    x"000007F0",
    x"000007ED",
    x"000007EA",
    x"000007E7",
    x"000007E4",
    x"000007E1",
    x"000007DE",
    x"000007DB",
    x"000007D8",
    x"000007D5",
    x"000007D2",
    x"000007CF",
    x"000007CC",
    x"000007C9",
    x"000007C6",
    x"000007C2",
    x"000007BF",
    x"000007BC",
    x"000007B9",
    x"000007B6",
    x"000007B3",
    x"000007B0",
    x"000007AD",
    x"000007AA",
    x"000007A7",
    x"000007A4",
    x"000007A1",
    x"0000079E",
    x"0000079B",
    x"00000798",
    x"00000796",
    x"00000793",
    x"00000790",
    x"0000078D",
    x"0000078A",
    x"00000787",
    x"00000784",
    x"00000781",
    x"0000077E",
    x"0000077B",
    x"00000778",
    x"00000775",
    x"00000772",
    x"0000076F",
    x"0000076C",
    x"0000076A",
    x"00000767",
    x"00000764",
    x"00000761",
    x"0000075E",
    x"0000075B",
    x"00000758",
    x"00000755",
    x"00000753",
    x"00000750",
    x"0000074D",
    x"0000074A",
    x"00000747",
    x"00000744",
    x"00000741",
    x"0000073F",
    x"0000073C",
    x"00000739",
    x"00000736",
    x"00000733",
    x"00000731",
    x"0000072E",
    x"0000072B",
    x"00000728",
    x"00000725",
    x"00000723",
    x"00000720",
    x"0000071D",
    x"0000071A",
    x"00000717",
    x"00000715",
    x"00000712",
    x"0000070F",
    x"0000070C",
    x"0000070A",
    x"00000707",
    x"00000704",
    x"00000701",
    x"000006FF",
    x"000006FC",
    x"000006F9",
    x"000006F7",
    x"000006F4",
    x"000006F1",
    x"000006EE",
    x"000006EC",
    x"000006E9",
    x"000006E6",
    x"000006E4",
    x"000006E1",
    x"000006DE",
    x"000006DC",
    x"000006D9",
    x"000006D6",
    x"000006D4",
    x"000006D1",
    x"000006CE",
    x"000006CC",
    x"000006C9",
    x"000006C6",
    x"000006C4",
    x"000006C1",
    x"000006BE",
    x"000006BC",
    x"000006B9",
    x"000006B6",
    x"000006B4",
    x"000006B1",
    x"000006AF",
    x"000006AC",
    x"000006A9",
    x"000006A7",
    x"000006A4",
    x"000006A2",
    x"0000069F",
    x"0000069C",
    x"0000069A",
    x"00000697",
    x"00000695",
    x"00000692",
    x"00000690",
    x"0000068D",
    x"0000068A",
    x"00000688",
    x"00000685",
    x"00000683",
    x"00000680",
    x"0000067E",
    x"0000067B",
    x"00000679",
    x"00000676",
    x"00000674",
    x"00000671",
    x"0000066F",
    x"0000066C",
    x"0000066A",
    x"00000667",
    x"00000665",
    x"00000662",
    x"00000660",
    x"0000065D",
    x"0000065B",
    x"00000658",
    x"00000656",
    x"00000653",
    x"00000651",
    x"0000064E",
    x"0000064C",
    x"00000649",
    x"00000647",
    x"00000644",
    x"00000642",
    x"0000063F",
    x"0000063D",
    x"0000063B",
    x"00000638",
    x"00000636",
    x"00000633",
    x"00000631",
    x"0000062E",
    x"0000062C",
    x"0000062A",
    x"00000627",
    x"00000625",
    x"00000622",
    x"00000620",
    x"0000061E",
    x"0000061B",
    x"00000619",
    x"00000617",
    x"00000614",
    x"00000612",
    x"0000060F",
    x"0000060D",
    x"0000060B",
    x"00000608",
    x"00000606",
    x"00000604",
    x"00000601",
    x"000005FF",
    x"000005FD",
    x"000005FA",
    x"000005F8",
    x"000005F6",
    x"000005F3",
    x"000005F1",
    x"000005EF",
    x"000005EC",
    x"000005EA",
    x"000005E8",
    x"000005E5",
    x"000005E3",
    x"000005E1",
    x"000005DE",
    x"000005DC",
    x"000005DA",
    x"000005D8",
    x"000005D5",
    x"000005D3",
    x"000005D1",
    x"000005CF",
    x"000005CC",
    x"000005CA",
    x"000005C8",
    x"000005C5",
    x"000005C3",
    x"000005C1",
    x"000005BF",
    x"000005BC",
    x"000005BA",
    x"000005B8",
    x"000005B6",
    x"000005B4",
    x"000005B1",
    x"000005AF",
    x"000005AD",
    x"000005AB",
    x"000005A8",
    x"000005A6",
    x"000005A4",
    x"000005A2",
    x"000005A0",
    x"0000059D",
    x"0000059B",
    x"00000599",
    x"00000597",
    x"00000595",
    x"00000593",
    x"00000590",
    x"0000058E",
    x"0000058C",
    x"0000058A",
    x"00000588",
    x"00000586",
    x"00000583",
    x"00000581",
    x"0000057F",
    x"0000057D",
    x"0000057B",
    x"00000579",
    x"00000577",
    x"00000574",
    x"00000572",
    x"00000570",
    x"0000056E",
    x"0000056C",
    x"0000056A",
    x"00000568",
    x"00000566",
    x"00000563",
    x"00000561",
    x"0000055F",
    x"0000055D",
    x"0000055B",
    x"00000559",
    x"00000557",
    x"00000555",
    x"00000553",
    x"00000551",
    x"0000054F",
    x"0000054C",
    x"0000054A",
    x"00000548",
    x"00000546",
    x"00000544",
    x"00000542",
    x"00000540",
    x"0000053E",
    x"0000053C",
    x"0000053A",
    x"00000538",
    x"00000536",
    x"00000534",
    x"00000532",
    x"00000530",
    x"0000052E",
    x"0000052C",
    x"0000052A",
    x"00000528",
    x"00000526",
    x"00000524",
    x"00000522",
    x"00000520",
    x"0000051E",
    x"0000051C",
    x"0000051A",
    x"00000518",
    x"00000516",
    x"00000514",
    x"00000512",
    x"00000510",
    x"0000050E",
    x"0000050C",
    x"0000050A",
    x"00000508",
    x"00000506",
    x"00000504",
    x"00000502",
    x"00000500",
    x"000004FE",
    x"000004FC",
    x"000004FA",
    x"000004F8",
    x"000004F6",
    x"000004F4",
    x"000004F2",
    x"000004F1",
    x"000004EF",
    x"000004ED",
    x"000004EB",
    x"000004E9",
    x"000004E7",
    x"000004E5",
    x"000004E3",
    x"000004E1",
    x"000004DF",
    x"000004DD",
    x"000004DB",
    x"000004DA",
    x"000004D8",
    x"000004D6",
    x"000004D4",
    x"000004D2",
    x"000004D0",
    x"000004CE",
    x"000004CC",
    x"000004CB",
    x"000004C9",
    x"000004C7",
    x"000004C5",
    x"000004C3",
    x"000004C1",
    x"000004BF",
    x"000004BD",
    x"000004BC",
    x"000004BA",
    x"000004B8",
    x"000004B6",
    x"000004B4",
    x"000004B2",
    x"000004B1",
    x"000004AF",
    x"000004AD",
    x"000004AB",
    x"000004A9",
    x"000004A7",
    x"000004A6",
    x"000004A4",
    x"000004A2",
    x"000004A0",
    x"0000049E",
    x"0000049D",
    x"0000049B",
    x"00000499",
    x"00000497",
    x"00000495",
    x"00000494",
    x"00000492",
    x"00000490",
    x"0000048E",
    x"0000048D",
    x"0000048B",
    x"00000489",
    x"00000487",
    x"00000485",
    x"00000484",
    x"00000482",
    x"00000480",
    x"0000047E",
    x"0000047D",
    x"0000047B",
    x"00000479",
    x"00000477",
    x"00000476",
    x"00000474",
    x"00000472",
    x"00000470",
    x"0000046F",
    x"0000046D",
    x"0000046B",
    x"0000046A",
    x"00000468",
    x"00000466",
    x"00000464",
    x"00000463",
    x"00000461",
    x"0000045F",
    x"0000045E",
    x"0000045C",
    x"0000045A",
    x"00000458",
    x"00000457",
    x"00000455",
    x"00000453",
    x"00000452",
    x"00000450",
    x"0000044E",
    x"0000044D",
    x"0000044B",
    x"00000449",
    x"00000448",
    x"00000446",
    x"00000444",
    x"00000443",
    x"00000441",
    x"0000043F",
    x"0000043E",
    x"0000043C",
    x"0000043A",
    x"00000439",
    x"00000437",
    x"00000435",
    x"00000434",
    x"00000432",
    x"00000430",
    x"0000042F",
    x"0000042D",
    x"0000042C",
    x"0000042A",
    x"00000428",
    x"00000427",
    x"00000425",
    x"00000423",
    x"00000422",
    x"00000420",
    x"0000041F",
    x"0000041D",
    x"0000041B",
    x"0000041A",
    x"00000418",
    x"00000417",
    x"00000415",
    x"00000413",
    x"00000412",
    x"00000410",
    x"0000040F",
    x"0000040D",
    x"0000040B",
    x"0000040A",
    x"00000408",
    x"00000407",
    x"00000405",
    x"00000404",
    x"00000402",
    x"00000400",
    x"000003FF",
    x"000003FD",
    x"000003FC",
    x"000003FA",
    x"000003F9",
    x"000003F7",
    x"000003F6",
    x"000003F4",
    x"000003F2",
    x"000003F1",
    x"000003EF",
    x"000003EE",
    x"000003EC",
    x"000003EB",
    x"000003E9",
    x"000003E8",
    x"000003E6",
    x"000003E5",
    x"000003E3",
    x"000003E2",
    x"000003E0",
    x"000003DF",
    x"000003DD",
    x"000003DC",
    x"000003DA",
    x"000003D9",
    x"000003D7",
    x"000003D6",
    x"000003D4",
    x"000003D3",
    x"000003D1",
    x"000003D0",
    x"000003CE",
    x"000003CD",
    x"000003CB",
    x"000003CA",
    x"000003C8",
    x"000003C7",
    x"000003C5",
    x"000003C4",
    x"000003C2",
    x"000003C1",
    x"000003BF",
    x"000003BE",
    x"000003BC",
    x"000003BB",
    x"000003BA",
    x"000003B8",
    x"000003B7",
    x"000003B5",
    x"000003B4",
    x"000003B2",
    x"000003B1",
    x"000003AF",
    x"000003AE",
    x"000003AD",
    x"000003AB",
    x"000003AA",
    x"000003A8",
    x"000003A7",
    x"000003A5",
    x"000003A4",
    x"000003A3",
    x"000003A1",
    x"000003A0",
    x"0000039E",
    x"0000039D",
    x"0000039B",
    x"0000039A",
    x"00000399",
    x"00000397",
    x"00000396",
    x"00000394",
    x"00000393",
    x"00000392",
    x"00000390",
    x"0000038F",
    x"0000038D",
    x"0000038C",
    x"0000038B",
    x"00000389",
    x"00000388",
    x"00000387",
    x"00000385",
    x"00000384",
    x"00000382",
    x"00000381",
    x"00000380",
    x"0000037E",
    x"0000037D",
    x"0000037C",
    x"0000037A",
    x"00000379",
    x"00000378",
    x"00000376",
    x"00000375",
    x"00000373",
    x"00000372",
    x"00000371",
    x"0000036F",
    x"0000036E",
    x"0000036D",
    x"0000036B",
    x"0000036A",
    x"00000369",
    x"00000367",
    x"00000366",
    x"00000365",
    x"00000363",
    x"00000362",
    x"00000361",
    x"0000035F",
    x"0000035E",
    x"0000035D",
    x"0000035C",
    x"0000035A",
    x"00000359",
    x"00000358",
    x"00000356",
    x"00000355",
    x"00000354",
    x"00000352",
    x"00000351",
    x"00000350",
    x"0000034F",
    x"0000034D",
    x"0000034C",
    x"0000034B",
    x"00000349",
    x"00000348",
    x"00000347",
    x"00000346",
    x"00000344",
    x"00000343",
    x"00000342",
    x"00000340",
    x"0000033F",
    x"0000033E",
    x"0000033D",
    x"0000033B",
    x"0000033A",
    x"00000339",
    x"00000338",
    x"00000336",
    x"00000335",
    x"00000334",
    x"00000333",
    x"00000331",
    x"00000330",
    x"0000032F",
    x"0000032E",
    x"0000032C",
    x"0000032B",
    x"0000032A",
    x"00000329",
    x"00000327",
    x"00000326",
    x"00000325",
    x"00000324",
    x"00000323",
    x"00000321",
    x"00000320",
    x"0000031F",
    x"0000031E",
    x"0000031C",
    x"0000031B",
    x"0000031A",
    x"00000319",
    x"00000318",
    x"00000316",
    x"00000315",
    x"00000314",
    x"00000313",
    x"00000312",
    x"00000310",
    x"0000030F",
    x"0000030E",
    x"0000030D",
    x"0000030C",
    x"0000030A",
    x"00000309",
    x"00000308",
    x"00000307",
    x"00000306",
    x"00000304",
    x"00000303",
    x"00000302",
    x"00000301",
    x"00000300",
    x"000002FF",
    x"000002FD",
    x"000002FC",
    x"000002FB",
    x"000002FA",
    x"000002F9",
    x"000002F8",
    x"000002F6",
    x"000002F5",
    x"000002F4",
    x"000002F3",
    x"000002F2",
    x"000002F1",
    x"000002F0",
    x"000002EE",
    x"000002ED",
    x"000002EC",
    x"000002EB",
    x"000002EA",
    x"000002E9",
    x"000002E8",
    x"000002E6",
    x"000002E5",
    x"000002E4",
    x"000002E3",
    x"000002E2",
    x"000002E1",
    x"000002E0",
    x"000002DF",
    x"000002DD",
    x"000002DC",
    x"000002DB",
    x"000002DA",
    x"000002D9",
    x"000002D8",
    x"000002D7",
    x"000002D6",
    x"000002D5",
    x"000002D3",
    x"000002D2",
    x"000002D1",
    x"000002D0",
    x"000002CF",
    x"000002CE",
    x"000002CD",
    x"000002CC",
    x"000002CB",
    x"000002CA",
    x"000002C8",
    x"000002C7",
    x"000002C6",
    x"000002C5",
    x"000002C4",
    x"000002C3",
    x"000002C2",
    x"000002C1",
    x"000002C0",
    x"000002BF",
    x"000002BE",
    x"000002BD",
    x"000002BC",
    x"000002BA",
    x"000002B9",
    x"000002B8",
    x"000002B7",
    x"000002B6",
    x"000002B5",
    x"000002B4",
    x"000002B3",
    x"000002B2",
    x"000002B1",
    x"000002B0",
    x"000002AF",
    x"000002AE",
    x"000002AD",
    x"000002AC",
    x"000002AB",
    x"000002AA",
    x"000002A9",
    x"000002A8",
    x"000002A7",
    x"000002A5",
    x"000002A4",
    x"000002A3",
    x"000002A2",
    x"000002A1",
    x"000002A0",
    x"0000029F",
    x"0000029E",
    x"0000029D",
    x"0000029C",
    x"0000029B",
    x"0000029A",
    x"00000299",
    x"00000298",
    x"00000297",
    x"00000296",
    x"00000295",
    x"00000294",
    x"00000293",
    x"00000292",
    x"00000291",
    x"00000290",
    x"0000028F",
    x"0000028E",
    x"0000028D",
    x"0000028C",
    x"0000028B",
    x"0000028A",
    x"00000289",
    x"00000288",
    x"00000287",
    x"00000286",
    x"00000285",
    x"00000284",
    x"00000283",
    x"00000282",
    x"00000281",
    x"00000280",
    x"0000027F",
    x"0000027E",
    x"0000027D",
    x"0000027C",
    x"0000027B",
    x"0000027A",
    x"00000279",
    x"00000279",
    x"00000278",
    x"00000277",
    x"00000276",
    x"00000275",
    x"00000274",
    x"00000273",
    x"00000272",
    x"00000271",
    x"00000270",
    x"0000026F",
    x"0000026E",
    x"0000026D",
    x"0000026C",
    x"0000026B",
    x"0000026A",
    x"00000269",
    x"00000268",
    x"00000267",
    x"00000266",
    x"00000266",
    x"00000265",
    x"00000264",
    x"00000263",
    x"00000262",
    x"00000261",
    x"00000260",
    x"0000025F",
    x"0000025E",
    x"0000025D",
    x"0000025C",
    x"0000025B",
    x"0000025A",
    x"00000259",
    x"00000259",
    x"00000258",
    x"00000257",
    x"00000256",
    x"00000255",
    x"00000254",
    x"00000253",
    x"00000252",
    x"00000251",
    x"00000250",
    x"0000024F",
    x"0000024F",
    x"0000024E",
    x"0000024D",
    x"0000024C",
    x"0000024B",
    x"0000024A",
    x"00000249",
    x"00000248",
    x"00000247",
    x"00000246",
    x"00000246",
    x"00000245",
    x"00000244",
    x"00000243",
    x"00000242",
    x"00000241",
    x"00000240",
    x"0000023F",
    x"0000023F",
    x"0000023E",
    x"0000023D",
    x"0000023C",
    x"0000023B",
    x"0000023A",
    x"00000239",
    x"00000238",
    x"00000238",
    x"00000237",
    x"00000236",
    x"00000235",
    x"00000234",
    x"00000233",
    x"00000232",
    x"00000232",
    x"00000231",
    x"00000230",
    x"0000022F",
    x"0000022E",
    x"0000022D",
    x"0000022C",
    x"0000022C",
    x"0000022B",
    x"0000022A",
    x"00000229",
    x"00000228",
    x"00000227",
    x"00000227",
    x"00000226",
    x"00000225",
    x"00000224",
    x"00000223",
    x"00000222",
    x"00000221",
    x"00000221",
    x"00000220",
    x"0000021F",
    x"0000021E",
    x"0000021D",
    x"0000021D",
    x"0000021C",
    x"0000021B",
    x"0000021A",
    x"00000219",
    x"00000218",
    x"00000218",
    x"00000217",
    x"00000216",
    x"00000215",
    x"00000214",
    x"00000214",
    x"00000213",
    x"00000212",
    x"00000211",
    x"00000210",
    x"0000020F",
    x"0000020F",
    x"0000020E",
    x"0000020D",
    x"0000020C",
    x"0000020B",
    x"0000020B",
    x"0000020A",
    x"00000209",
    x"00000208",
    x"00000208",
    x"00000207",
    x"00000206",
    x"00000205",
    x"00000204",
    x"00000204",
    x"00000203",
    x"00000202",
    x"00000201",
    x"00000200",
    x"00000200",
    x"000001FF",
    x"000001FE",
    x"000001FD",
    x"000001FD",
    x"000001FC",
    x"000001FB",
    x"000001FA",
    x"000001F9",
    x"000001F9",
    x"000001F8",
    x"000001F7",
    x"000001F6",
    x"000001F6",
    x"000001F5",
    x"000001F4",
    x"000001F3",
    x"000001F3",
    x"000001F2",
    x"000001F1",
    x"000001F0",
    x"000001EF",
    x"000001EF",
    x"000001EE",
    x"000001ED",
    x"000001EC",
    x"000001EC",
    x"000001EB",
    x"000001EA",
    x"000001E9",
    x"000001E9",
    x"000001E8",
    x"000001E7",
    x"000001E7",
    x"000001E6",
    x"000001E5",
    x"000001E4",
    x"000001E4",
    x"000001E3",
    x"000001E2",
    x"000001E1",
    x"000001E1",
    x"000001E0",
    x"000001DF",
    x"000001DE",
    x"000001DE",
    x"000001DD",
    x"000001DC",
    x"000001DC",
    x"000001DB",
    x"000001DA",
    x"000001D9",
    x"000001D9",
    x"000001D8",
    x"000001D7",
    x"000001D6",
    x"000001D6",
    x"000001D5",
    x"000001D4",
    x"000001D4",
    x"000001D3",
    x"000001D2",
    x"000001D1",
    x"000001D1",
    x"000001D0",
    x"000001CF",
    x"000001CF",
    x"000001CE",
    x"000001CD",
    x"000001CD",
    x"000001CC",
    x"000001CB",
    x"000001CA",
    x"000001CA",
    x"000001C9",
    x"000001C8",
    x"000001C8",
    x"000001C7",
    x"000001C6",
    x"000001C6",
    x"000001C5",
    x"000001C4",
    x"000001C3",
    x"000001C3",
    x"000001C2",
    x"000001C1",
    x"000001C1",
    x"000001C0",
    x"000001BF",
    x"000001BF",
    x"000001BE",
    x"000001BD",
    x"000001BD",
    x"000001BC",
    x"000001BB",
    x"000001BB",
    x"000001BA",
    x"000001B9",
    x"000001B9",
    x"000001B8",
    x"000001B7",
    x"000001B7",
    x"000001B6",
    x"000001B5",
    x"000001B5",
    x"000001B4",
    x"000001B3",
    x"000001B3",
    x"000001B2",
    x"000001B1",
    x"000001B1",
    x"000001B0",
    x"000001AF",
    x"000001AF",
    x"000001AE",
    x"000001AD",
    x"000001AD",
    x"000001AC",
    x"000001AB",
    x"000001AB",
    x"000001AA",
    x"000001A9",
    x"000001A9",
    x"000001A8",
    x"000001A7",
    x"000001A7",
    x"000001A6",
    x"000001A6",
    x"000001A5",
    x"000001A4",
    x"000001A4",
    x"000001A3",
    x"000001A2",
    x"000001A2",
    x"000001A1",
    x"000001A0",
    x"000001A0",
    x"0000019F",
    x"0000019E",
    x"0000019E",
    x"0000019D",
    x"0000019D",
    x"0000019C",
    x"0000019B",
    x"0000019B",
    x"0000019A",
    x"00000199",
    x"00000199",
    x"00000198",
    x"00000198",
    x"00000197",
    x"00000196",
    x"00000196",
    x"00000195",
    x"00000194",
    x"00000194",
    x"00000193",
    x"00000193",
    x"00000192",
    x"00000191",
    x"00000191",
    x"00000190",
    x"00000190",
    x"0000018F",
    x"0000018E",
    x"0000018E",
    x"0000018D",
    x"0000018D",
    x"0000018C",
    x"0000018B",
    x"0000018B",
    x"0000018A",
    x"0000018A",
    x"00000189",
    x"00000188",
    x"00000188",
    x"00000187",
    x"00000187",
    x"00000186",
    x"00000185",
    x"00000185",
    x"00000184",
    x"00000184",
    x"00000183",
    x"00000182",
    x"00000182",
    x"00000181",
    x"00000181",
    x"00000180",
    x"0000017F",
    x"0000017F",
    x"0000017E",
    x"0000017E",
    x"0000017D",
    x"0000017D",
    x"0000017C",
    x"0000017B",
    x"0000017B",
    x"0000017A",
    x"0000017A",
    x"00000179",
    x"00000178",
    x"00000178",
    x"00000177",
    x"00000177",
    x"00000176",
    x"00000176",
    x"00000175",
    x"00000174",
    x"00000174",
    x"00000173",
    x"00000173",
    x"00000172",
    x"00000172",
    x"00000171",
    x"00000171",
    x"00000170",
    x"0000016F",
    x"0000016F",
    x"0000016E",
    x"0000016E",
    x"0000016D",
    x"0000016D",
    x"0000016C",
    x"0000016C",
    x"0000016B",
    x"0000016A",
    x"0000016A",
    x"00000169",
    x"00000169",
    x"00000168",
    x"00000168",
    x"00000167",
    x"00000167",
    x"00000166",
    x"00000165",
    x"00000165",
    x"00000164",
    x"00000164",
    x"00000163",
    x"00000163",
    x"00000162",
    x"00000162",
    x"00000161",
    x"00000161",
    x"00000160",
    x"00000160",
    x"0000015F",
    x"0000015E",
    x"0000015E",
    x"0000015D",
    x"0000015D",
    x"0000015C",
    x"0000015C",
    x"0000015B",
    x"0000015B",
    x"0000015A",
    x"0000015A",
    x"00000159",
    x"00000159",
    x"00000158",
    x"00000158",
    x"00000157",
    x"00000157",
    x"00000156",
    x"00000155",
    x"00000155",
    x"00000154",
    x"00000154",
    x"00000153",
    x"00000153",
    x"00000152",
    x"00000152",
    x"00000151",
    x"00000151",
    x"00000150",
    x"00000150",
    x"0000014F",
    x"0000014F",
    x"0000014E",
    x"0000014E",
    x"0000014D",
    x"0000014D",
    x"0000014C",
    x"0000014C",
    x"0000014B",
    x"0000014B",
    x"0000014A",
    x"0000014A",
    x"00000149",
    x"00000149",
    x"00000148",
    x"00000148",
    x"00000147",
    x"00000147",
    x"00000146",
    x"00000146",
    x"00000145",
    x"00000145",
    x"00000144",
    x"00000144",
    x"00000143",
    x"00000143",
    x"00000142",
    x"00000142",
    x"00000141",
    x"00000141",
    x"00000140",
    x"00000140",
    x"0000013F",
    x"0000013F",
    x"0000013E",
    x"0000013E",
    x"0000013D",
    x"0000013D",
    x"0000013C",
    x"0000013C",
    x"0000013B",
    x"0000013B",
    x"0000013A",
    x"0000013A",
    x"0000013A",
    x"00000139",
    x"00000139",
    x"00000138",
    x"00000138",
    x"00000137",
    x"00000137",
    x"00000136",
    x"00000136",
    x"00000135",
    x"00000135",
    x"00000134",
    x"00000134",
    x"00000133",
    x"00000133",
    x"00000132",
    x"00000132",
    x"00000131",
    x"00000131",
    x"00000131",
    x"00000130",
    x"00000130",
    x"0000012F",
    x"0000012F",
    x"0000012E",
    x"0000012E",
    x"0000012D",
    x"0000012D",
    x"0000012C",
    x"0000012C",
    x"0000012B",
    x"0000012B",
    x"0000012B",
    x"0000012A",
    x"0000012A",
    x"00000129",
    x"00000129",
    x"00000128",
    x"00000128",
    x"00000127",
    x"00000127",
    x"00000126",
    x"00000126",
    x"00000126",
    x"00000125",
    x"00000125",
    x"00000124",
    x"00000124",
    x"00000123",
    x"00000123",
    x"00000122",
    x"00000122",
    x"00000122",
    x"00000121",
    x"00000121",
    x"00000120",
    x"00000120",
    x"0000011F",
    x"0000011F",
    x"0000011F",
    x"0000011E",
    x"0000011E",
    x"0000011D",
    x"0000011D",
    x"0000011C",
    x"0000011C",
    x"0000011B",
    x"0000011B",
    x"0000011B",
    x"0000011A",
    x"0000011A",
    x"00000119",
    x"00000119",
    x"00000118",
    x"00000118",
    x"00000118",
    x"00000117",
    x"00000117",
    x"00000116",
    x"00000116",
    x"00000115",
    x"00000115",
    x"00000115",
    x"00000114",
    x"00000114",
    x"00000113",
    x"00000113",
    x"00000113",
    x"00000112",
    x"00000112",
    x"00000111",
    x"00000111",
    x"00000110",
    x"00000110",
    x"00000110",
    x"0000010F",
    x"0000010F",
    x"0000010E",
    x"0000010E",
    x"0000010E",
    x"0000010D",
    x"0000010D",
    x"0000010C",
    x"0000010C",
    x"0000010B",
    x"0000010B",
    x"0000010B",
    x"0000010A",
    x"0000010A",
    x"00000109",
    x"00000109",
    x"00000109",
    x"00000108",
    x"00000108",
    x"00000107",
    x"00000107",
    x"00000107",
    x"00000106",
    x"00000106",
    x"00000105",
    x"00000105",
    x"00000105",
    x"00000104",
    x"00000104",
    x"00000103",
    x"00000103",
    x"00000103",
    x"00000102",
    x"00000102",
    x"00000101",
    x"00000101",
    x"00000101",
    x"00000100",
    x"00000100",
    x"00000100",
    x"000000FF",
    x"000000FF",
    x"000000FE",
    x"000000FE",
    x"000000FE",
    x"000000FD",
    x"000000FD",
    x"000000FC",
    x"000000FC",
    x"000000FC",
    x"000000FB",
    x"000000FB",
    x"000000FB",
    x"000000FA",
    x"000000FA",
    x"000000F9",
    x"000000F9",
    x"000000F9",
    x"000000F8",
    x"000000F8",
    x"000000F7",
    x"000000F7",
    x"000000F7",
    x"000000F6",
    x"000000F6",
    x"000000F6",
    x"000000F5",
    x"000000F5",
    x"000000F4",
    x"000000F4",
    x"000000F4",
    x"000000F3",
    x"000000F3",
    x"000000F3",
    x"000000F2",
    x"000000F2",
    x"000000F2",
    x"000000F1",
    x"000000F1",
    x"000000F0",
    x"000000F0",
    x"000000F0",
    x"000000EF",
    x"000000EF",
    x"000000EF",
    x"000000EE",
    x"000000EE",
    x"000000ED",
    x"000000ED",
    x"000000ED",
    x"000000EC",
    x"000000EC",
    x"000000EC",
    x"000000EB",
    x"000000EB",
    x"000000EB",
    x"000000EA",
    x"000000EA",
    x"000000EA",
    x"000000E9",
    x"000000E9",
    x"000000E8",
    x"000000E8",
    x"000000E8",
    x"000000E7",
    x"000000E7",
    x"000000E7",
    x"000000E6",
    x"000000E6",
    x"000000E6",
    x"000000E5",
    x"000000E5",
    x"000000E5",
    x"000000E4",
    x"000000E4",
    x"000000E4",
    x"000000E3",
    x"000000E3",
    x"000000E3",
    x"000000E2",
    x"000000E2",
    x"000000E1",
    x"000000E1",
    x"000000E1",
    x"000000E0",
    x"000000E0",
    x"000000E0",
    x"000000DF",
    x"000000DF",
    x"000000DF",
    x"000000DE",
    x"000000DE",
    x"000000DE",
    x"000000DD",
    x"000000DD",
    x"000000DD",
    x"000000DC",
    x"000000DC",
    x"000000DC",
    x"000000DB",
    x"000000DB",
    x"000000DB",
    x"000000DA",
    x"000000DA",
    x"000000DA",
    x"000000D9",
    x"000000D9",
    x"000000D9",
    x"000000D8",
    x"000000D8",
    x"000000D8",
    x"000000D7",
    x"000000D7",
    x"000000D7",
    x"000000D6",
    x"000000D6",
    x"000000D6",
    x"000000D5",
    x"000000D5",
    x"000000D5",
    x"000000D4",
    x"000000D4",
    x"000000D4",
    x"000000D3",
    x"000000D3",
    x"000000D3",
    x"000000D3",
    x"000000D2",
    x"000000D2",
    x"000000D2",
    x"000000D1",
    x"000000D1",
    x"000000D1",
    x"000000D0",
    x"000000D0",
    x"000000D0",
    x"000000CF",
    x"000000CF",
    x"000000CF",
    x"000000CE",
    x"000000CE",
    x"000000CE",
    x"000000CD",
    x"000000CD",
    x"000000CD",
    x"000000CC",
    x"000000CC",
    x"000000CC",
    x"000000CC",
    x"000000CB",
    x"000000CB",
    x"000000CB",
    x"000000CA",
    x"000000CA",
    x"000000CA",
    x"000000C9",
    x"000000C9",
    x"000000C9",
    x"000000C8",
    x"000000C8",
    x"000000C8",
    x"000000C8",
    x"000000C7",
    x"000000C7",
    x"000000C7",
    x"000000C6",
    x"000000C6",
    x"000000C6",
    x"000000C5",
    x"000000C5",
    x"000000C5",
    x"000000C5",
    x"000000C4",
    x"000000C4",
    x"000000C4",
    x"000000C3",
    x"000000C3",
    x"000000C3",
    x"000000C2",
    x"000000C2",
    x"000000C2",
    x"000000C2",
    x"000000C1",
    x"000000C1",
    x"000000C1",
    x"000000C0",
    x"000000C0",
    x"000000C0",
    x"000000C0",
    x"000000BF",
    x"000000BF",
    x"000000BF",
    x"000000BE",
    x"000000BE",
    x"000000BE",
    x"000000BD",
    x"000000BD",
    x"000000BD",
    x"000000BD",
    x"000000BC",
    x"000000BC",
    x"000000BC",
    x"000000BB",
    x"000000BB",
    x"000000BB",
    x"000000BB",
    x"000000BA",
    x"000000BA",
    x"000000BA",
    x"000000B9",
    x"000000B9",
    x"000000B9",
    x"000000B9",
    x"000000B8",
    x"000000B8",
    x"000000B8",
    x"000000B8",
    x"000000B7",
    x"000000B7",
    x"000000B7",
    x"000000B6",
    x"000000B6",
    x"000000B6",
    x"000000B6",
    x"000000B5",
    x"000000B5",
    x"000000B5",
    x"000000B4",
    x"000000B4",
    x"000000B4",
    x"000000B4",
    x"000000B3",
    x"000000B3",
    x"000000B3",
    x"000000B3",
    x"000000B2",
    x"000000B2",
    x"000000B2",
    x"000000B1",
    x"000000B1",
    x"000000B1",
    x"000000B1",
    x"000000B0",
    x"000000B0",
    x"000000B0",
    x"000000B0",
    x"000000AF",
    x"000000AF",
    x"000000AF",
    x"000000AE",
    x"000000AE",
    x"000000AE",
    x"000000AE",
    x"000000AD",
    x"000000AD",
    x"000000AD",
    x"000000AD",
    x"000000AC",
    x"000000AC",
    x"000000AC",
    x"000000AC",
    x"000000AB",
    x"000000AB",
    x"000000AB",
    x"000000AB",
    x"000000AA",
    x"000000AA",
    x"000000AA",
    x"000000AA",
    x"000000A9",
    x"000000A9",
    x"000000A9",
    x"000000A8",
    x"000000A8",
    x"000000A8",
    x"000000A8",
    x"000000A7",
    x"000000A7",
    x"000000A7",
    x"000000A7",
    x"000000A6",
    x"000000A6",
    x"000000A6",
    x"000000A6",
    x"000000A5",
    x"000000A5",
    x"000000A5",
    x"000000A5",
    x"000000A4",
    x"000000A4",
    x"000000A4",
    x"000000A4",
    x"000000A3",
    x"000000A3",
    x"000000A3",
    x"000000A3",
    x"000000A2",
    x"000000A2",
    x"000000A2",
    x"000000A2",
    x"000000A1",
    x"000000A1",
    x"000000A1",
    x"000000A1",
    x"000000A0",
    x"000000A0",
    x"000000A0",
    x"000000A0",
    x"0000009F",
    x"0000009F",
    x"0000009F",
    x"0000009F",
    x"0000009E",
    x"0000009E",
    x"0000009E",
    x"0000009E",
    x"0000009E",
    x"0000009D",
    x"0000009D",
    x"0000009D",
    x"0000009D",
    x"0000009C",
    x"0000009C",
    x"0000009C",
    x"0000009C",
    x"0000009B",
    x"0000009B",
    x"0000009B",
    x"0000009B",
    x"0000009A",
    x"0000009A",
    x"0000009A",
    x"0000009A",
    x"00000099",
    x"00000099",
    x"00000099",
    x"00000099",
    x"00000099",
    x"00000098",
    x"00000098",
    x"00000098",
    x"00000098",
    x"00000097",
    x"00000097",
    x"00000097",
    x"00000097",
    x"00000096",
    x"00000096",
    x"00000096",
    x"00000096",
    x"00000096",
    x"00000095",
    x"00000095",
    x"00000095",
    x"00000095",
    x"00000094",
    x"00000094",
    x"00000094",
    x"00000094",
    x"00000094",
    x"00000093",
    x"00000093",
    x"00000093",
    x"00000093",
    x"00000092",
    x"00000092",
    x"00000092",
    x"00000092",
    x"00000092",
    x"00000091",
    x"00000091",
    x"00000091",
    x"00000091",
    x"00000090",
    x"00000090",
    x"00000090",
    x"00000090",
    x"00000090",
    x"0000008F",
    x"0000008F",
    x"0000008F",
    x"0000008F",
    x"0000008E",
    x"0000008E",
    x"0000008E",
    x"0000008E",
    x"0000008E",
    x"0000008D",
    x"0000008D",
    x"0000008D",
    x"0000008D",
    x"0000008C",
    x"0000008C",
    x"0000008C",
    x"0000008C",
    x"0000008C",
    x"0000008B",
    x"0000008B",
    x"0000008B",
    x"0000008B",
    x"0000008B",
    x"0000008A",
    x"0000008A",
    x"0000008A",
    x"0000008A",
    x"0000008A",
    x"00000089",
    x"00000089",
    x"00000089",
    x"00000089",
    x"00000088",
    x"00000088",
    x"00000088",
    x"00000088",
    x"00000088",
    x"00000087",
    x"00000087",
    x"00000087",
    x"00000087",
    x"00000087",
    x"00000086",
    x"00000086",
    x"00000086",
    x"00000086",
    x"00000086",
    x"00000085",
    x"00000085",
    x"00000085",
    x"00000085",
    x"00000085",
    x"00000084",
    x"00000084",
    x"00000084",
    x"00000084",
    x"00000084",
    x"00000083",
    x"00000083",
    x"00000083",
    x"00000083",
    x"00000083",
    x"00000082",
    x"00000082",
    x"00000082",
    x"00000082",
    x"00000082",
    x"00000081",
    x"00000081",
    x"00000081",
    x"00000081",
    x"00000081",
    x"00000080",
    x"00000080",
    x"00000080",
    x"00000080",
    x"00000080",
    x"0000007F",
    x"0000007F",
    x"0000007F",
    x"0000007F",
    x"0000007F",
    x"0000007E",
    x"0000007E",
    x"0000007E",
    x"0000007E",
    x"0000007E",
    x"0000007D",
    x"0000007D",
    x"0000007D",
    x"0000007D",
    x"0000007D",
    x"0000007D",
    x"0000007C",
    x"0000007C",
    x"0000007C",
    x"0000007C",
    x"0000007C",
    x"0000007B",
    x"0000007B",
    x"0000007B",
    x"0000007B",
    x"0000007B",
    x"0000007A",
    x"0000007A",
    x"0000007A",
    x"0000007A",
    x"0000007A",
    x"0000007A",
    x"00000079",
    x"00000079",
    x"00000079",
    x"00000079",
    x"00000079",
    x"00000078",
    x"00000078",
    x"00000078",
    x"00000078",
    x"00000078",
    x"00000078",
    x"00000077",
    x"00000077",
    x"00000077",
    x"00000077",
    x"00000077",
    x"00000076",
    x"00000076",
    x"00000076",
    x"00000076",
    x"00000076",
    x"00000076",
    x"00000075",
    x"00000075",
    x"00000075",
    x"00000075",
    x"00000075",
    x"00000074",
    x"00000074",
    x"00000074",
    x"00000074",
    x"00000074",
    x"00000074",
    x"00000073",
    x"00000073",
    x"00000073",
    x"00000073",
    x"00000073",
    x"00000073",
    x"00000072",
    x"00000072",
    x"00000072",
    x"00000072",
    x"00000072",
    x"00000071",
    x"00000071",
    x"00000071",
    x"00000071",
    x"00000071",
    x"00000071",
    x"00000070",
    x"00000070",
    x"00000070",
    x"00000070",
    x"00000070",
    x"00000070",
    x"0000006F",
    x"0000006F",
    x"0000006F",
    x"0000006F",
    x"0000006F",
    x"0000006F",
    x"0000006E",
    x"0000006E",
    x"0000006E",
    x"0000006E",
    x"0000006E",
    x"0000006E",
    x"0000006D",
    x"0000006D",
    x"0000006D",
    x"0000006D",
    x"0000006D",
    x"0000006D",
    x"0000006C",
    x"0000006C",
    x"0000006C",
    x"0000006C",
    x"0000006C",
    x"0000006C",
    x"0000006B",
    x"0000006B",
    x"0000006B",
    x"0000006B",
    x"0000006B",
    x"0000006B",
    x"0000006A",
    x"0000006A",
    x"0000006A",
    x"0000006A",
    x"0000006A",
    x"0000006A",
    x"00000069",
    x"00000069",
    x"00000069",
    x"00000069",
    x"00000069",
    x"00000069",
    x"00000068",
    x"00000068",
    x"00000068",
    x"00000068",
    x"00000068",
    x"00000068",
    x"00000068",
    x"00000067",
    x"00000067",
    x"00000067",
    x"00000067",
    x"00000067",
    x"00000067",
    x"00000066",
    x"00000066",
    x"00000066",
    x"00000066",
    x"00000066",
    x"00000066",
    x"00000066",
    x"00000065",
    x"00000065",
    x"00000065",
    x"00000065",
    x"00000065",
    x"00000065",
    x"00000064",
    x"00000064",
    x"00000064",
    x"00000064",
    x"00000064",
    x"00000064",
    x"00000064",
    x"00000063",
    x"00000063",
    x"00000063",
    x"00000063",
    x"00000063",
    x"00000063",
    x"00000062",
    x"00000062",
    x"00000062",
    x"00000062",
    x"00000062",
    x"00000062",
    x"00000062",
    x"00000061",
    x"00000061",
    x"00000061",
    x"00000061",
    x"00000061",
    x"00000061",
    x"00000061",
    x"00000060",
    x"00000060",
    x"00000060",
    x"00000060",
    x"00000060",
    x"00000060",
    x"00000060",
    x"0000005F",
    x"0000005F",
    x"0000005F",
    x"0000005F",
    x"0000005F",
    x"0000005F",
    x"0000005E",
    x"0000005E",
    x"0000005E",
    x"0000005E",
    x"0000005E",
    x"0000005E",
    x"0000005E",
    x"0000005D",
    x"0000005D",
    x"0000005D",
    x"0000005D",
    x"0000005D",
    x"0000005D",
    x"0000005D",
    x"0000005C",
    x"0000005C",
    x"0000005C",
    x"0000005C",
    x"0000005C",
    x"0000005C",
    x"0000005C",
    x"0000005C",
    x"0000005B",
    x"0000005B",
    x"0000005B",
    x"0000005B",
    x"0000005B",
    x"0000005B",
    x"0000005B",
    x"0000005A",
    x"0000005A",
    x"0000005A",
    x"0000005A",
    x"0000005A",
    x"0000005A",
    x"0000005A",
    x"00000059",
    x"00000059",
    x"00000059",
    x"00000059",
    x"00000059",
    x"00000059",
    x"00000059",
    x"00000058",
    x"00000058",
    x"00000058",
    x"00000058",
    x"00000058",
    x"00000058",
    x"00000058",
    x"00000058",
    x"00000057",
    x"00000057",
    x"00000057",
    x"00000057",
    x"00000057",
    x"00000057",
    x"00000057",
    x"00000056",
    x"00000056",
    x"00000056",
    x"00000056",
    x"00000056",
    x"00000056",
    x"00000056",
    x"00000056",
    x"00000055",
    x"00000055",
    x"00000055",
    x"00000055",
    x"00000055",
    x"00000055",
    x"00000055",
    x"00000055",
    x"00000054",
    x"00000054",
    x"00000054",
    x"00000054",
    x"00000054",
    x"00000054",
    x"00000054",
    x"00000054",
    x"00000053",
    x"00000053",
    x"00000053",
    x"00000053",
    x"00000053",
    x"00000053",
    x"00000053",
    x"00000052",
    x"00000052",
    x"00000052",
    x"00000052",
    x"00000052",
    x"00000052",
    x"00000052",
    x"00000052",
    x"00000051",
    x"00000051",
    x"00000051",
    x"00000051",
    x"00000051",
    x"00000051",
    x"00000051",
    x"00000051",
    x"00000050",
    x"00000050",
    x"00000050",
    x"00000050",
    x"00000050",
    x"00000050",
    x"00000050",
    x"00000050",
    x"00000050",
    x"0000004F",
    x"0000004F",
    x"0000004F",
    x"0000004F",
    x"0000004F",
    x"0000004F",
    x"0000004F",
    x"0000004F",
    x"0000004E",
    x"0000004E",
    x"0000004E",
    x"0000004E",
    x"0000004E",
    x"0000004E",
    x"0000004E",
    x"0000004E",
    x"0000004D",
    x"0000004D",
    x"0000004D",
    x"0000004D",
    x"0000004D",
    x"0000004D",
    x"0000004D",
    x"0000004D",
    x"0000004D",
    x"0000004C",
    x"0000004C",
    x"0000004C",
    x"0000004C",
    x"0000004C",
    x"0000004C",
    x"0000004C",
    x"0000004C",
    x"0000004C",
    x"0000004B",
    x"0000004B",
    x"0000004B",
    x"0000004B",
    x"0000004B",
    x"0000004B",
    x"0000004B",
    x"0000004B",
    x"0000004A",
    x"0000004A",
    x"0000004A",
    x"0000004A",
    x"0000004A",
    x"0000004A",
    x"0000004A",
    x"0000004A",
    x"0000004A",
    x"00000049",
    x"00000049",
    x"00000049",
    x"00000049",
    x"00000049",
    x"00000049",
    x"00000049",
    x"00000049",
    x"00000049",
    x"00000048",
    x"00000048",
    x"00000048",
    x"00000048",
    x"00000048",
    x"00000048",
    x"00000048",
    x"00000048",
    x"00000048",
    x"00000047",
    x"00000047",
    x"00000047",
    x"00000047",
    x"00000047",
    x"00000047",
    x"00000047",
    x"00000047",
    x"00000047",
    x"00000046",
    x"00000046",
    x"00000046",
    x"00000046",
    x"00000046",
    x"00000046",
    x"00000046",
    x"00000046",
    x"00000046",
    x"00000046",
    x"00000045",
    x"00000045",
    x"00000045",
    x"00000045",
    x"00000045",
    x"00000045",
    x"00000045",
    x"00000045",
    x"00000045",
    x"00000044",
    x"00000044",
    x"00000044",
    x"00000044",
    x"00000044",
    x"00000044",
    x"00000044",
    x"00000044",
    x"00000044",
    x"00000044",
    x"00000043",
    x"00000043",
    x"00000043",
    x"00000043",
    x"00000043",
    x"00000043",
    x"00000043",
    x"00000043",
    x"00000043",
    x"00000043",
    x"00000042",
    x"00000042",
    x"00000042",
    x"00000042",
    x"00000042",
    x"00000042",
    x"00000042",
    x"00000042",
    x"00000042",
    x"00000042",
    x"00000041",
    x"00000041",
    x"00000041",
    x"00000041",
    x"00000041",
    x"00000041",
    x"00000041",
    x"00000041",
    x"00000041",
    x"00000041",
    x"00000040",
    x"00000040",
    x"00000040",
    x"00000040",
    x"00000040",
    x"00000040",
    x"00000040",
    x"00000040",
    x"00000040",
    x"00000040",
    x"0000003F",
    x"0000003F",
    x"0000003F",
    x"0000003F",
    x"0000003F",
    x"0000003F",
    x"0000003F",
    x"0000003F",
    x"0000003F",
    x"0000003F",
    x"0000003E",
    x"0000003E",
    x"0000003E",
    x"0000003E",
    x"0000003E",
    x"0000003E",
    x"0000003E",
    x"0000003E",
    x"0000003E",
    x"0000003E",
    x"0000003E",
    x"0000003D",
    x"0000003D",
    x"0000003D",
    x"0000003D",
    x"0000003D",
    x"0000003D",
    x"0000003D",
    x"0000003D",
    x"0000003D",
    x"0000003D",
    x"0000003D",
    x"0000003C",
    x"0000003C",
    x"0000003C",
    x"0000003C",
    x"0000003C",
    x"0000003C",
    x"0000003C",
    x"0000003C",
    x"0000003C",
    x"0000003C",
    x"0000003C",
    x"0000003B",
    x"0000003B",
    x"0000003B",
    x"0000003B",
    x"0000003B",
    x"0000003B",
    x"0000003B",
    x"0000003B",
    x"0000003B",
    x"0000003B",
    x"0000003B",
    x"0000003A",
    x"0000003A",
    x"0000003A",
    x"0000003A",
    x"0000003A",
    x"0000003A",
    x"0000003A",
    x"0000003A",
    x"0000003A",
    x"0000003A",
    x"0000003A",
    x"00000039",
    x"00000039",
    x"00000039",
    x"00000039",
    x"00000039",
    x"00000039",
    x"00000039",
    x"00000039",
    x"00000039",
    x"00000039",
    x"00000039",
    x"00000038",
    x"00000038",
    x"00000038",
    x"00000038",
    x"00000038",
    x"00000038",
    x"00000038",
    x"00000038",
    x"00000038",
    x"00000038",
    x"00000038",
    x"00000038",
    x"00000037",
    x"00000037",
    x"00000037",
    x"00000037",
    x"00000037",
    x"00000037",
    x"00000037",
    x"00000037",
    x"00000037",
    x"00000037",
    x"00000037",
    x"00000037",
    x"00000036",
    x"00000036",
    x"00000036",
    x"00000036",
    x"00000036",
    x"00000036",
    x"00000036",
    x"00000036",
    x"00000036",
    x"00000036",
    x"00000036",
    x"00000036",
    x"00000035",
    x"00000035",
    x"00000035",
    x"00000035",
    x"00000035",
    x"00000035",
    x"00000035",
    x"00000035",
    x"00000035",
    x"00000035",
    x"00000035",
    x"00000035",
    x"00000035",
    x"00000034",
    x"00000034",
    x"00000034",
    x"00000034",
    x"00000034",
    x"00000034",
    x"00000034",
    x"00000034",
    x"00000034",
    x"00000034",
    x"00000034",
    x"00000034",
    x"00000033",
    x"00000033",
    x"00000033",
    x"00000033",
    x"00000033",
    x"00000033",
    x"00000033",
    x"00000033",
    x"00000033",
    x"00000033",
    x"00000033",
    x"00000033",
    x"00000033",
    x"00000032",
    x"00000032",
    x"00000032",
    x"00000032",
    x"00000032",
    x"00000032",
    x"00000032",
    x"00000032",
    x"00000032",
    x"00000032",
    x"00000032",
    x"00000032",
    x"00000032",
    x"00000031",
    x"00000031",
    x"00000031",
    x"00000031",
    x"00000031",
    x"00000031",
    x"00000031",
    x"00000031",
    x"00000031",
    x"00000031",
    x"00000031",
    x"00000031",
    x"00000031",
    x"00000031",
    x"00000030",
    x"00000030",
    x"00000030",
    x"00000030",
    x"00000030",
    x"00000030",
    x"00000030",
    x"00000030",
    x"00000030",
    x"00000030",
    x"00000030",
    x"00000030",
    x"00000030",
    x"0000002F",
    x"0000002F",
    x"0000002F",
    x"0000002F",
    x"0000002F",
    x"0000002F",
    x"0000002F",
    x"0000002F",
    x"0000002F",
    x"0000002F",
    x"0000002F",
    x"0000002F",
    x"0000002F",
    x"0000002F",
    x"0000002E",
    x"0000002E",
    x"0000002E",
    x"0000002E",
    x"0000002E",
    x"0000002E",
    x"0000002E",
    x"0000002E",
    x"0000002E",
    x"0000002E",
    x"0000002E",
    x"0000002E",
    x"0000002E",
    x"0000002E",
    x"0000002D",
    x"0000002D",
    x"0000002D",
    x"0000002D",
    x"0000002D",
    x"0000002D",
    x"0000002D",
    x"0000002D",
    x"0000002D",
    x"0000002D",
    x"0000002D",
    x"0000002D",
    x"0000002D",
    x"0000002D",
    x"0000002D",
    x"0000002C",
    x"0000002C",
    x"0000002C",
    x"0000002C",
    x"0000002C",
    x"0000002C",
    x"0000002C",
    x"0000002C",
    x"0000002C",
    x"0000002C",
    x"0000002C",
    x"0000002C",
    x"0000002C",
    x"0000002C",
    x"0000002C",
    x"0000002B",
    x"0000002B",
    x"0000002B",
    x"0000002B",
    x"0000002B",
    x"0000002B",
    x"0000002B",
    x"0000002B",
    x"0000002B",
    x"0000002B",
    x"0000002B",
    x"0000002B",
    x"0000002B",
    x"0000002B",
    x"0000002B",
    x"0000002A",
    x"0000002A",
    x"0000002A",
    x"0000002A",
    x"0000002A",
    x"0000002A",
    x"0000002A",
    x"0000002A",
    x"0000002A",
    x"0000002A",
    x"0000002A",
    x"0000002A",
    x"0000002A",
    x"0000002A",
    x"0000002A",
    x"0000002A",
    x"00000029",
    x"00000029",
    x"00000029",
    x"00000029",
    x"00000029",
    x"00000029",
    x"00000029",
    x"00000029",
    x"00000029",
    x"00000029",
    x"00000029",
    x"00000029",
    x"00000029",
    x"00000029",
    x"00000029",
    x"00000029",
    x"00000028",
    x"00000028",
    x"00000028",
    x"00000028",
    x"00000028",
    x"00000028",
    x"00000028",
    x"00000028",
    x"00000028",
    x"00000028",
    x"00000028",
    x"00000028",
    x"00000028",
    x"00000028",
    x"00000028",
    x"00000028",
    x"00000027",
    x"00000027",
    x"00000027",
    x"00000027",
    x"00000027",
    x"00000027",
    x"00000027",
    x"00000027",
    x"00000027",
    x"00000027",
    x"00000027",
    x"00000027",
    x"00000027",
    x"00000027",
    x"00000027",
    x"00000027",
    x"00000027",
    x"00000026",
    x"00000026",
    x"00000026",
    x"00000026",
    x"00000026",
    x"00000026",
    x"00000026",
    x"00000026",
    x"00000026",
    x"00000026",
    x"00000026",
    x"00000026",
    x"00000026",
    x"00000026",
    x"00000026",
    x"00000026",
    x"00000026",
    x"00000025",
    x"00000025",
    x"00000025",
    x"00000025",
    x"00000025",
    x"00000025",
    x"00000025",
    x"00000025",
    x"00000025",
    x"00000025",
    x"00000025",
    x"00000025",
    x"00000025",
    x"00000025",
    x"00000025",
    x"00000025",
    x"00000025",
    x"00000025",
    x"00000024",
    x"00000024",
    x"00000024",
    x"00000024",
    x"00000024",
    x"00000024",
    x"00000024",
    x"00000024",
    x"00000024",
    x"00000024",
    x"00000024",
    x"00000024",
    x"00000024",
    x"00000024",
    x"00000024",
    x"00000024",
    x"00000024",
    x"00000024",
    x"00000023",
    x"00000023",
    x"00000023",
    x"00000023",
    x"00000023",
    x"00000023",
    x"00000023",
    x"00000023",
    x"00000023",
    x"00000023",
    x"00000023",
    x"00000023",
    x"00000023",
    x"00000023",
    x"00000023",
    x"00000023",
    x"00000023",
    x"00000023",
    x"00000023",
    x"00000022",
    x"00000022",
    x"00000022",
    x"00000022",
    x"00000022",
    x"00000022",
    x"00000022",
    x"00000022",
    x"00000022",
    x"00000022",
    x"00000022",
    x"00000022",
    x"00000022",
    x"00000022",
    x"00000022",
    x"00000022",
    x"00000022",
    x"00000022",
    x"00000022",
    x"00000021",
    x"00000021",
    x"00000021",
    x"00000021",
    x"00000021",
    x"00000021",
    x"00000021",
    x"00000021",
    x"00000021",
    x"00000021",
    x"00000021",
    x"00000021",
    x"00000021",
    x"00000021",
    x"00000021",
    x"00000021",
    x"00000021",
    x"00000021",
    x"00000021",
    x"00000021",
    x"00000020",
    x"00000020",
    x"00000020",
    x"00000020",
    x"00000020",
    x"00000020",
    x"00000020",
    x"00000020",
    x"00000020",
    x"00000020",
    x"00000020",
    x"00000020",
    x"00000020",
    x"00000020",
    x"00000020",
    x"00000020",
    x"00000020",
    x"00000020",
    x"00000020",
    x"00000020",
    x"0000001F",
    x"0000001F",
    x"0000001F",
    x"0000001F",
    x"0000001F",
    x"0000001F",
    x"0000001F",
    x"0000001F",
    x"0000001F",
    x"0000001F",
    x"0000001F",
    x"0000001F",
    x"0000001F",
    x"0000001F",
    x"0000001F",
    x"0000001F",
    x"0000001F",
    x"0000001F",
    x"0000001F",
    x"0000001F",
    x"0000001F",
    x"0000001F",
    x"0000001E",
    x"0000001E",
    x"0000001E",
    x"0000001E",
    x"0000001E",
    x"0000001E",
    x"0000001E",
    x"0000001E",
    x"0000001E",
    x"0000001E",
    x"0000001E",
    x"0000001E",
    x"0000001E",
    x"0000001E",
    x"0000001E",
    x"0000001E",
    x"0000001E",
    x"0000001E",
    x"0000001E",
    x"0000001E",
    x"0000001E",
    x"0000001D",
    x"0000001D",
    x"0000001D",
    x"0000001D",
    x"0000001D",
    x"0000001D",
    x"0000001D",
    x"0000001D",
    x"0000001D",
    x"0000001D",
    x"0000001D",
    x"0000001D",
    x"0000001D",
    x"0000001D",
    x"0000001D",
    x"0000001D",
    x"0000001D",
    x"0000001D",
    x"0000001D",
    x"0000001D",
    x"0000001D",
    x"0000001D",
    x"0000001D",
    x"0000001C",
    x"0000001C",
    x"0000001C",
    x"0000001C",
    x"0000001C",
    x"0000001C",
    x"0000001C",
    x"0000001C",
    x"0000001C",
    x"0000001C",
    x"0000001C",
    x"0000001C",
    x"0000001C",
    x"0000001C",
    x"0000001C",
    x"0000001C",
    x"0000001C",
    x"0000001C",
    x"0000001C",
    x"0000001C",
    x"0000001C",
    x"0000001C",
    x"0000001C",
    x"0000001B",
    x"0000001B",
    x"0000001B",
    x"0000001B",
    x"0000001B",
    x"0000001B",
    x"0000001B",
    x"0000001B",
    x"0000001B",
    x"0000001B",
    x"0000001B",
    x"0000001B",
    x"0000001B",
    x"0000001B",
    x"0000001B",
    x"0000001B",
    x"0000001B",
    x"0000001B",
    x"0000001B",
    x"0000001B",
    x"0000001B",
    x"0000001B",
    x"0000001B"
  );

begin

  p_mem_read : process (clk) begin
    if rising_edge(clk) then
      data_out <= mem(to_integer(unsigned(address)));
    end if;
  end process;

end architecture;
