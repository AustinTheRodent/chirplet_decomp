
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sine_rom is
  port
  (
    clk       : in  std_logic;
    address   : in  std_logic_vector(13 downto 0);
    data_out  : out std_logic_vector(31 downto 0)
  );
end entity;

architecture rtl of sine_rom is

  constant C_DATA_WIDTH  : integer := 32;
  constant C_ADDR_WIDTH  : integer := 14;

  constant RAM_DEPTH :integer := 2**C_ADDR_WIDTH;

  type RAM is array (integer range <>) of std_logic_vector (C_DATA_WIDTH-1 downto 0);
  signal mem : RAM (0 to RAM_DEPTH-1) :=
  (
    x"00000000",
    x"38C90FDB",
    x"39490FDB",
    x"3996CBE4",
    x"39C90FDA",
    x"39FB53D1",
    x"3A16CBE3",
    x"3A2FEDDE",
    x"3A490FD9",
    x"3A6231D4",
    x"3A7B53CF",
    x"3A8A3AE5",
    x"3A96CBE2",
    x"3AA35CDF",
    x"3AAFEDDC",
    x"3ABC7ED9",
    x"3AC90FD5",
    x"3AD5A0D2",
    x"3AE231CF",
    x"3AEEC2CB",
    x"3AFB53C7",
    x"3B03F262",
    x"3B0A3AE0",
    x"3B10835D",
    x"3B16CBDB",
    x"3B1D1459",
    x"3B235CD7",
    x"3B29A554",
    x"3B2FEDD1",
    x"3B36364F",
    x"3B3C7ECC",
    x"3B42C749",
    x"3B490FC6",
    x"3B4F5843",
    x"3B55A0C0",
    x"3B5BE93C",
    x"3B6231B9",
    x"3B687A35",
    x"3B6EC2B1",
    x"3B750B2D",
    x"3B7B53A9",
    x"3B80CE12",
    x"3B83F250",
    x"3B87168E",
    x"3B8A3ACB",
    x"3B8D5F09",
    x"3B908346",
    x"3B93A784",
    x"3B96CBC1",
    x"3B99EFFE",
    x"3B9D143B",
    x"3BA03878",
    x"3BA35CB5",
    x"3BA680F2",
    x"3BA9A52F",
    x"3BACC96B",
    x"3BAFEDA8",
    x"3BB311E4",
    x"3BB63621",
    x"3BB95A5D",
    x"3BBC7E99",
    x"3BBFA2D5",
    x"3BC2C711",
    x"3BC5EB4C",
    x"3BC90F88",
    x"3BCC33C3",
    x"3BCF57FF",
    x"3BD27C3A",
    x"3BD5A075",
    x"3BD8C4B0",
    x"3BDBE8EB",
    x"3BDF0D26",
    x"3BE23160",
    x"3BE5559B",
    x"3BE879D5",
    x"3BEB9E0F",
    x"3BEEC249",
    x"3BF1E683",
    x"3BF50ABD",
    x"3BF82EF6",
    x"3BFB5330",
    x"3BFE7769",
    x"3C00CDD1",
    x"3C025FEE",
    x"3C03F20A",
    x"3C058426",
    x"3C071643",
    x"3C08A85F",
    x"3C0A3A7B",
    x"3C0BCC97",
    x"3C0D5EB3",
    x"3C0EF0CF",
    x"3C1082EA",
    x"3C121506",
    x"3C13A722",
    x"3C15393D",
    x"3C16CB58",
    x"3C185D74",
    x"3C19EF8F",
    x"3C1B81AA",
    x"3C1D13C5",
    x"3C1EA5E0",
    x"3C2037FB",
    x"3C21CA16",
    x"3C235C30",
    x"3C24EE4B",
    x"3C268065",
    x"3C281280",
    x"3C29A49A",
    x"3C2B36B4",
    x"3C2CC8CE",
    x"3C2E5AE8",
    x"3C2FED02",
    x"3C317F1B",
    x"3C331135",
    x"3C34A34F",
    x"3C363568",
    x"3C37C781",
    x"3C39599A",
    x"3C3AEBB4",
    x"3C3C7DCC",
    x"3C3E0FE5",
    x"3C3FA1FE",
    x"3C413417",
    x"3C42C62F",
    x"3C445847",
    x"3C45EA60",
    x"3C477C78",
    x"3C490E90",
    x"3C4AA0A8",
    x"3C4C32C0",
    x"3C4DC4D7",
    x"3C4F56EF",
    x"3C50E906",
    x"3C527B1D",
    x"3C540D35",
    x"3C559F4C",
    x"3C573162",
    x"3C58C379",
    x"3C5A5590",
    x"3C5BE7A6",
    x"3C5D79BD",
    x"3C5F0BD3",
    x"3C609DE9",
    x"3C622FFF",
    x"3C63C215",
    x"3C65542B",
    x"3C66E640",
    x"3C687856",
    x"3C6A0A6B",
    x"3C6B9C80",
    x"3C6D2E95",
    x"3C6EC0AA",
    x"3C7052BF",
    x"3C71E4D3",
    x"3C7376E7",
    x"3C7508FC",
    x"3C769B10",
    x"3C782D24",
    x"3C79BF38",
    x"3C7B514B",
    x"3C7CE35F",
    x"3C7E7572",
    x"3C8003C3",
    x"3C80CCCC",
    x"3C8195D6",
    x"3C825EDF",
    x"3C8327E8",
    x"3C83F0F2",
    x"3C84B9FB",
    x"3C858304",
    x"3C864C0D",
    x"3C871516",
    x"3C87DE1E",
    x"3C88A727",
    x"3C897030",
    x"3C8A3938",
    x"3C8B0241",
    x"3C8BCB49",
    x"3C8C9452",
    x"3C8D5D5A",
    x"3C8E2662",
    x"3C8EEF6A",
    x"3C8FB872",
    x"3C90817A",
    x"3C914A82",
    x"3C921389",
    x"3C92DC91",
    x"3C93A599",
    x"3C946EA0",
    x"3C9537A7",
    x"3C9600AF",
    x"3C96C9B6",
    x"3C9792BD",
    x"3C985BC4",
    x"3C9924CB",
    x"3C99EDD2",
    x"3C9AB6D8",
    x"3C9B7FDF",
    x"3C9C48E6",
    x"3C9D11EC",
    x"3C9DDAF2",
    x"3C9EA3F9",
    x"3C9F6CFF",
    x"3CA03605",
    x"3CA0FF0B",
    x"3CA1C811",
    x"3CA29116",
    x"3CA35A1C",
    x"3CA42322",
    x"3CA4EC27",
    x"3CA5B52C",
    x"3CA67E32",
    x"3CA74737",
    x"3CA8103C",
    x"3CA8D941",
    x"3CA9A246",
    x"3CAA6B4B",
    x"3CAB344F",
    x"3CABFD54",
    x"3CACC658",
    x"3CAD8F5D",
    x"3CAE5861",
    x"3CAF2165",
    x"3CAFEA69",
    x"3CB0B36D",
    x"3CB17C71",
    x"3CB24575",
    x"3CB30E78",
    x"3CB3D77C",
    x"3CB4A07F",
    x"3CB56982",
    x"3CB63286",
    x"3CB6FB89",
    x"3CB7C48C",
    x"3CB88D8E",
    x"3CB95691",
    x"3CBA1F94",
    x"3CBAE896",
    x"3CBBB199",
    x"3CBC7A9B",
    x"3CBD439D",
    x"3CBE0C9F",
    x"3CBED5A1",
    x"3CBF9EA3",
    x"3CC067A5",
    x"3CC130A6",
    x"3CC1F9A8",
    x"3CC2C2A9",
    x"3CC38BAA",
    x"3CC454AB",
    x"3CC51DAC",
    x"3CC5E6AD",
    x"3CC6AFAE",
    x"3CC778AF",
    x"3CC841AF",
    x"3CC90AB0",
    x"3CC9D3B0",
    x"3CCA9CB0",
    x"3CCB65B0",
    x"3CCC2EB0",
    x"3CCCF7B0",
    x"3CCDC0B0",
    x"3CCE89AF",
    x"3CCF52AF",
    x"3CD01BAE",
    x"3CD0E4AD",
    x"3CD1ADAC",
    x"3CD276AB",
    x"3CD33FAA",
    x"3CD408A9",
    x"3CD4D1A7",
    x"3CD59AA6",
    x"3CD663A4",
    x"3CD72CA2",
    x"3CD7F5A0",
    x"3CD8BE9E",
    x"3CD9879C",
    x"3CDA5099",
    x"3CDB1997",
    x"3CDBE294",
    x"3CDCAB91",
    x"3CDD748F",
    x"3CDE3D8C",
    x"3CDF0688",
    x"3CDFCF85",
    x"3CE09882",
    x"3CE1617E",
    x"3CE22A7A",
    x"3CE2F377",
    x"3CE3BC73",
    x"3CE4856E",
    x"3CE54E6A",
    x"3CE61766",
    x"3CE6E061",
    x"3CE7A95D",
    x"3CE87258",
    x"3CE93B53",
    x"3CEA044E",
    x"3CEACD49",
    x"3CEB9643",
    x"3CEC5F3E",
    x"3CED2838",
    x"3CEDF132",
    x"3CEEBA2C",
    x"3CEF8326",
    x"3CF04C20",
    x"3CF1151A",
    x"3CF1DE13",
    x"3CF2A70D",
    x"3CF37006",
    x"3CF438FF",
    x"3CF501F8",
    x"3CF5CAF0",
    x"3CF693E9",
    x"3CF75CE2",
    x"3CF825DA",
    x"3CF8EED2",
    x"3CF9B7CA",
    x"3CFA80C2",
    x"3CFB49BA",
    x"3CFC12B1",
    x"3CFCDBA9",
    x"3CFDA4A0",
    x"3CFE6D97",
    x"3CFF368E",
    x"3CFFFF85",
    x"3D00643E",
    x"3D00C8B9",
    x"3D012D34",
    x"3D0191AF",
    x"3D01F62A",
    x"3D025AA5",
    x"3D02BF20",
    x"3D03239B",
    x"3D038815",
    x"3D03EC90",
    x"3D04510B",
    x"3D04B585",
    x"3D0519FF",
    x"3D057E7A",
    x"3D05E2F4",
    x"3D06476E",
    x"3D06ABE8",
    x"3D071062",
    x"3D0774DC",
    x"3D07D956",
    x"3D083DCF",
    x"3D08A249",
    x"3D0906C3",
    x"3D096B3C",
    x"3D09CFB6",
    x"3D0A342F",
    x"3D0A98A8",
    x"3D0AFD21",
    x"3D0B619A",
    x"3D0BC613",
    x"3D0C2A8C",
    x"3D0C8F05",
    x"3D0CF37E",
    x"3D0D57F6",
    x"3D0DBC6F",
    x"3D0E20E7",
    x"3D0E8560",
    x"3D0EE9D8",
    x"3D0F4E50",
    x"3D0FB2C8",
    x"3D101740",
    x"3D107BB8",
    x"3D10E030",
    x"3D1144A8",
    x"3D11A920",
    x"3D120D97",
    x"3D12720F",
    x"3D12D686",
    x"3D133AFE",
    x"3D139F75",
    x"3D1403EC",
    x"3D146863",
    x"3D14CCDA",
    x"3D153151",
    x"3D1595C8",
    x"3D15FA3F",
    x"3D165EB5",
    x"3D16C32C",
    x"3D1727A2",
    x"3D178C18",
    x"3D17F08F",
    x"3D185505",
    x"3D18B97B",
    x"3D191DF1",
    x"3D198267",
    x"3D19E6DD",
    x"3D1A4B52",
    x"3D1AAFC8",
    x"3D1B143D",
    x"3D1B78B3",
    x"3D1BDD28",
    x"3D1C419D",
    x"3D1CA613",
    x"3D1D0A88",
    x"3D1D6EFD",
    x"3D1DD372",
    x"3D1E37E6",
    x"3D1E9C5B",
    x"3D1F00D0",
    x"3D1F6544",
    x"3D1FC9B8",
    x"3D202E2D",
    x"3D2092A1",
    x"3D20F715",
    x"3D215B89",
    x"3D21BFFD",
    x"3D222471",
    x"3D2288E4",
    x"3D22ED58",
    x"3D2351CB",
    x"3D23B63F",
    x"3D241AB2",
    x"3D247F25",
    x"3D24E399",
    x"3D25480C",
    x"3D25AC7E",
    x"3D2610F1",
    x"3D267564",
    x"3D26D9D7",
    x"3D273E49",
    x"3D27A2BC",
    x"3D28072E",
    x"3D286BA0",
    x"3D28D012",
    x"3D293484",
    x"3D2998F6",
    x"3D29FD68",
    x"3D2A61DA",
    x"3D2AC64B",
    x"3D2B2ABD",
    x"3D2B8F2E",
    x"3D2BF39F",
    x"3D2C5811",
    x"3D2CBC82",
    x"3D2D20F3",
    x"3D2D8564",
    x"3D2DE9D4",
    x"3D2E4E45",
    x"3D2EB2B6",
    x"3D2F1726",
    x"3D2F7B96",
    x"3D2FE007",
    x"3D304477",
    x"3D30A8E7",
    x"3D310D57",
    x"3D3171C6",
    x"3D31D636",
    x"3D323AA6",
    x"3D329F15",
    x"3D330385",
    x"3D3367F4",
    x"3D33CC63",
    x"3D3430D2",
    x"3D349541",
    x"3D34F9B0",
    x"3D355E1F",
    x"3D35C28D",
    x"3D3626FC",
    x"3D368B6A",
    x"3D36EFD9",
    x"3D375447",
    x"3D37B8B5",
    x"3D381D23",
    x"3D388191",
    x"3D38E5FE",
    x"3D394A6C",
    x"3D39AEDA",
    x"3D3A1347",
    x"3D3A77B4",
    x"3D3ADC22",
    x"3D3B408F",
    x"3D3BA4FC",
    x"3D3C0968",
    x"3D3C6DD5",
    x"3D3CD242",
    x"3D3D36AE",
    x"3D3D9B1B",
    x"3D3DFF87",
    x"3D3E63F3",
    x"3D3EC85F",
    x"3D3F2CCB",
    x"3D3F9137",
    x"3D3FF5A3",
    x"3D405A0E",
    x"3D40BE7A",
    x"3D4122E5",
    x"3D418750",
    x"3D41EBBB",
    x"3D425026",
    x"3D42B491",
    x"3D4318FC",
    x"3D437D67",
    x"3D43E1D1",
    x"3D44463C",
    x"3D44AAA6",
    x"3D450F10",
    x"3D45737A",
    x"3D45D7E4",
    x"3D463C4E",
    x"3D46A0B8",
    x"3D470521",
    x"3D47698B",
    x"3D47CDF4",
    x"3D48325D",
    x"3D4896C7",
    x"3D48FB30",
    x"3D495F98",
    x"3D49C401",
    x"3D4A286A",
    x"3D4A8CD2",
    x"3D4AF13B",
    x"3D4B55A3",
    x"3D4BBA0B",
    x"3D4C1E73",
    x"3D4C82DB",
    x"3D4CE743",
    x"3D4D4BAA",
    x"3D4DB012",
    x"3D4E1479",
    x"3D4E78E1",
    x"3D4EDD48",
    x"3D4F41AF",
    x"3D4FA616",
    x"3D500A7C",
    x"3D506EE3",
    x"3D50D34A",
    x"3D5137B0",
    x"3D519C16",
    x"3D52007C",
    x"3D5264E2",
    x"3D52C948",
    x"3D532DAE",
    x"3D539214",
    x"3D53F679",
    x"3D545ADF",
    x"3D54BF44",
    x"3D5523A9",
    x"3D55880E",
    x"3D55EC73",
    x"3D5650D8",
    x"3D56B53C",
    x"3D5719A1",
    x"3D577E05",
    x"3D57E269",
    x"3D5846CD",
    x"3D58AB31",
    x"3D590F95",
    x"3D5973F9",
    x"3D59D85C",
    x"3D5A3CC0",
    x"3D5AA123",
    x"3D5B0586",
    x"3D5B69E9",
    x"3D5BCE4C",
    x"3D5C32AF",
    x"3D5C9712",
    x"3D5CFB74",
    x"3D5D5FD7",
    x"3D5DC439",
    x"3D5E289B",
    x"3D5E8CFD",
    x"3D5EF15F",
    x"3D5F55C0",
    x"3D5FBA22",
    x"3D601E83",
    x"3D6082E5",
    x"3D60E746",
    x"3D614BA7",
    x"3D61B008",
    x"3D621469",
    x"3D6278C9",
    x"3D62DD2A",
    x"3D63418A",
    x"3D63A5EA",
    x"3D640A4A",
    x"3D646EAA",
    x"3D64D30A",
    x"3D65376A",
    x"3D659BC9",
    x"3D660029",
    x"3D666488",
    x"3D66C8E7",
    x"3D672D46",
    x"3D6791A5",
    x"3D67F604",
    x"3D685A62",
    x"3D68BEC1",
    x"3D69231F",
    x"3D69877D",
    x"3D69EBDB",
    x"3D6A5039",
    x"3D6AB496",
    x"3D6B18F4",
    x"3D6B7D51",
    x"3D6BE1AF",
    x"3D6C460C",
    x"3D6CAA69",
    x"3D6D0EC6",
    x"3D6D7323",
    x"3D6DD77F",
    x"3D6E3BDC",
    x"3D6EA038",
    x"3D6F0494",
    x"3D6F68F0",
    x"3D6FCD4C",
    x"3D7031A8",
    x"3D709603",
    x"3D70FA5E",
    x"3D715EBA",
    x"3D71C315",
    x"3D722770",
    x"3D728BCB",
    x"3D72F025",
    x"3D735480",
    x"3D73B8DA",
    x"3D741D35",
    x"3D74818F",
    x"3D74E5E9",
    x"3D754A42",
    x"3D75AE9C",
    x"3D7612F6",
    x"3D76774F",
    x"3D76DBA8",
    x"3D774001",
    x"3D77A45A",
    x"3D7808B3",
    x"3D786D0C",
    x"3D78D164",
    x"3D7935BC",
    x"3D799A15",
    x"3D79FE6D",
    x"3D7A62C5",
    x"3D7AC71C",
    x"3D7B2B74",
    x"3D7B8FCB",
    x"3D7BF422",
    x"3D7C587A",
    x"3D7CBCD1",
    x"3D7D2127",
    x"3D7D857E",
    x"3D7DE9D5",
    x"3D7E4E2B",
    x"3D7EB281",
    x"3D7F16D7",
    x"3D7F7B2D",
    x"3D7FDF83",
    x"3D8021EC",
    x"3D805417",
    x"3D808642",
    x"3D80B86C",
    x"3D80EA97",
    x"3D811CC1",
    x"3D814EEB",
    x"3D818116",
    x"3D81B340",
    x"3D81E56A",
    x"3D821794",
    x"3D8249BE",
    x"3D827BE8",
    x"3D82AE11",
    x"3D82E03B",
    x"3D831265",
    x"3D83448E",
    x"3D8376B8",
    x"3D83A8E1",
    x"3D83DB0A",
    x"3D840D34",
    x"3D843F5D",
    x"3D847186",
    x"3D84A3AF",
    x"3D84D5D8",
    x"3D850801",
    x"3D853A29",
    x"3D856C52",
    x"3D859E7B",
    x"3D85D0A3",
    x"3D8602CC",
    x"3D8634F4",
    x"3D86671C",
    x"3D869944",
    x"3D86CB6C",
    x"3D86FD94",
    x"3D872FBC",
    x"3D8761E4",
    x"3D87940C",
    x"3D87C634",
    x"3D87F85B",
    x"3D882A83",
    x"3D885CAA",
    x"3D888ED2",
    x"3D88C0F9",
    x"3D88F320",
    x"3D892547",
    x"3D89576E",
    x"3D898995",
    x"3D89BBBC",
    x"3D89EDE3",
    x"3D8A200A",
    x"3D8A5230",
    x"3D8A8457",
    x"3D8AB67D",
    x"3D8AE8A4",
    x"3D8B1ACA",
    x"3D8B4CF0",
    x"3D8B7F16",
    x"3D8BB13C",
    x"3D8BE362",
    x"3D8C1588",
    x"3D8C47AE",
    x"3D8C79D4",
    x"3D8CABF9",
    x"3D8CDE1F",
    x"3D8D1044",
    x"3D8D426A",
    x"3D8D748F",
    x"3D8DA6B4",
    x"3D8DD8D9",
    x"3D8E0AFE",
    x"3D8E3D23",
    x"3D8E6F48",
    x"3D8EA16D",
    x"3D8ED391",
    x"3D8F05B6",
    x"3D8F37DA",
    x"3D8F69FF",
    x"3D8F9C23",
    x"3D8FCE47",
    x"3D90006C",
    x"3D903290",
    x"3D9064B4",
    x"3D9096D8",
    x"3D90C8FB",
    x"3D90FB1F",
    x"3D912D43",
    x"3D915F66",
    x"3D91918A",
    x"3D91C3AD",
    x"3D91F5D0",
    x"3D9227F4",
    x"3D925A17",
    x"3D928C3A",
    x"3D92BE5D",
    x"3D92F07F",
    x"3D9322A2",
    x"3D9354C5",
    x"3D9386E7",
    x"3D93B90A",
    x"3D93EB2C",
    x"3D941D4F",
    x"3D944F71",
    x"3D948193",
    x"3D94B3B5",
    x"3D94E5D7",
    x"3D9517F9",
    x"3D954A1B",
    x"3D957C3C",
    x"3D95AE5E",
    x"3D95E07F",
    x"3D9612A1",
    x"3D9644C2",
    x"3D9676E3",
    x"3D96A905",
    x"3D96DB26",
    x"3D970D47",
    x"3D973F67",
    x"3D977188",
    x"3D97A3A9",
    x"3D97D5CA",
    x"3D9807EA",
    x"3D983A0A",
    x"3D986C2B",
    x"3D989E4B",
    x"3D98D06B",
    x"3D99028B",
    x"3D9934AB",
    x"3D9966CB",
    x"3D9998EB",
    x"3D99CB0A",
    x"3D99FD2A",
    x"3D9A2F4A",
    x"3D9A6169",
    x"3D9A9388",
    x"3D9AC5A7",
    x"3D9AF7C7",
    x"3D9B29E6",
    x"3D9B5C05",
    x"3D9B8E23",
    x"3D9BC042",
    x"3D9BF261",
    x"3D9C247F",
    x"3D9C569E",
    x"3D9C88BC",
    x"3D9CBADA",
    x"3D9CECF9",
    x"3D9D1F17",
    x"3D9D5135",
    x"3D9D8353",
    x"3D9DB570",
    x"3D9DE78E",
    x"3D9E19AC",
    x"3D9E4BC9",
    x"3D9E7DE7",
    x"3D9EB004",
    x"3D9EE221",
    x"3D9F143E",
    x"3D9F465B",
    x"3D9F7878",
    x"3D9FAA95",
    x"3D9FDCB2",
    x"3DA00ECF",
    x"3DA040EB",
    x"3DA07308",
    x"3DA0A524",
    x"3DA0D740",
    x"3DA1095C",
    x"3DA13B78",
    x"3DA16D94",
    x"3DA19FB0",
    x"3DA1D1CC",
    x"3DA203E8",
    x"3DA23603",
    x"3DA2681F",
    x"3DA29A3A",
    x"3DA2CC55",
    x"3DA2FE71",
    x"3DA3308C",
    x"3DA362A7",
    x"3DA394C2",
    x"3DA3C6DC",
    x"3DA3F8F7",
    x"3DA42B12",
    x"3DA45D2C",
    x"3DA48F47",
    x"3DA4C161",
    x"3DA4F37B",
    x"3DA52595",
    x"3DA557AF",
    x"3DA589C9",
    x"3DA5BBE3",
    x"3DA5EDFD",
    x"3DA62016",
    x"3DA65230",
    x"3DA68449",
    x"3DA6B663",
    x"3DA6E87C",
    x"3DA71A95",
    x"3DA74CAE",
    x"3DA77EC7",
    x"3DA7B0E0",
    x"3DA7E2F8",
    x"3DA81511",
    x"3DA84729",
    x"3DA87942",
    x"3DA8AB5A",
    x"3DA8DD72",
    x"3DA90F8A",
    x"3DA941A2",
    x"3DA973BA",
    x"3DA9A5D2",
    x"3DA9D7EA",
    x"3DAA0A01",
    x"3DAA3C19",
    x"3DAA6E30",
    x"3DAAA048",
    x"3DAAD25F",
    x"3DAB0476",
    x"3DAB368D",
    x"3DAB68A4",
    x"3DAB9ABA",
    x"3DABCCD1",
    x"3DABFEE8",
    x"3DAC30FE",
    x"3DAC6314",
    x"3DAC952B",
    x"3DACC741",
    x"3DACF957",
    x"3DAD2B6D",
    x"3DAD5D83",
    x"3DAD8F98",
    x"3DADC1AE",
    x"3DADF3C3",
    x"3DAE25D9",
    x"3DAE57EE",
    x"3DAE8A03",
    x"3DAEBC18",
    x"3DAEEE2D",
    x"3DAF2042",
    x"3DAF5257",
    x"3DAF846C",
    x"3DAFB680",
    x"3DAFE895",
    x"3DB01AA9",
    x"3DB04CBD",
    x"3DB07ED2",
    x"3DB0B0E6",
    x"3DB0E2FA",
    x"3DB1150D",
    x"3DB14721",
    x"3DB17935",
    x"3DB1AB48",
    x"3DB1DD5C",
    x"3DB20F6F",
    x"3DB24182",
    x"3DB27395",
    x"3DB2A5A8",
    x"3DB2D7BB",
    x"3DB309CE",
    x"3DB33BE0",
    x"3DB36DF3",
    x"3DB3A005",
    x"3DB3D218",
    x"3DB4042A",
    x"3DB4363C",
    x"3DB4684E",
    x"3DB49A60",
    x"3DB4CC72",
    x"3DB4FE83",
    x"3DB53095",
    x"3DB562A6",
    x"3DB594B8",
    x"3DB5C6C9",
    x"3DB5F8DA",
    x"3DB62AEB",
    x"3DB65CFC",
    x"3DB68F0D",
    x"3DB6C11D",
    x"3DB6F32E",
    x"3DB7253E",
    x"3DB7574F",
    x"3DB7895F",
    x"3DB7BB6F",
    x"3DB7ED7F",
    x"3DB81F8F",
    x"3DB8519F",
    x"3DB883AF",
    x"3DB8B5BE",
    x"3DB8E7CE",
    x"3DB919DD",
    x"3DB94BEC",
    x"3DB97DFB",
    x"3DB9B00A",
    x"3DB9E219",
    x"3DBA1428",
    x"3DBA4637",
    x"3DBA7845",
    x"3DBAAA54",
    x"3DBADC62",
    x"3DBB0E70",
    x"3DBB407E",
    x"3DBB728C",
    x"3DBBA49A",
    x"3DBBD6A8",
    x"3DBC08B6",
    x"3DBC3AC3",
    x"3DBC6CD1",
    x"3DBC9EDE",
    x"3DBCD0EB",
    x"3DBD02F8",
    x"3DBD3505",
    x"3DBD6712",
    x"3DBD991F",
    x"3DBDCB2C",
    x"3DBDFD38",
    x"3DBE2F45",
    x"3DBE6151",
    x"3DBE935D",
    x"3DBEC569",
    x"3DBEF775",
    x"3DBF2981",
    x"3DBF5B8D",
    x"3DBF8D98",
    x"3DBFBFA4",
    x"3DBFF1AF",
    x"3DC023BA",
    x"3DC055C6",
    x"3DC087D1",
    x"3DC0B9DC",
    x"3DC0EBE6",
    x"3DC11DF1",
    x"3DC14FFC",
    x"3DC18206",
    x"3DC1B410",
    x"3DC1E61B",
    x"3DC21825",
    x"3DC24A2F",
    x"3DC27C39",
    x"3DC2AE42",
    x"3DC2E04C",
    x"3DC31255",
    x"3DC3445F",
    x"3DC37668",
    x"3DC3A871",
    x"3DC3DA7A",
    x"3DC40C83",
    x"3DC43E8C",
    x"3DC47095",
    x"3DC4A29D",
    x"3DC4D4A6",
    x"3DC506AE",
    x"3DC538B6",
    x"3DC56ABE",
    x"3DC59CC6",
    x"3DC5CECE",
    x"3DC600D6",
    x"3DC632DE",
    x"3DC664E5",
    x"3DC696ED",
    x"3DC6C8F4",
    x"3DC6FAFB",
    x"3DC72D02",
    x"3DC75F09",
    x"3DC79110",
    x"3DC7C316",
    x"3DC7F51D",
    x"3DC82723",
    x"3DC8592A",
    x"3DC88B30",
    x"3DC8BD36",
    x"3DC8EF3C",
    x"3DC92142",
    x"3DC95347",
    x"3DC9854D",
    x"3DC9B752",
    x"3DC9E958",
    x"3DCA1B5D",
    x"3DCA4D62",
    x"3DCA7F67",
    x"3DCAB16C",
    x"3DCAE371",
    x"3DCB1575",
    x"3DCB477A",
    x"3DCB797E",
    x"3DCBAB82",
    x"3DCBDD86",
    x"3DCC0F8A",
    x"3DCC418E",
    x"3DCC7392",
    x"3DCCA596",
    x"3DCCD799",
    x"3DCD099C",
    x"3DCD3BA0",
    x"3DCD6DA3",
    x"3DCD9FA6",
    x"3DCDD1A9",
    x"3DCE03AB",
    x"3DCE35AE",
    x"3DCE67B1",
    x"3DCE99B3",
    x"3DCECBB5",
    x"3DCEFDB7",
    x"3DCF2FB9",
    x"3DCF61BB",
    x"3DCF93BD",
    x"3DCFC5BF",
    x"3DCFF7C0",
    x"3DD029C2",
    x"3DD05BC3",
    x"3DD08DC4",
    x"3DD0BFC5",
    x"3DD0F1C6",
    x"3DD123C7",
    x"3DD155C7",
    x"3DD187C8",
    x"3DD1B9C8",
    x"3DD1EBC8",
    x"3DD21DC8",
    x"3DD24FC8",
    x"3DD281C8",
    x"3DD2B3C8",
    x"3DD2E5C8",
    x"3DD317C7",
    x"3DD349C7",
    x"3DD37BC6",
    x"3DD3ADC5",
    x"3DD3DFC4",
    x"3DD411C3",
    x"3DD443C1",
    x"3DD475C0",
    x"3DD4A7BE",
    x"3DD4D9BD",
    x"3DD50BBB",
    x"3DD53DB9",
    x"3DD56FB7",
    x"3DD5A1B5",
    x"3DD5D3B3",
    x"3DD605B0",
    x"3DD637AE",
    x"3DD669AB",
    x"3DD69BA8",
    x"3DD6CDA5",
    x"3DD6FFA2",
    x"3DD7319F",
    x"3DD7639C",
    x"3DD79598",
    x"3DD7C795",
    x"3DD7F991",
    x"3DD82B8D",
    x"3DD85D89",
    x"3DD88F85",
    x"3DD8C181",
    x"3DD8F37C",
    x"3DD92578",
    x"3DD95773",
    x"3DD9896E",
    x"3DD9BB69",
    x"3DD9ED64",
    x"3DDA1F5F",
    x"3DDA515A",
    x"3DDA8354",
    x"3DDAB54F",
    x"3DDAE749",
    x"3DDB1943",
    x"3DDB4B3D",
    x"3DDB7D37",
    x"3DDBAF31",
    x"3DDBE12B",
    x"3DDC1324",
    x"3DDC451E",
    x"3DDC7717",
    x"3DDCA910",
    x"3DDCDB09",
    x"3DDD0D02",
    x"3DDD3EFB",
    x"3DDD70F3",
    x"3DDDA2EC",
    x"3DDDD4E4",
    x"3DDE06DC",
    x"3DDE38D4",
    x"3DDE6ACC",
    x"3DDE9CC4",
    x"3DDECEBC",
    x"3DDF00B3",
    x"3DDF32AB",
    x"3DDF64A2",
    x"3DDF9699",
    x"3DDFC890",
    x"3DDFFA87",
    x"3DE02C7D",
    x"3DE05E74",
    x"3DE0906A",
    x"3DE0C261",
    x"3DE0F457",
    x"3DE1264D",
    x"3DE15843",
    x"3DE18A39",
    x"3DE1BC2E",
    x"3DE1EE24",
    x"3DE22019",
    x"3DE2520E",
    x"3DE28403",
    x"3DE2B5F8",
    x"3DE2E7ED",
    x"3DE319E2",
    x"3DE34BD6",
    x"3DE37DCB",
    x"3DE3AFBF",
    x"3DE3E1B3",
    x"3DE413A7",
    x"3DE4459B",
    x"3DE4778F",
    x"3DE4A982",
    x"3DE4DB76",
    x"3DE50D69",
    x"3DE53F5C",
    x"3DE5714F",
    x"3DE5A342",
    x"3DE5D535",
    x"3DE60727",
    x"3DE6391A",
    x"3DE66B0C",
    x"3DE69CFE",
    x"3DE6CEF0",
    x"3DE700E2",
    x"3DE732D4",
    x"3DE764C6",
    x"3DE796B7",
    x"3DE7C8A9",
    x"3DE7FA9A",
    x"3DE82C8B",
    x"3DE85E7C",
    x"3DE8906D",
    x"3DE8C25D",
    x"3DE8F44E",
    x"3DE9263E",
    x"3DE9582E",
    x"3DE98A1F",
    x"3DE9BC0E",
    x"3DE9EDFE",
    x"3DEA1FEE",
    x"3DEA51DE",
    x"3DEA83CD",
    x"3DEAB5BC",
    x"3DEAE7AB",
    x"3DEB199A",
    x"3DEB4B89",
    x"3DEB7D78",
    x"3DEBAF66",
    x"3DEBE155",
    x"3DEC1343",
    x"3DEC4531",
    x"3DEC771F",
    x"3DECA90D",
    x"3DECDAFB",
    x"3DED0CE8",
    x"3DED3ED5",
    x"3DED70C3",
    x"3DEDA2B0",
    x"3DEDD49D",
    x"3DEE068A",
    x"3DEE3876",
    x"3DEE6A63",
    x"3DEE9C4F",
    x"3DEECE3C",
    x"3DEF0028",
    x"3DEF3214",
    x"3DEF63FF",
    x"3DEF95EB",
    x"3DEFC7D7",
    x"3DEFF9C2",
    x"3DF02BAD",
    x"3DF05D98",
    x"3DF08F83",
    x"3DF0C16E",
    x"3DF0F359",
    x"3DF12543",
    x"3DF1572E",
    x"3DF18918",
    x"3DF1BB02",
    x"3DF1ECEC",
    x"3DF21ED6",
    x"3DF250BF",
    x"3DF282A9",
    x"3DF2B492",
    x"3DF2E67C",
    x"3DF31865",
    x"3DF34A4E",
    x"3DF37C36",
    x"3DF3AE1F",
    x"3DF3E007",
    x"3DF411F0",
    x"3DF443D8",
    x"3DF475C0",
    x"3DF4A7A8",
    x"3DF4D990",
    x"3DF50B77",
    x"3DF53D5F",
    x"3DF56F46",
    x"3DF5A12D",
    x"3DF5D314",
    x"3DF604FB",
    x"3DF636E2",
    x"3DF668C8",
    x"3DF69AAF",
    x"3DF6CC95",
    x"3DF6FE7B",
    x"3DF73061",
    x"3DF76247",
    x"3DF7942C",
    x"3DF7C612",
    x"3DF7F7F7",
    x"3DF829DD",
    x"3DF85BC2",
    x"3DF88DA7",
    x"3DF8BF8B",
    x"3DF8F170",
    x"3DF92354",
    x"3DF95539",
    x"3DF9871D",
    x"3DF9B901",
    x"3DF9EAE5",
    x"3DFA1CC8",
    x"3DFA4EAC",
    x"3DFA808F",
    x"3DFAB273",
    x"3DFAE456",
    x"3DFB1639",
    x"3DFB481C",
    x"3DFB79FE",
    x"3DFBABE1",
    x"3DFBDDC3",
    x"3DFC0FA5",
    x"3DFC4187",
    x"3DFC7369",
    x"3DFCA54B",
    x"3DFCD72D",
    x"3DFD090E",
    x"3DFD3AEF",
    x"3DFD6CD1",
    x"3DFD9EB2",
    x"3DFDD092",
    x"3DFE0273",
    x"3DFE3454",
    x"3DFE6634",
    x"3DFE9814",
    x"3DFEC9F4",
    x"3DFEFBD4",
    x"3DFF2DB4",
    x"3DFF5F94",
    x"3DFF9173",
    x"3DFFC352",
    x"3DFFF531",
    x"3E001388",
    x"3E002C78",
    x"3E004567",
    x"3E005E56",
    x"3E007745",
    x"3E009035",
    x"3E00A924",
    x"3E00C213",
    x"3E00DB01",
    x"3E00F3F0",
    x"3E010CDF",
    x"3E0125CE",
    x"3E013EBC",
    x"3E0157AB",
    x"3E017099",
    x"3E018987",
    x"3E01A276",
    x"3E01BB64",
    x"3E01D452",
    x"3E01ED40",
    x"3E02062E",
    x"3E021F1C",
    x"3E02380A",
    x"3E0250F7",
    x"3E0269E5",
    x"3E0282D2",
    x"3E029BC0",
    x"3E02B4AD",
    x"3E02CD9B",
    x"3E02E688",
    x"3E02FF75",
    x"3E031862",
    x"3E03314F",
    x"3E034A3C",
    x"3E036329",
    x"3E037C16",
    x"3E039502",
    x"3E03ADEF",
    x"3E03C6DB",
    x"3E03DFC8",
    x"3E03F8B4",
    x"3E0411A0",
    x"3E042A8D",
    x"3E044379",
    x"3E045C65",
    x"3E047551",
    x"3E048E3D",
    x"3E04A729",
    x"3E04C014",
    x"3E04D900",
    x"3E04F1EB",
    x"3E050AD7",
    x"3E0523C2",
    x"3E053CAE",
    x"3E055599",
    x"3E056E84",
    x"3E05876F",
    x"3E05A05A",
    x"3E05B945",
    x"3E05D230",
    x"3E05EB1B",
    x"3E060405",
    x"3E061CF0",
    x"3E0635DB",
    x"3E064EC5",
    x"3E0667AF",
    x"3E06809A",
    x"3E069984",
    x"3E06B26E",
    x"3E06CB58",
    x"3E06E442",
    x"3E06FD2C",
    x"3E071616",
    x"3E072EFF",
    x"3E0747E9",
    x"3E0760D2",
    x"3E0779BC",
    x"3E0792A5",
    x"3E07AB8F",
    x"3E07C478",
    x"3E07DD61",
    x"3E07F64A",
    x"3E080F33",
    x"3E08281C",
    x"3E084105",
    x"3E0859ED",
    x"3E0872D6",
    x"3E088BBF",
    x"3E08A4A7",
    x"3E08BD90",
    x"3E08D678",
    x"3E08EF60",
    x"3E090848",
    x"3E092130",
    x"3E093A18",
    x"3E095300",
    x"3E096BE8",
    x"3E0984D0",
    x"3E099DB7",
    x"3E09B69F",
    x"3E09CF86",
    x"3E09E86E",
    x"3E0A0155",
    x"3E0A1A3C",
    x"3E0A3324",
    x"3E0A4C0B",
    x"3E0A64F2",
    x"3E0A7DD9",
    x"3E0A96BF",
    x"3E0AAFA6",
    x"3E0AC88D",
    x"3E0AE173",
    x"3E0AFA5A",
    x"3E0B1340",
    x"3E0B2C27",
    x"3E0B450D",
    x"3E0B5DF3",
    x"3E0B76D9",
    x"3E0B8FBF",
    x"3E0BA8A5",
    x"3E0BC18B",
    x"3E0BDA71",
    x"3E0BF356",
    x"3E0C0C3C",
    x"3E0C2521",
    x"3E0C3E07",
    x"3E0C56EC",
    x"3E0C6FD1",
    x"3E0C88B6",
    x"3E0CA19B",
    x"3E0CBA80",
    x"3E0CD365",
    x"3E0CEC4A",
    x"3E0D052F",
    x"3E0D1E13",
    x"3E0D36F8",
    x"3E0D4FDC",
    x"3E0D68C1",
    x"3E0D81A5",
    x"3E0D9A89",
    x"3E0DB36D",
    x"3E0DCC51",
    x"3E0DE535",
    x"3E0DFE19",
    x"3E0E16FD",
    x"3E0E2FE1",
    x"3E0E48C4",
    x"3E0E61A8",
    x"3E0E7A8B",
    x"3E0E936F",
    x"3E0EAC52",
    x"3E0EC535",
    x"3E0EDE18",
    x"3E0EF6FB",
    x"3E0F0FDE",
    x"3E0F28C1",
    x"3E0F41A4",
    x"3E0F5A86",
    x"3E0F7369",
    x"3E0F8C4B",
    x"3E0FA52E",
    x"3E0FBE10",
    x"3E0FD6F2",
    x"3E0FEFD5",
    x"3E1008B7",
    x"3E102199",
    x"3E103A7B",
    x"3E10535C",
    x"3E106C3E",
    x"3E108520",
    x"3E109E01",
    x"3E10B6E3",
    x"3E10CFC4",
    x"3E10E8A5",
    x"3E110186",
    x"3E111A68",
    x"3E113349",
    x"3E114C2A",
    x"3E11650A",
    x"3E117DEB",
    x"3E1196CC",
    x"3E11AFAC",
    x"3E11C88D",
    x"3E11E16D",
    x"3E11FA4E",
    x"3E12132E",
    x"3E122C0E",
    x"3E1244EE",
    x"3E125DCE",
    x"3E1276AE",
    x"3E128F8E",
    x"3E12A86D",
    x"3E12C14D",
    x"3E12DA2C",
    x"3E12F30C",
    x"3E130BEB",
    x"3E1324CA",
    x"3E133DAA",
    x"3E135689",
    x"3E136F68",
    x"3E138847",
    x"3E13A125",
    x"3E13BA04",
    x"3E13D2E3",
    x"3E13EBC1",
    x"3E1404A0",
    x"3E141D7E",
    x"3E14365C",
    x"3E144F3B",
    x"3E146819",
    x"3E1480F7",
    x"3E1499D5",
    x"3E14B2B2",
    x"3E14CB90",
    x"3E14E46E",
    x"3E14FD4B",
    x"3E151629",
    x"3E152F06",
    x"3E1547E4",
    x"3E1560C1",
    x"3E15799E",
    x"3E15927B",
    x"3E15AB58",
    x"3E15C435",
    x"3E15DD11",
    x"3E15F5EE",
    x"3E160ECB",
    x"3E1627A7",
    x"3E164083",
    x"3E165960",
    x"3E16723C",
    x"3E168B18",
    x"3E16A3F4",
    x"3E16BCD0",
    x"3E16D5AC",
    x"3E16EE88",
    x"3E170763",
    x"3E17203F",
    x"3E17391A",
    x"3E1751F6",
    x"3E176AD1",
    x"3E1783AC",
    x"3E179C87",
    x"3E17B562",
    x"3E17CE3D",
    x"3E17E718",
    x"3E17FFF3",
    x"3E1818CE",
    x"3E1831A8",
    x"3E184A83",
    x"3E18635D",
    x"3E187C37",
    x"3E189511",
    x"3E18ADEC",
    x"3E18C6C6",
    x"3E18DFA0",
    x"3E18F879",
    x"3E191153",
    x"3E192A2D",
    x"3E194306",
    x"3E195BE0",
    x"3E1974B9",
    x"3E198D92",
    x"3E19A66C",
    x"3E19BF45",
    x"3E19D81E",
    x"3E19F0F7",
    x"3E1A09CF",
    x"3E1A22A8",
    x"3E1A3B81",
    x"3E1A5459",
    x"3E1A6D32",
    x"3E1A860A",
    x"3E1A9EE2",
    x"3E1AB7BB",
    x"3E1AD093",
    x"3E1AE96B",
    x"3E1B0242",
    x"3E1B1B1A",
    x"3E1B33F2",
    x"3E1B4CCA",
    x"3E1B65A1",
    x"3E1B7E79",
    x"3E1B9750",
    x"3E1BB027",
    x"3E1BC8FE",
    x"3E1BE1D5",
    x"3E1BFAAC",
    x"3E1C1383",
    x"3E1C2C5A",
    x"3E1C4530",
    x"3E1C5E07",
    x"3E1C76DE",
    x"3E1C8FB4",
    x"3E1CA88A",
    x"3E1CC160",
    x"3E1CDA36",
    x"3E1CF30D",
    x"3E1D0BE2",
    x"3E1D24B8",
    x"3E1D3D8E",
    x"3E1D5664",
    x"3E1D6F39",
    x"3E1D880F",
    x"3E1DA0E4",
    x"3E1DB9B9",
    x"3E1DD28E",
    x"3E1DEB63",
    x"3E1E0438",
    x"3E1E1D0D",
    x"3E1E35E2",
    x"3E1E4EB7",
    x"3E1E678B",
    x"3E1E8060",
    x"3E1E9934",
    x"3E1EB208",
    x"3E1ECADD",
    x"3E1EE3B1",
    x"3E1EFC85",
    x"3E1F1559",
    x"3E1F2E2C",
    x"3E1F4700",
    x"3E1F5FD4",
    x"3E1F78A7",
    x"3E1F917B",
    x"3E1FAA4E",
    x"3E1FC321",
    x"3E1FDBF4",
    x"3E1FF4C8",
    x"3E200D9A",
    x"3E20266D",
    x"3E203F40",
    x"3E205813",
    x"3E2070E5",
    x"3E2089B8",
    x"3E20A28A",
    x"3E20BB5C",
    x"3E20D42F",
    x"3E20ED01",
    x"3E2105D3",
    x"3E211EA5",
    x"3E213776",
    x"3E215048",
    x"3E21691A",
    x"3E2181EB",
    x"3E219ABD",
    x"3E21B38E",
    x"3E21CC5F",
    x"3E21E530",
    x"3E21FE01",
    x"3E2216D2",
    x"3E222FA3",
    x"3E224874",
    x"3E226144",
    x"3E227A15",
    x"3E2292E5",
    x"3E22ABB6",
    x"3E22C486",
    x"3E22DD56",
    x"3E22F626",
    x"3E230EF6",
    x"3E2327C6",
    x"3E234095",
    x"3E235965",
    x"3E237235",
    x"3E238B04",
    x"3E23A3D3",
    x"3E23BCA3",
    x"3E23D572",
    x"3E23EE41",
    x"3E240710",
    x"3E241FDF",
    x"3E2438AD",
    x"3E24517C",
    x"3E246A4B",
    x"3E248319",
    x"3E249BE7",
    x"3E24B4B6",
    x"3E24CD84",
    x"3E24E652",
    x"3E24FF20",
    x"3E2517EE",
    x"3E2530BC",
    x"3E254989",
    x"3E256257",
    x"3E257B24",
    x"3E2593F2",
    x"3E25ACBF",
    x"3E25C58C",
    x"3E25DE59",
    x"3E25F726",
    x"3E260FF3",
    x"3E2628C0",
    x"3E26418C",
    x"3E265A59",
    x"3E267325",
    x"3E268BF2",
    x"3E26A4BE",
    x"3E26BD8A",
    x"3E26D656",
    x"3E26EF22",
    x"3E2707EE",
    x"3E2720BA",
    x"3E273985",
    x"3E275251",
    x"3E276B1C",
    x"3E2783E8",
    x"3E279CB3",
    x"3E27B57E",
    x"3E27CE49",
    x"3E27E714",
    x"3E27FFDF",
    x"3E2818AA",
    x"3E283174",
    x"3E284A3F",
    x"3E286309",
    x"3E287BD4",
    x"3E28949E",
    x"3E28AD68",
    x"3E28C632",
    x"3E28DEFC",
    x"3E28F7C6",
    x"3E291090",
    x"3E292959",
    x"3E294223",
    x"3E295AEC",
    x"3E2973B6",
    x"3E298C7F",
    x"3E29A548",
    x"3E29BE11",
    x"3E29D6DA",
    x"3E29EFA3",
    x"3E2A086B",
    x"3E2A2134",
    x"3E2A39FD",
    x"3E2A52C5",
    x"3E2A6B8D",
    x"3E2A8456",
    x"3E2A9D1E",
    x"3E2AB5E6",
    x"3E2ACEAE",
    x"3E2AE775",
    x"3E2B003D",
    x"3E2B1905",
    x"3E2B31CC",
    x"3E2B4A93",
    x"3E2B635B",
    x"3E2B7C22",
    x"3E2B94E9",
    x"3E2BADB0",
    x"3E2BC677",
    x"3E2BDF3E",
    x"3E2BF804",
    x"3E2C10CB",
    x"3E2C2991",
    x"3E2C4258",
    x"3E2C5B1E",
    x"3E2C73E4",
    x"3E2C8CAA",
    x"3E2CA570",
    x"3E2CBE36",
    x"3E2CD6FB",
    x"3E2CEFC1",
    x"3E2D0887",
    x"3E2D214C",
    x"3E2D3A11",
    x"3E2D52D6",
    x"3E2D6B9C",
    x"3E2D8461",
    x"3E2D9D25",
    x"3E2DB5EA",
    x"3E2DCEAF",
    x"3E2DE773",
    x"3E2E0038",
    x"3E2E18FC",
    x"3E2E31C1",
    x"3E2E4A85",
    x"3E2E6349",
    x"3E2E7C0D",
    x"3E2E94D1",
    x"3E2EAD94",
    x"3E2EC658",
    x"3E2EDF1B",
    x"3E2EF7DF",
    x"3E2F10A2",
    x"3E2F2965",
    x"3E2F4228",
    x"3E2F5AEB",
    x"3E2F73AE",
    x"3E2F8C71",
    x"3E2FA534",
    x"3E2FBDF6",
    x"3E2FD6B9",
    x"3E2FEF7B",
    x"3E30083D",
    x"3E302100",
    x"3E3039C2",
    x"3E305284",
    x"3E306B45",
    x"3E308407",
    x"3E309CC9",
    x"3E30B58A",
    x"3E30CE4C",
    x"3E30E70D",
    x"3E30FFCE",
    x"3E31188F",
    x"3E313150",
    x"3E314A11",
    x"3E3162D2",
    x"3E317B92",
    x"3E319453",
    x"3E31AD13",
    x"3E31C5D4",
    x"3E31DE94",
    x"3E31F754",
    x"3E321014",
    x"3E3228D4",
    x"3E324194",
    x"3E325A54",
    x"3E327313",
    x"3E328BD3",
    x"3E32A492",
    x"3E32BD51",
    x"3E32D610",
    x"3E32EECF",
    x"3E33078E",
    x"3E33204D",
    x"3E33390C",
    x"3E3351CB",
    x"3E336A89",
    x"3E338348",
    x"3E339C06",
    x"3E33B4C4",
    x"3E33CD82",
    x"3E33E640",
    x"3E33FEFE",
    x"3E3417BC",
    x"3E343079",
    x"3E344937",
    x"3E3461F4",
    x"3E347AB2",
    x"3E34936F",
    x"3E34AC2C",
    x"3E34C4E9",
    x"3E34DDA6",
    x"3E34F662",
    x"3E350F1F",
    x"3E3527DC",
    x"3E354098",
    x"3E355954",
    x"3E357211",
    x"3E358ACD",
    x"3E35A389",
    x"3E35BC45",
    x"3E35D501",
    x"3E35EDBC",
    x"3E360678",
    x"3E361F33",
    x"3E3637EF",
    x"3E3650AA",
    x"3E366965",
    x"3E368220",
    x"3E369ADB",
    x"3E36B396",
    x"3E36CC50",
    x"3E36E50B",
    x"3E36FDC5",
    x"3E371680",
    x"3E372F3A",
    x"3E3747F4",
    x"3E3760AE",
    x"3E377968",
    x"3E379222",
    x"3E37AADC",
    x"3E37C395",
    x"3E37DC4F",
    x"3E37F508",
    x"3E380DC1",
    x"3E38267A",
    x"3E383F33",
    x"3E3857EC",
    x"3E3870A5",
    x"3E38895E",
    x"3E38A217",
    x"3E38BACF",
    x"3E38D387",
    x"3E38EC40",
    x"3E3904F8",
    x"3E391DB0",
    x"3E393668",
    x"3E394F20",
    x"3E3967D7",
    x"3E39808F",
    x"3E399946",
    x"3E39B1FE",
    x"3E39CAB5",
    x"3E39E36C",
    x"3E39FC23",
    x"3E3A14DA",
    x"3E3A2D91",
    x"3E3A4647",
    x"3E3A5EFE",
    x"3E3A77B4",
    x"3E3A906B",
    x"3E3AA921",
    x"3E3AC1D7",
    x"3E3ADA8D",
    x"3E3AF343",
    x"3E3B0BF9",
    x"3E3B24AF",
    x"3E3B3D64",
    x"3E3B561A",
    x"3E3B6ECF",
    x"3E3B8784",
    x"3E3BA039",
    x"3E3BB8EE",
    x"3E3BD1A3",
    x"3E3BEA58",
    x"3E3C030D",
    x"3E3C1BC1",
    x"3E3C3476",
    x"3E3C4D2A",
    x"3E3C65DE",
    x"3E3C7E92",
    x"3E3C9746",
    x"3E3CAFFA",
    x"3E3CC8AE",
    x"3E3CE161",
    x"3E3CFA15",
    x"3E3D12C8",
    x"3E3D2B7C",
    x"3E3D442F",
    x"3E3D5CE2",
    x"3E3D7595",
    x"3E3D8E48",
    x"3E3DA6FA",
    x"3E3DBFAD",
    x"3E3DD860",
    x"3E3DF112",
    x"3E3E09C4",
    x"3E3E2276",
    x"3E3E3B28",
    x"3E3E53DA",
    x"3E3E6C8C",
    x"3E3E853E",
    x"3E3E9DEF",
    x"3E3EB6A1",
    x"3E3ECF52",
    x"3E3EE804",
    x"3E3F00B5",
    x"3E3F1966",
    x"3E3F3217",
    x"3E3F4AC7",
    x"3E3F6378",
    x"3E3F7C29",
    x"3E3F94D9",
    x"3E3FAD89",
    x"3E3FC639",
    x"3E3FDEEA",
    x"3E3FF79A",
    x"3E401049",
    x"3E4028F9",
    x"3E4041A9",
    x"3E405A58",
    x"3E407308",
    x"3E408BB7",
    x"3E40A466",
    x"3E40BD15",
    x"3E40D5C4",
    x"3E40EE73",
    x"3E410722",
    x"3E411FD0",
    x"3E41387F",
    x"3E41512D",
    x"3E4169DB",
    x"3E418289",
    x"3E419B37",
    x"3E41B3E5",
    x"3E41CC93",
    x"3E41E541",
    x"3E41FDEE",
    x"3E42169B",
    x"3E422F49",
    x"3E4247F6",
    x"3E4260A3",
    x"3E427950",
    x"3E4291FD",
    x"3E42AAAA",
    x"3E42C356",
    x"3E42DC03",
    x"3E42F4AF",
    x"3E430D5B",
    x"3E432607",
    x"3E433EB3",
    x"3E43575F",
    x"3E43700B",
    x"3E4388B7",
    x"3E43A162",
    x"3E43BA0E",
    x"3E43D2B9",
    x"3E43EB64",
    x"3E44040F",
    x"3E441CBA",
    x"3E443565",
    x"3E444E10",
    x"3E4466BA",
    x"3E447F65",
    x"3E44980F",
    x"3E44B0B9",
    x"3E44C963",
    x"3E44E20D",
    x"3E44FAB7",
    x"3E451361",
    x"3E452C0B",
    x"3E4544B4",
    x"3E455D5E",
    x"3E457607",
    x"3E458EB0",
    x"3E45A759",
    x"3E45C002",
    x"3E45D8AB",
    x"3E45F153",
    x"3E4609FC",
    x"3E4622A5",
    x"3E463B4D",
    x"3E4653F5",
    x"3E466C9D",
    x"3E468545",
    x"3E469DED",
    x"3E46B695",
    x"3E46CF3C",
    x"3E46E7E4",
    x"3E47008B",
    x"3E471932",
    x"3E4731DA",
    x"3E474A81",
    x"3E476328",
    x"3E477BCE",
    x"3E479475",
    x"3E47AD1B",
    x"3E47C5C2",
    x"3E47DE68",
    x"3E47F70E",
    x"3E480FB4",
    x"3E48285A",
    x"3E484100",
    x"3E4859A6",
    x"3E48724B",
    x"3E488AF1",
    x"3E48A396",
    x"3E48BC3B",
    x"3E48D4E0",
    x"3E48ED85",
    x"3E49062A",
    x"3E491ECF",
    x"3E493774",
    x"3E495018",
    x"3E4968BC",
    x"3E498161",
    x"3E499A05",
    x"3E49B2A9",
    x"3E49CB4D",
    x"3E49E3F0",
    x"3E49FC94",
    x"3E4A1538",
    x"3E4A2DDB",
    x"3E4A467E",
    x"3E4A5F21",
    x"3E4A77C4",
    x"3E4A9067",
    x"3E4AA90A",
    x"3E4AC1AD",
    x"3E4ADA4F",
    x"3E4AF2F2",
    x"3E4B0B94",
    x"3E4B2436",
    x"3E4B3CD8",
    x"3E4B557A",
    x"3E4B6E1C",
    x"3E4B86BE",
    x"3E4B9F5F",
    x"3E4BB801",
    x"3E4BD0A2",
    x"3E4BE943",
    x"3E4C01E4",
    x"3E4C1A85",
    x"3E4C3326",
    x"3E4C4BC7",
    x"3E4C6467",
    x"3E4C7D08",
    x"3E4C95A8",
    x"3E4CAE48",
    x"3E4CC6E8",
    x"3E4CDF88",
    x"3E4CF828",
    x"3E4D10C8",
    x"3E4D2967",
    x"3E4D4207",
    x"3E4D5AA6",
    x"3E4D7345",
    x"3E4D8BE4",
    x"3E4DA483",
    x"3E4DBD22",
    x"3E4DD5C1",
    x"3E4DEE60",
    x"3E4E06FE",
    x"3E4E1F9C",
    x"3E4E383B",
    x"3E4E50D9",
    x"3E4E6977",
    x"3E4E8215",
    x"3E4E9AB2",
    x"3E4EB350",
    x"3E4ECBED",
    x"3E4EE48B",
    x"3E4EFD28",
    x"3E4F15C5",
    x"3E4F2E62",
    x"3E4F46FF",
    x"3E4F5F9C",
    x"3E4F7838",
    x"3E4F90D5",
    x"3E4FA971",
    x"3E4FC20D",
    x"3E4FDAA9",
    x"3E4FF345",
    x"3E500BE1",
    x"3E50247D",
    x"3E503D19",
    x"3E5055B4",
    x"3E506E4F",
    x"3E5086EB",
    x"3E509F86",
    x"3E50B821",
    x"3E50D0BC",
    x"3E50E956",
    x"3E5101F1",
    x"3E511A8B",
    x"3E513326",
    x"3E514BC0",
    x"3E51645A",
    x"3E517CF4",
    x"3E51958E",
    x"3E51AE28",
    x"3E51C6C1",
    x"3E51DF5B",
    x"3E51F7F4",
    x"3E52108D",
    x"3E522926",
    x"3E5241BF",
    x"3E525A58",
    x"3E5272F1",
    x"3E528B89",
    x"3E52A422",
    x"3E52BCBA",
    x"3E52D552",
    x"3E52EDEA",
    x"3E530682",
    x"3E531F1A",
    x"3E5337B2",
    x"3E535049",
    x"3E5368E1",
    x"3E538178",
    x"3E539A0F",
    x"3E53B2A6",
    x"3E53CB3D",
    x"3E53E3D4",
    x"3E53FC6B",
    x"3E541501",
    x"3E542D98",
    x"3E54462E",
    x"3E545EC4",
    x"3E54775A",
    x"3E548FF0",
    x"3E54A886",
    x"3E54C11B",
    x"3E54D9B1",
    x"3E54F246",
    x"3E550ADC",
    x"3E552371",
    x"3E553C06",
    x"3E55549B",
    x"3E556D2F",
    x"3E5585C4",
    x"3E559E58",
    x"3E55B6ED",
    x"3E55CF81",
    x"3E55E815",
    x"3E5600A9",
    x"3E56193D",
    x"3E5631D1",
    x"3E564A64",
    x"3E5662F8",
    x"3E567B8B",
    x"3E56941E",
    x"3E56ACB1",
    x"3E56C544",
    x"3E56DDD7",
    x"3E56F66A",
    x"3E570EFC",
    x"3E57278F",
    x"3E574021",
    x"3E5758B3",
    x"3E577145",
    x"3E5789D7",
    x"3E57A269",
    x"3E57BAFB",
    x"3E57D38C",
    x"3E57EC1D",
    x"3E5804AF",
    x"3E581D40",
    x"3E5835D1",
    x"3E584E62",
    x"3E5866F2",
    x"3E587F83",
    x"3E589813",
    x"3E58B0A4",
    x"3E58C934",
    x"3E58E1C4",
    x"3E58FA54",
    x"3E5912E4",
    x"3E592B74",
    x"3E594403",
    x"3E595C93",
    x"3E597522",
    x"3E598DB1",
    x"3E59A640",
    x"3E59BECF",
    x"3E59D75E",
    x"3E59EFEC",
    x"3E5A087B",
    x"3E5A2109",
    x"3E5A3997",
    x"3E5A5226",
    x"3E5A6AB4",
    x"3E5A8341",
    x"3E5A9BCF",
    x"3E5AB45D",
    x"3E5ACCEA",
    x"3E5AE578",
    x"3E5AFE05",
    x"3E5B1692",
    x"3E5B2F1F",
    x"3E5B47AC",
    x"3E5B6038",
    x"3E5B78C5",
    x"3E5B9151",
    x"3E5BA9DD",
    x"3E5BC26A",
    x"3E5BDAF6",
    x"3E5BF381",
    x"3E5C0C0D",
    x"3E5C2499",
    x"3E5C3D24",
    x"3E5C55B0",
    x"3E5C6E3B",
    x"3E5C86C6",
    x"3E5C9F51",
    x"3E5CB7DC",
    x"3E5CD066",
    x"3E5CE8F1",
    x"3E5D017B",
    x"3E5D1A05",
    x"3E5D3290",
    x"3E5D4B1A",
    x"3E5D63A4",
    x"3E5D7C2D",
    x"3E5D94B7",
    x"3E5DAD40",
    x"3E5DC5CA",
    x"3E5DDE53",
    x"3E5DF6DC",
    x"3E5E0F65",
    x"3E5E27EE",
    x"3E5E4076",
    x"3E5E58FF",
    x"3E5E7187",
    x"3E5E8A10",
    x"3E5EA298",
    x"3E5EBB20",
    x"3E5ED3A8",
    x"3E5EEC2F",
    x"3E5F04B7",
    x"3E5F1D3E",
    x"3E5F35C6",
    x"3E5F4E4D",
    x"3E5F66D4",
    x"3E5F7F5B",
    x"3E5F97E2",
    x"3E5FB068",
    x"3E5FC8EF",
    x"3E5FE175",
    x"3E5FF9FC",
    x"3E601282",
    x"3E602B08",
    x"3E60438E",
    x"3E605C13",
    x"3E607499",
    x"3E608D1E",
    x"3E60A5A4",
    x"3E60BE29",
    x"3E60D6AE",
    x"3E60EF33",
    x"3E6107B8",
    x"3E61203C",
    x"3E6138C1",
    x"3E615145",
    x"3E6169C9",
    x"3E61824D",
    x"3E619AD1",
    x"3E61B355",
    x"3E61CBD9",
    x"3E61E45C",
    x"3E61FCE0",
    x"3E621563",
    x"3E622DE6",
    x"3E624669",
    x"3E625EEC",
    x"3E62776F",
    x"3E628FF1",
    x"3E62A874",
    x"3E62C0F6",
    x"3E62D978",
    x"3E62F1FA",
    x"3E630A7C",
    x"3E6322FE",
    x"3E633B80",
    x"3E635401",
    x"3E636C83",
    x"3E638504",
    x"3E639D85",
    x"3E63B606",
    x"3E63CE87",
    x"3E63E707",
    x"3E63FF88",
    x"3E641808",
    x"3E643089",
    x"3E644909",
    x"3E646189",
    x"3E647A09",
    x"3E649288",
    x"3E64AB08",
    x"3E64C387",
    x"3E64DC07",
    x"3E64F486",
    x"3E650D05",
    x"3E652584",
    x"3E653E02",
    x"3E655681",
    x"3E656F00",
    x"3E65877E",
    x"3E659FFC",
    x"3E65B87A",
    x"3E65D0F8",
    x"3E65E976",
    x"3E6601F3",
    x"3E661A71",
    x"3E6632EE",
    x"3E664B6C",
    x"3E6663E9",
    x"3E667C66",
    x"3E6694E2",
    x"3E66AD5F",
    x"3E66C5DC",
    x"3E66DE58",
    x"3E66F6D4",
    x"3E670F50",
    x"3E6727CC",
    x"3E674048",
    x"3E6758C4",
    x"3E67713F",
    x"3E6789BB",
    x"3E67A236",
    x"3E67BAB1",
    x"3E67D32C",
    x"3E67EBA7",
    x"3E680422",
    x"3E681C9C",
    x"3E683517",
    x"3E684D91",
    x"3E68660B",
    x"3E687E85",
    x"3E6896FF",
    x"3E68AF79",
    x"3E68C7F3",
    x"3E68E06C",
    x"3E68F8E5",
    x"3E69115F",
    x"3E6929D8",
    x"3E694251",
    x"3E695AC9",
    x"3E697342",
    x"3E698BBA",
    x"3E69A433",
    x"3E69BCAB",
    x"3E69D523",
    x"3E69ED9B",
    x"3E6A0613",
    x"3E6A1E8A",
    x"3E6A3702",
    x"3E6A4F79",
    x"3E6A67F0",
    x"3E6A8067",
    x"3E6A98DE",
    x"3E6AB155",
    x"3E6AC9CC",
    x"3E6AE242",
    x"3E6AFAB9",
    x"3E6B132F",
    x"3E6B2BA5",
    x"3E6B441B",
    x"3E6B5C91",
    x"3E6B7506",
    x"3E6B8D7C",
    x"3E6BA5F1",
    x"3E6BBE66",
    x"3E6BD6DC",
    x"3E6BEF51",
    x"3E6C07C5",
    x"3E6C203A",
    x"3E6C38AF",
    x"3E6C5123",
    x"3E6C6997",
    x"3E6C820B",
    x"3E6C9A7F",
    x"3E6CB2F3",
    x"3E6CCB67",
    x"3E6CE3DA",
    x"3E6CFC4E",
    x"3E6D14C1",
    x"3E6D2D34",
    x"3E6D45A7",
    x"3E6D5E1A",
    x"3E6D768C",
    x"3E6D8EFF",
    x"3E6DA771",
    x"3E6DBFE3",
    x"3E6DD856",
    x"3E6DF0C7",
    x"3E6E0939",
    x"3E6E21AB",
    x"3E6E3A1C",
    x"3E6E528E",
    x"3E6E6AFF",
    x"3E6E8370",
    x"3E6E9BE1",
    x"3E6EB452",
    x"3E6ECCC3",
    x"3E6EE533",
    x"3E6EFDA3",
    x"3E6F1614",
    x"3E6F2E84",
    x"3E6F46F4",
    x"3E6F5F63",
    x"3E6F77D3",
    x"3E6F9043",
    x"3E6FA8B2",
    x"3E6FC121",
    x"3E6FD990",
    x"3E6FF1FF",
    x"3E700A6E",
    x"3E7022DD",
    x"3E703B4B",
    x"3E7053B9",
    x"3E706C28",
    x"3E708496",
    x"3E709D04",
    x"3E70B571",
    x"3E70CDDF",
    x"3E70E64C",
    x"3E70FEBA",
    x"3E711727",
    x"3E712F94",
    x"3E714801",
    x"3E71606E",
    x"3E7178DA",
    x"3E719147",
    x"3E71A9B3",
    x"3E71C21F",
    x"3E71DA8B",
    x"3E71F2F7",
    x"3E720B63",
    x"3E7223CE",
    x"3E723C3A",
    x"3E7254A5",
    x"3E726D10",
    x"3E72857B",
    x"3E729DE6",
    x"3E72B651",
    x"3E72CEBC",
    x"3E72E726",
    x"3E72FF90",
    x"3E7317FA",
    x"3E733064",
    x"3E7348CE",
    x"3E736138",
    x"3E7379A1",
    x"3E73920B",
    x"3E73AA74",
    x"3E73C2DD",
    x"3E73DB46",
    x"3E73F3AF",
    x"3E740C18",
    x"3E742480",
    x"3E743CE8",
    x"3E745551",
    x"3E746DB9",
    x"3E748621",
    x"3E749E88",
    x"3E74B6F0",
    x"3E74CF57",
    x"3E74E7BF",
    x"3E750026",
    x"3E75188D",
    x"3E7530F4",
    x"3E75495B",
    x"3E7561C1",
    x"3E757A28",
    x"3E75928E",
    x"3E75AAF4",
    x"3E75C35A",
    x"3E75DBC0",
    x"3E75F426",
    x"3E760C8B",
    x"3E7624F1",
    x"3E763D56",
    x"3E7655BB",
    x"3E766E20",
    x"3E768685",
    x"3E769EEA",
    x"3E76B74E",
    x"3E76CFB2",
    x"3E76E817",
    x"3E77007B",
    x"3E7718DF",
    x"3E773142",
    x"3E7749A6",
    x"3E77620A",
    x"3E777A6D",
    x"3E7792D0",
    x"3E77AB33",
    x"3E77C396",
    x"3E77DBF9",
    x"3E77F45B",
    x"3E780CBE",
    x"3E782520",
    x"3E783D82",
    x"3E7855E4",
    x"3E786E46",
    x"3E7886A8",
    x"3E789F09",
    x"3E78B76B",
    x"3E78CFCC",
    x"3E78E82D",
    x"3E79008E",
    x"3E7918EF",
    x"3E79314F",
    x"3E7949B0",
    x"3E796210",
    x"3E797A70",
    x"3E7992D0",
    x"3E79AB30",
    x"3E79C390",
    x"3E79DBF0",
    x"3E79F44F",
    x"3E7A0CAE",
    x"3E7A250D",
    x"3E7A3D6C",
    x"3E7A55CB",
    x"3E7A6E2A",
    x"3E7A8688",
    x"3E7A9EE7",
    x"3E7AB745",
    x"3E7ACFA3",
    x"3E7AE801",
    x"3E7B005F",
    x"3E7B18BC",
    x"3E7B311A",
    x"3E7B4977",
    x"3E7B61D4",
    x"3E7B7A31",
    x"3E7B928E",
    x"3E7BAAEB",
    x"3E7BC348",
    x"3E7BDBA4",
    x"3E7BF400",
    x"3E7C0C5C",
    x"3E7C24B8",
    x"3E7C3D14",
    x"3E7C5570",
    x"3E7C6DCB",
    x"3E7C8627",
    x"3E7C9E82",
    x"3E7CB6DD",
    x"3E7CCF38",
    x"3E7CE793",
    x"3E7CFFED",
    x"3E7D1848",
    x"3E7D30A2",
    x"3E7D48FC",
    x"3E7D6156",
    x"3E7D79B0",
    x"3E7D9209",
    x"3E7DAA63",
    x"3E7DC2BC",
    x"3E7DDB16",
    x"3E7DF36F",
    x"3E7E0BC8",
    x"3E7E2420",
    x"3E7E3C79",
    x"3E7E54D1",
    x"3E7E6D2A",
    x"3E7E8582",
    x"3E7E9DDA",
    x"3E7EB632",
    x"3E7ECE89",
    x"3E7EE6E1",
    x"3E7EFF38",
    x"3E7F178F",
    x"3E7F2FE7",
    x"3E7F483D",
    x"3E7F6094",
    x"3E7F78EB",
    x"3E7F9141",
    x"3E7FA998",
    x"3E7FC1EE",
    x"3E7FDA44",
    x"3E7FF29A",
    x"3E800578",
    x"3E8011A2",
    x"3E801DCD",
    x"3E8029F8",
    x"3E803622",
    x"3E80424D",
    x"3E804E77",
    x"3E805AA1",
    x"3E8066CC",
    x"3E8072F6",
    x"3E807F20",
    x"3E808B4A",
    x"3E809774",
    x"3E80A39E",
    x"3E80AFC7",
    x"3E80BBF1",
    x"3E80C81B",
    x"3E80D444",
    x"3E80E06E",
    x"3E80EC97",
    x"3E80F8C0",
    x"3E8104E9",
    x"3E811113",
    x"3E811D3C",
    x"3E812965",
    x"3E81358E",
    x"3E8141B6",
    x"3E814DDF",
    x"3E815A08",
    x"3E816630",
    x"3E817259",
    x"3E817E81",
    x"3E818AAA",
    x"3E8196D2",
    x"3E81A2FA",
    x"3E81AF22",
    x"3E81BB4A",
    x"3E81C772",
    x"3E81D39A",
    x"3E81DFC2",
    x"3E81EBEA",
    x"3E81F811",
    x"3E820439",
    x"3E821060",
    x"3E821C88",
    x"3E8228AF",
    x"3E8234D7",
    x"3E8240FE",
    x"3E824D25",
    x"3E82594C",
    x"3E826573",
    x"3E82719A",
    x"3E827DC0",
    x"3E8289E7",
    x"3E82960E",
    x"3E82A234",
    x"3E82AE5B",
    x"3E82BA81",
    x"3E82C6A8",
    x"3E82D2CE",
    x"3E82DEF4",
    x"3E82EB1A",
    x"3E82F740",
    x"3E830366",
    x"3E830F8C",
    x"3E831BB2",
    x"3E8327D7",
    x"3E8333FD",
    x"3E834022",
    x"3E834C48",
    x"3E83586D",
    x"3E836493",
    x"3E8370B8",
    x"3E837CDD",
    x"3E838902",
    x"3E839527",
    x"3E83A14C",
    x"3E83AD71",
    x"3E83B995",
    x"3E83C5BA",
    x"3E83D1DF",
    x"3E83DE03",
    x"3E83EA28",
    x"3E83F64C",
    x"3E840270",
    x"3E840E94",
    x"3E841AB8",
    x"3E8426DD",
    x"3E843300",
    x"3E843F24",
    x"3E844B48",
    x"3E84576C",
    x"3E84638F",
    x"3E846FB3",
    x"3E847BD6",
    x"3E8487FA",
    x"3E84941D",
    x"3E84A040",
    x"3E84AC64",
    x"3E84B887",
    x"3E84C4AA",
    x"3E84D0CC",
    x"3E84DCEF",
    x"3E84E912",
    x"3E84F535",
    x"3E850157",
    x"3E850D7A",
    x"3E85199C",
    x"3E8525BF",
    x"3E8531E1",
    x"3E853E03",
    x"3E854A25",
    x"3E855647",
    x"3E856269",
    x"3E856E8B",
    x"3E857AAD",
    x"3E8586CE",
    x"3E8592F0",
    x"3E859F12",
    x"3E85AB33",
    x"3E85B755",
    x"3E85C376",
    x"3E85CF97",
    x"3E85DBB8",
    x"3E85E7D9",
    x"3E85F3FA",
    x"3E86001B",
    x"3E860C3C",
    x"3E86185D",
    x"3E86247D",
    x"3E86309E",
    x"3E863CBE",
    x"3E8648DF",
    x"3E8654FF",
    x"3E86611F",
    x"3E866D40",
    x"3E867960",
    x"3E868580",
    x"3E8691A0",
    x"3E869DBF",
    x"3E86A9DF",
    x"3E86B5FF",
    x"3E86C21F",
    x"3E86CE3E",
    x"3E86DA5D",
    x"3E86E67D",
    x"3E86F29C",
    x"3E86FEBB",
    x"3E870ADA",
    x"3E8716F9",
    x"3E872318",
    x"3E872F37",
    x"3E873B56",
    x"3E874775",
    x"3E875393",
    x"3E875FB2",
    x"3E876BD0",
    x"3E8777EF",
    x"3E87840D",
    x"3E87902B",
    x"3E879C49",
    x"3E87A868",
    x"3E87B486",
    x"3E87C0A3",
    x"3E87CCC1",
    x"3E87D8DF",
    x"3E87E4FD",
    x"3E87F11A",
    x"3E87FD38",
    x"3E880955",
    x"3E881572",
    x"3E882190",
    x"3E882DAD",
    x"3E8839CA",
    x"3E8845E7",
    x"3E885204",
    x"3E885E21",
    x"3E886A3D",
    x"3E88765A",
    x"3E888277",
    x"3E888E93",
    x"3E889AB0",
    x"3E88A6CC",
    x"3E88B2E8",
    x"3E88BF04",
    x"3E88CB20",
    x"3E88D73C",
    x"3E88E358",
    x"3E88EF74",
    x"3E88FB90",
    x"3E8907AC",
    x"3E8913C7",
    x"3E891FE3",
    x"3E892BFE",
    x"3E893819",
    x"3E894435",
    x"3E895050",
    x"3E895C6B",
    x"3E896886",
    x"3E8974A1",
    x"3E8980BC",
    x"3E898CD7",
    x"3E8998F1",
    x"3E89A50C",
    x"3E89B126",
    x"3E89BD41",
    x"3E89C95B",
    x"3E89D575",
    x"3E89E190",
    x"3E89EDAA",
    x"3E89F9C4",
    x"3E8A05DE",
    x"3E8A11F7",
    x"3E8A1E11",
    x"3E8A2A2B",
    x"3E8A3645",
    x"3E8A425E",
    x"3E8A4E78",
    x"3E8A5A91",
    x"3E8A66AA",
    x"3E8A72C3",
    x"3E8A7EDC",
    x"3E8A8AF5",
    x"3E8A970E",
    x"3E8AA327",
    x"3E8AAF40",
    x"3E8ABB59",
    x"3E8AC771",
    x"3E8AD38A",
    x"3E8ADFA2",
    x"3E8AEBBB",
    x"3E8AF7D3",
    x"3E8B03EB",
    x"3E8B1003",
    x"3E8B1C1B",
    x"3E8B2833",
    x"3E8B344B",
    x"3E8B4063",
    x"3E8B4C7A",
    x"3E8B5892",
    x"3E8B64AA",
    x"3E8B70C1",
    x"3E8B7CD8",
    x"3E8B88F0",
    x"3E8B9507",
    x"3E8BA11E",
    x"3E8BAD35",
    x"3E8BB94C",
    x"3E8BC563",
    x"3E8BD179",
    x"3E8BDD90",
    x"3E8BE9A7",
    x"3E8BF5BD",
    x"3E8C01D4",
    x"3E8C0DEA",
    x"3E8C1A00",
    x"3E8C2616",
    x"3E8C322C",
    x"3E8C3E42",
    x"3E8C4A58",
    x"3E8C566E",
    x"3E8C6284",
    x"3E8C6E9A",
    x"3E8C7AAF",
    x"3E8C86C5",
    x"3E8C92DA",
    x"3E8C9EEF",
    x"3E8CAB05",
    x"3E8CB71A",
    x"3E8CC32F",
    x"3E8CCF44",
    x"3E8CDB59",
    x"3E8CE76D",
    x"3E8CF382",
    x"3E8CFF97",
    x"3E8D0BAB",
    x"3E8D17C0",
    x"3E8D23D4",
    x"3E8D2FE9",
    x"3E8D3BFD",
    x"3E8D4811",
    x"3E8D5425",
    x"3E8D6039",
    x"3E8D6C4D",
    x"3E8D7861",
    x"3E8D8474",
    x"3E8D9088",
    x"3E8D9C9B",
    x"3E8DA8AF",
    x"3E8DB4C2",
    x"3E8DC0D6",
    x"3E8DCCE9",
    x"3E8DD8FC",
    x"3E8DE50F",
    x"3E8DF122",
    x"3E8DFD35",
    x"3E8E0947",
    x"3E8E155A",
    x"3E8E216D",
    x"3E8E2D7F",
    x"3E8E3992",
    x"3E8E45A4",
    x"3E8E51B6",
    x"3E8E5DC8",
    x"3E8E69DB",
    x"3E8E75ED",
    x"3E8E81FE",
    x"3E8E8E10",
    x"3E8E9A22",
    x"3E8EA634",
    x"3E8EB245",
    x"3E8EBE57",
    x"3E8ECA68",
    x"3E8ED679",
    x"3E8EE28B",
    x"3E8EEE9C",
    x"3E8EFAAD",
    x"3E8F06BE",
    x"3E8F12CF",
    x"3E8F1EDF",
    x"3E8F2AF0",
    x"3E8F3701",
    x"3E8F4311",
    x"3E8F4F22",
    x"3E8F5B32",
    x"3E8F6742",
    x"3E8F7353",
    x"3E8F7F63",
    x"3E8F8B73",
    x"3E8F9783",
    x"3E8FA392",
    x"3E8FAFA2",
    x"3E8FBBB2",
    x"3E8FC7C1",
    x"3E8FD3D1",
    x"3E8FDFE0",
    x"3E8FEBF0",
    x"3E8FF7FF",
    x"3E90040E",
    x"3E90101D",
    x"3E901C2C",
    x"3E90283B",
    x"3E90344A",
    x"3E904059",
    x"3E904C67",
    x"3E905876",
    x"3E906484",
    x"3E907093",
    x"3E907CA1",
    x"3E9088AF",
    x"3E9094BD",
    x"3E90A0CB",
    x"3E90ACD9",
    x"3E90B8E7",
    x"3E90C4F5",
    x"3E90D102",
    x"3E90DD10",
    x"3E90E91D",
    x"3E90F52B",
    x"3E910138",
    x"3E910D45",
    x"3E911953",
    x"3E912560",
    x"3E91316D",
    x"3E913D79",
    x"3E914986",
    x"3E915593",
    x"3E9161A0",
    x"3E916DAC",
    x"3E9179B9",
    x"3E9185C5",
    x"3E9191D1",
    x"3E919DDD",
    x"3E91A9E9",
    x"3E91B5F5",
    x"3E91C201",
    x"3E91CE0D",
    x"3E91DA19",
    x"3E91E625",
    x"3E91F230",
    x"3E91FE3C",
    x"3E920A47",
    x"3E921652",
    x"3E92225E",
    x"3E922E69",
    x"3E923A74",
    x"3E92467F",
    x"3E92528A",
    x"3E925E94",
    x"3E926A9F",
    x"3E9276AA",
    x"3E9282B4",
    x"3E928EBF",
    x"3E929AC9",
    x"3E92A6D3",
    x"3E92B2DD",
    x"3E92BEE7",
    x"3E92CAF1",
    x"3E92D6FB",
    x"3E92E305",
    x"3E92EF0F",
    x"3E92FB18",
    x"3E930722",
    x"3E93132B",
    x"3E931F35",
    x"3E932B3E",
    x"3E933747",
    x"3E934350",
    x"3E934F59",
    x"3E935B62",
    x"3E93676B",
    x"3E937374",
    x"3E937F7D",
    x"3E938B85",
    x"3E93978E",
    x"3E93A396",
    x"3E93AF9E",
    x"3E93BBA6",
    x"3E93C7AF",
    x"3E93D3B7",
    x"3E93DFBF",
    x"3E93EBC6",
    x"3E93F7CE",
    x"3E9403D6",
    x"3E940FDD",
    x"3E941BE5",
    x"3E9427EC",
    x"3E9433F4",
    x"3E943FFB",
    x"3E944C02",
    x"3E945809",
    x"3E946410",
    x"3E947017",
    x"3E947C1E",
    x"3E948824",
    x"3E94942B",
    x"3E94A031",
    x"3E94AC38",
    x"3E94B83E",
    x"3E94C444",
    x"3E94D04B",
    x"3E94DC51",
    x"3E94E857",
    x"3E94F45D",
    x"3E950062",
    x"3E950C68",
    x"3E95186E",
    x"3E952473",
    x"3E953079",
    x"3E953C7E",
    x"3E954883",
    x"3E955488",
    x"3E95608D",
    x"3E956C92",
    x"3E957897",
    x"3E95849C",
    x"3E9590A1",
    x"3E959CA6",
    x"3E95A8AA",
    x"3E95B4AE",
    x"3E95C0B3",
    x"3E95CCB7",
    x"3E95D8BB",
    x"3E95E4BF",
    x"3E95F0C3",
    x"3E95FCC7",
    x"3E9608CB",
    x"3E9614CF",
    x"3E9620D2",
    x"3E962CD6",
    x"3E9638D9",
    x"3E9644DD",
    x"3E9650E0",
    x"3E965CE3",
    x"3E9668E6",
    x"3E9674E9",
    x"3E9680EC",
    x"3E968CEF",
    x"3E9698F2",
    x"3E96A4F4",
    x"3E96B0F7",
    x"3E96BCF9",
    x"3E96C8FC",
    x"3E96D4FE",
    x"3E96E100",
    x"3E96ED02",
    x"3E96F904",
    x"3E970506",
    x"3E971108",
    x"3E971D0A",
    x"3E97290B",
    x"3E97350D",
    x"3E97410E",
    x"3E974D10",
    x"3E975911",
    x"3E976512",
    x"3E977113",
    x"3E977D14",
    x"3E978915",
    x"3E979516",
    x"3E97A117",
    x"3E97AD17",
    x"3E97B918",
    x"3E97C518",
    x"3E97D119",
    x"3E97DD19",
    x"3E97E919",
    x"3E97F519",
    x"3E980119",
    x"3E980D19",
    x"3E981919",
    x"3E982519",
    x"3E983118",
    x"3E983D18",
    x"3E984917",
    x"3E985517",
    x"3E986116",
    x"3E986D15",
    x"3E987914",
    x"3E988513",
    x"3E989112",
    x"3E989D11",
    x"3E98A910",
    x"3E98B50E",
    x"3E98C10D",
    x"3E98CD0B",
    x"3E98D90A",
    x"3E98E508",
    x"3E98F106",
    x"3E98FD04",
    x"3E990902",
    x"3E991500",
    x"3E9920FE",
    x"3E992CFB",
    x"3E9938F9",
    x"3E9944F7",
    x"3E9950F4",
    x"3E995CF1",
    x"3E9968EE",
    x"3E9974EC",
    x"3E9980E9",
    x"3E998CE6",
    x"3E9998E3",
    x"3E99A4DF",
    x"3E99B0DC",
    x"3E99BCD9",
    x"3E99C8D5",
    x"3E99D4D1",
    x"3E99E0CE",
    x"3E99ECCA",
    x"3E99F8C6",
    x"3E9A04C2",
    x"3E9A10BE",
    x"3E9A1CBA",
    x"3E9A28B6",
    x"3E9A34B1",
    x"3E9A40AD",
    x"3E9A4CA8",
    x"3E9A58A4",
    x"3E9A649F",
    x"3E9A709A",
    x"3E9A7C95",
    x"3E9A8890",
    x"3E9A948B",
    x"3E9AA086",
    x"3E9AAC81",
    x"3E9AB87B",
    x"3E9AC476",
    x"3E9AD070",
    x"3E9ADC6B",
    x"3E9AE865",
    x"3E9AF45F",
    x"3E9B0059",
    x"3E9B0C53",
    x"3E9B184D",
    x"3E9B2447",
    x"3E9B3041",
    x"3E9B3C3A",
    x"3E9B4834",
    x"3E9B542D",
    x"3E9B6027",
    x"3E9B6C20",
    x"3E9B7819",
    x"3E9B8412",
    x"3E9B900B",
    x"3E9B9C04",
    x"3E9BA7FD",
    x"3E9BB3F5",
    x"3E9BBFEE",
    x"3E9BCBE6",
    x"3E9BD7DF",
    x"3E9BE3D7",
    x"3E9BEFCF",
    x"3E9BFBC7",
    x"3E9C07BF",
    x"3E9C13B7",
    x"3E9C1FAF",
    x"3E9C2BA7",
    x"3E9C379E",
    x"3E9C4396",
    x"3E9C4F8D",
    x"3E9C5B85",
    x"3E9C677C",
    x"3E9C7373",
    x"3E9C7F6A",
    x"3E9C8B61",
    x"3E9C9758",
    x"3E9CA34F",
    x"3E9CAF46",
    x"3E9CBB3C",
    x"3E9CC733",
    x"3E9CD329",
    x"3E9CDF20",
    x"3E9CEB16",
    x"3E9CF70C",
    x"3E9D0302",
    x"3E9D0EF8",
    x"3E9D1AEE",
    x"3E9D26E3",
    x"3E9D32D9",
    x"3E9D3ECF",
    x"3E9D4AC4",
    x"3E9D56BA",
    x"3E9D62AF",
    x"3E9D6EA4",
    x"3E9D7A99",
    x"3E9D868E",
    x"3E9D9283",
    x"3E9D9E78",
    x"3E9DAA6D",
    x"3E9DB661",
    x"3E9DC256",
    x"3E9DCE4A",
    x"3E9DDA3E",
    x"3E9DE633",
    x"3E9DF227",
    x"3E9DFE1B",
    x"3E9E0A0F",
    x"3E9E1603",
    x"3E9E21F6",
    x"3E9E2DEA",
    x"3E9E39DE",
    x"3E9E45D1",
    x"3E9E51C4",
    x"3E9E5DB8",
    x"3E9E69AB",
    x"3E9E759E",
    x"3E9E8191",
    x"3E9E8D84",
    x"3E9E9977",
    x"3E9EA569",
    x"3E9EB15C",
    x"3E9EBD4F",
    x"3E9EC941",
    x"3E9ED533",
    x"3E9EE126",
    x"3E9EED18",
    x"3E9EF90A",
    x"3E9F04FC",
    x"3E9F10EE",
    x"3E9F1CDF",
    x"3E9F28D1",
    x"3E9F34C3",
    x"3E9F40B4",
    x"3E9F4CA5",
    x"3E9F5897",
    x"3E9F6488",
    x"3E9F7079",
    x"3E9F7C6A",
    x"3E9F885B",
    x"3E9F944C",
    x"3E9FA03C",
    x"3E9FAC2D",
    x"3E9FB81D",
    x"3E9FC40E",
    x"3E9FCFFE",
    x"3E9FDBEE",
    x"3E9FE7DE",
    x"3E9FF3CE",
    x"3E9FFFBE",
    x"3EA00BAE",
    x"3EA0179E",
    x"3EA0238E",
    x"3EA02F7D",
    x"3EA03B6D",
    x"3EA0475C",
    x"3EA0534B",
    x"3EA05F3A",
    x"3EA06B29",
    x"3EA07718",
    x"3EA08307",
    x"3EA08EF6",
    x"3EA09AE5",
    x"3EA0A6D3",
    x"3EA0B2C2",
    x"3EA0BEB0",
    x"3EA0CA9E",
    x"3EA0D68D",
    x"3EA0E27B",
    x"3EA0EE69",
    x"3EA0FA57",
    x"3EA10644",
    x"3EA11232",
    x"3EA11E20",
    x"3EA12A0D",
    x"3EA135FB",
    x"3EA141E8",
    x"3EA14DD5",
    x"3EA159C2",
    x"3EA165AF",
    x"3EA1719C",
    x"3EA17D89",
    x"3EA18976",
    x"3EA19562",
    x"3EA1A14F",
    x"3EA1AD3B",
    x"3EA1B928",
    x"3EA1C514",
    x"3EA1D100",
    x"3EA1DCEC",
    x"3EA1E8D8",
    x"3EA1F4C4",
    x"3EA200B0",
    x"3EA20C9B",
    x"3EA21887",
    x"3EA22472",
    x"3EA2305E",
    x"3EA23C49",
    x"3EA24834",
    x"3EA2541F",
    x"3EA2600A",
    x"3EA26BF5",
    x"3EA277E0",
    x"3EA283CB",
    x"3EA28FB5",
    x"3EA29BA0",
    x"3EA2A78A",
    x"3EA2B374",
    x"3EA2BF5E",
    x"3EA2CB49",
    x"3EA2D733",
    x"3EA2E31C",
    x"3EA2EF06",
    x"3EA2FAF0",
    x"3EA306DA",
    x"3EA312C3",
    x"3EA31EAD",
    x"3EA32A96",
    x"3EA3367F",
    x"3EA34268",
    x"3EA34E51",
    x"3EA35A3A",
    x"3EA36623",
    x"3EA3720C",
    x"3EA37DF4",
    x"3EA389DD",
    x"3EA395C5",
    x"3EA3A1AD",
    x"3EA3AD96",
    x"3EA3B97E",
    x"3EA3C566",
    x"3EA3D14E",
    x"3EA3DD36",
    x"3EA3E91D",
    x"3EA3F505",
    x"3EA400ED",
    x"3EA40CD4",
    x"3EA418BB",
    x"3EA424A3",
    x"3EA4308A",
    x"3EA43C71",
    x"3EA44858",
    x"3EA4543F",
    x"3EA46025",
    x"3EA46C0C",
    x"3EA477F2",
    x"3EA483D9",
    x"3EA48FBF",
    x"3EA49BA6",
    x"3EA4A78C",
    x"3EA4B372",
    x"3EA4BF58",
    x"3EA4CB3E",
    x"3EA4D723",
    x"3EA4E309",
    x"3EA4EEEE",
    x"3EA4FAD4",
    x"3EA506B9",
    x"3EA5129F",
    x"3EA51E84",
    x"3EA52A69",
    x"3EA5364E",
    x"3EA54233",
    x"3EA54E17",
    x"3EA559FC",
    x"3EA565E1",
    x"3EA571C5",
    x"3EA57DA9",
    x"3EA5898E",
    x"3EA59572",
    x"3EA5A156",
    x"3EA5AD3A",
    x"3EA5B91E",
    x"3EA5C501",
    x"3EA5D0E5",
    x"3EA5DCC9",
    x"3EA5E8AC",
    x"3EA5F48F",
    x"3EA60073",
    x"3EA60C56",
    x"3EA61839",
    x"3EA6241C",
    x"3EA62FFF",
    x"3EA63BE2",
    x"3EA647C4",
    x"3EA653A7",
    x"3EA65F89",
    x"3EA66B6C",
    x"3EA6774E",
    x"3EA68330",
    x"3EA68F12",
    x"3EA69AF4",
    x"3EA6A6D6",
    x"3EA6B2B8",
    x"3EA6BE99",
    x"3EA6CA7B",
    x"3EA6D65C",
    x"3EA6E23E",
    x"3EA6EE1F",
    x"3EA6FA00",
    x"3EA705E1",
    x"3EA711C2",
    x"3EA71DA3",
    x"3EA72984",
    x"3EA73564",
    x"3EA74145",
    x"3EA74D25",
    x"3EA75906",
    x"3EA764E6",
    x"3EA770C6",
    x"3EA77CA6",
    x"3EA78886",
    x"3EA79466",
    x"3EA7A046",
    x"3EA7AC25",
    x"3EA7B805",
    x"3EA7C3E4",
    x"3EA7CFC4",
    x"3EA7DBA3",
    x"3EA7E782",
    x"3EA7F361",
    x"3EA7FF40",
    x"3EA80B1F",
    x"3EA816FE",
    x"3EA822DC",
    x"3EA82EBB",
    x"3EA83A99",
    x"3EA84678",
    x"3EA85256",
    x"3EA85E34",
    x"3EA86A12",
    x"3EA875F0",
    x"3EA881CE",
    x"3EA88DAB",
    x"3EA89989",
    x"3EA8A567",
    x"3EA8B144",
    x"3EA8BD21",
    x"3EA8C8FE",
    x"3EA8D4DC",
    x"3EA8E0B9",
    x"3EA8EC95",
    x"3EA8F872",
    x"3EA9044F",
    x"3EA9102C",
    x"3EA91C08",
    x"3EA927E5",
    x"3EA933C1",
    x"3EA93F9D",
    x"3EA94B79",
    x"3EA95755",
    x"3EA96331",
    x"3EA96F0D",
    x"3EA97AE8",
    x"3EA986C4",
    x"3EA992A0",
    x"3EA99E7B",
    x"3EA9AA56",
    x"3EA9B631",
    x"3EA9C20C",
    x"3EA9CDE7",
    x"3EA9D9C2",
    x"3EA9E59D",
    x"3EA9F178",
    x"3EA9FD52",
    x"3EAA092D",
    x"3EAA1507",
    x"3EAA20E1",
    x"3EAA2CBB",
    x"3EAA3895",
    x"3EAA446F",
    x"3EAA5049",
    x"3EAA5C23",
    x"3EAA67FD",
    x"3EAA73D6",
    x"3EAA7FB0",
    x"3EAA8B89",
    x"3EAA9762",
    x"3EAAA33B",
    x"3EAAAF14",
    x"3EAABAED",
    x"3EAAC6C6",
    x"3EAAD29F",
    x"3EAADE77",
    x"3EAAEA50",
    x"3EAAF628",
    x"3EAB0201",
    x"3EAB0DD9",
    x"3EAB19B1",
    x"3EAB2589",
    x"3EAB3161",
    x"3EAB3D39",
    x"3EAB4910",
    x"3EAB54E8",
    x"3EAB60BF",
    x"3EAB6C97",
    x"3EAB786E",
    x"3EAB8445",
    x"3EAB901C",
    x"3EAB9BF3",
    x"3EABA7CA",
    x"3EABB3A1",
    x"3EABBF77",
    x"3EABCB4E",
    x"3EABD724",
    x"3EABE2FB",
    x"3EABEED1",
    x"3EABFAA7",
    x"3EAC067D",
    x"3EAC1253",
    x"3EAC1E29",
    x"3EAC29FF",
    x"3EAC35D4",
    x"3EAC41AA",
    x"3EAC4D7F",
    x"3EAC5954",
    x"3EAC652A",
    x"3EAC70FF",
    x"3EAC7CD4",
    x"3EAC88A9",
    x"3EAC947D",
    x"3EACA052",
    x"3EACAC27",
    x"3EACB7FB",
    x"3EACC3CF",
    x"3EACCFA4",
    x"3EACDB78",
    x"3EACE74C",
    x"3EACF320",
    x"3EACFEF4",
    x"3EAD0AC7",
    x"3EAD169B",
    x"3EAD226F",
    x"3EAD2E42",
    x"3EAD3A15",
    x"3EAD45E9",
    x"3EAD51BC",
    x"3EAD5D8F",
    x"3EAD6962",
    x"3EAD7534",
    x"3EAD8107",
    x"3EAD8CDA",
    x"3EAD98AC",
    x"3EADA47F",
    x"3EADB051",
    x"3EADBC23",
    x"3EADC7F5",
    x"3EADD3C7",
    x"3EADDF99",
    x"3EADEB6B",
    x"3EADF73C",
    x"3EAE030E",
    x"3EAE0EDF",
    x"3EAE1AB1",
    x"3EAE2682",
    x"3EAE3253",
    x"3EAE3E24",
    x"3EAE49F5",
    x"3EAE55C6",
    x"3EAE6197",
    x"3EAE6D67",
    x"3EAE7938",
    x"3EAE8508",
    x"3EAE90D8",
    x"3EAE9CA8",
    x"3EAEA879",
    x"3EAEB449",
    x"3EAEC018",
    x"3EAECBE8",
    x"3EAED7B8",
    x"3EAEE387",
    x"3EAEEF57",
    x"3EAEFB26",
    x"3EAF06F5",
    x"3EAF12C5",
    x"3EAF1E94",
    x"3EAF2A62",
    x"3EAF3631",
    x"3EAF4200",
    x"3EAF4DCF",
    x"3EAF599D",
    x"3EAF656B",
    x"3EAF713A",
    x"3EAF7D08",
    x"3EAF88D6",
    x"3EAF94A4",
    x"3EAFA072",
    x"3EAFAC40",
    x"3EAFB80D",
    x"3EAFC3DB",
    x"3EAFCFA8",
    x"3EAFDB76",
    x"3EAFE743",
    x"3EAFF310",
    x"3EAFFEDD",
    x"3EB00AAA",
    x"3EB01677",
    x"3EB02243",
    x"3EB02E10",
    x"3EB039DC",
    x"3EB045A9",
    x"3EB05175",
    x"3EB05D41",
    x"3EB0690D",
    x"3EB074D9",
    x"3EB080A5",
    x"3EB08C71",
    x"3EB0983C",
    x"3EB0A408",
    x"3EB0AFD3",
    x"3EB0BB9F",
    x"3EB0C76A",
    x"3EB0D335",
    x"3EB0DF00",
    x"3EB0EACB",
    x"3EB0F696",
    x"3EB10260",
    x"3EB10E2B",
    x"3EB119F5",
    x"3EB125C0",
    x"3EB1318A",
    x"3EB13D54",
    x"3EB1491E",
    x"3EB154E8",
    x"3EB160B2",
    x"3EB16C7C",
    x"3EB17845",
    x"3EB1840F",
    x"3EB18FD8",
    x"3EB19BA1",
    x"3EB1A76B",
    x"3EB1B334",
    x"3EB1BEFD",
    x"3EB1CAC5",
    x"3EB1D68E",
    x"3EB1E257",
    x"3EB1EE1F",
    x"3EB1F9E8",
    x"3EB205B0",
    x"3EB21178",
    x"3EB21D41",
    x"3EB22909",
    x"3EB234D0",
    x"3EB24098",
    x"3EB24C60",
    x"3EB25827",
    x"3EB263EF",
    x"3EB26FB6",
    x"3EB27B7E",
    x"3EB28745",
    x"3EB2930C",
    x"3EB29ED3",
    x"3EB2AA99",
    x"3EB2B660",
    x"3EB2C227",
    x"3EB2CDED",
    x"3EB2D9B4",
    x"3EB2E57A",
    x"3EB2F140",
    x"3EB2FD06",
    x"3EB308CC",
    x"3EB31492",
    x"3EB32058",
    x"3EB32C1D",
    x"3EB337E3",
    x"3EB343A8",
    x"3EB34F6E",
    x"3EB35B33",
    x"3EB366F8",
    x"3EB372BD",
    x"3EB37E82",
    x"3EB38A47",
    x"3EB3960B",
    x"3EB3A1D0",
    x"3EB3AD94",
    x"3EB3B959",
    x"3EB3C51D",
    x"3EB3D0E1",
    x"3EB3DCA5",
    x"3EB3E869",
    x"3EB3F42D",
    x"3EB3FFF0",
    x"3EB40BB4",
    x"3EB41777",
    x"3EB4233B",
    x"3EB42EFE",
    x"3EB43AC1",
    x"3EB44684",
    x"3EB45247",
    x"3EB45E0A",
    x"3EB469CD",
    x"3EB4758F",
    x"3EB48152",
    x"3EB48D14",
    x"3EB498D6",
    x"3EB4A499",
    x"3EB4B05B",
    x"3EB4BC1D",
    x"3EB4C7DE",
    x"3EB4D3A0",
    x"3EB4DF62",
    x"3EB4EB23",
    x"3EB4F6E5",
    x"3EB502A6",
    x"3EB50E67",
    x"3EB51A28",
    x"3EB525E9",
    x"3EB531AA",
    x"3EB53D6B",
    x"3EB5492B",
    x"3EB554EC",
    x"3EB560AC",
    x"3EB56C6D",
    x"3EB5782D",
    x"3EB583ED",
    x"3EB58FAD",
    x"3EB59B6D",
    x"3EB5A72D",
    x"3EB5B2EC",
    x"3EB5BEAC",
    x"3EB5CA6B",
    x"3EB5D62B",
    x"3EB5E1EA",
    x"3EB5EDA9",
    x"3EB5F968",
    x"3EB60527",
    x"3EB610E6",
    x"3EB61CA4",
    x"3EB62863",
    x"3EB63421",
    x"3EB63FE0",
    x"3EB64B9E",
    x"3EB6575C",
    x"3EB6631A",
    x"3EB66ED8",
    x"3EB67A96",
    x"3EB68653",
    x"3EB69211",
    x"3EB69DCE",
    x"3EB6A98C",
    x"3EB6B549",
    x"3EB6C106",
    x"3EB6CCC3",
    x"3EB6D880",
    x"3EB6E43D",
    x"3EB6EFFA",
    x"3EB6FBB6",
    x"3EB70773",
    x"3EB7132F",
    x"3EB71EEB",
    x"3EB72AA7",
    x"3EB73663",
    x"3EB7421F",
    x"3EB74DDB",
    x"3EB75997",
    x"3EB76552",
    x"3EB7710E",
    x"3EB77CC9",
    x"3EB78884",
    x"3EB79440",
    x"3EB79FFB",
    x"3EB7ABB6",
    x"3EB7B770",
    x"3EB7C32B",
    x"3EB7CEE6",
    x"3EB7DAA0",
    x"3EB7E65B",
    x"3EB7F215",
    x"3EB7FDCF",
    x"3EB80989",
    x"3EB81543",
    x"3EB820FD",
    x"3EB82CB6",
    x"3EB83870",
    x"3EB8442A",
    x"3EB84FE3",
    x"3EB85B9C",
    x"3EB86755",
    x"3EB8730E",
    x"3EB87EC7",
    x"3EB88A80",
    x"3EB89639",
    x"3EB8A1F1",
    x"3EB8ADAA",
    x"3EB8B962",
    x"3EB8C51B",
    x"3EB8D0D3",
    x"3EB8DC8B",
    x"3EB8E843",
    x"3EB8F3FA",
    x"3EB8FFB2",
    x"3EB90B6A",
    x"3EB91721",
    x"3EB922D9",
    x"3EB92E90",
    x"3EB93A47",
    x"3EB945FE",
    x"3EB951B5",
    x"3EB95D6C",
    x"3EB96923",
    x"3EB974D9",
    x"3EB98090",
    x"3EB98C46",
    x"3EB997FC",
    x"3EB9A3B2",
    x"3EB9AF68",
    x"3EB9BB1E",
    x"3EB9C6D4",
    x"3EB9D28A",
    x"3EB9DE3F",
    x"3EB9E9F5",
    x"3EB9F5AA",
    x"3EBA015F",
    x"3EBA0D15",
    x"3EBA18CA",
    x"3EBA247F",
    x"3EBA3033",
    x"3EBA3BE8",
    x"3EBA479D",
    x"3EBA5351",
    x"3EBA5F05",
    x"3EBA6ABA",
    x"3EBA766E",
    x"3EBA8222",
    x"3EBA8DD6",
    x"3EBA9989",
    x"3EBAA53D",
    x"3EBAB0F1",
    x"3EBABCA4",
    x"3EBAC857",
    x"3EBAD40B",
    x"3EBADFBE",
    x"3EBAEB71",
    x"3EBAF724",
    x"3EBB02D6",
    x"3EBB0E89",
    x"3EBB1A3C",
    x"3EBB25EE",
    x"3EBB31A0",
    x"3EBB3D53",
    x"3EBB4905",
    x"3EBB54B7",
    x"3EBB6069",
    x"3EBB6C1A",
    x"3EBB77CC",
    x"3EBB837E",
    x"3EBB8F2F",
    x"3EBB9AE0",
    x"3EBBA692",
    x"3EBBB243",
    x"3EBBBDF4",
    x"3EBBC9A4",
    x"3EBBD555",
    x"3EBBE106",
    x"3EBBECB6",
    x"3EBBF867",
    x"3EBC0417",
    x"3EBC0FC7",
    x"3EBC1B77",
    x"3EBC2727",
    x"3EBC32D7",
    x"3EBC3E87",
    x"3EBC4A36",
    x"3EBC55E6",
    x"3EBC6195",
    x"3EBC6D45",
    x"3EBC78F4",
    x"3EBC84A3",
    x"3EBC9052",
    x"3EBC9C00",
    x"3EBCA7AF",
    x"3EBCB35E",
    x"3EBCBF0C",
    x"3EBCCABB",
    x"3EBCD669",
    x"3EBCE217",
    x"3EBCEDC5",
    x"3EBCF973",
    x"3EBD0521",
    x"3EBD10CE",
    x"3EBD1C7C",
    x"3EBD2829",
    x"3EBD33D7",
    x"3EBD3F84",
    x"3EBD4B31",
    x"3EBD56DE",
    x"3EBD628B",
    x"3EBD6E38",
    x"3EBD79E4",
    x"3EBD8591",
    x"3EBD913D",
    x"3EBD9CEA",
    x"3EBDA896",
    x"3EBDB442",
    x"3EBDBFEE",
    x"3EBDCB9A",
    x"3EBDD746",
    x"3EBDE2F1",
    x"3EBDEE9D",
    x"3EBDFA48",
    x"3EBE05F3",
    x"3EBE119E",
    x"3EBE1D4A",
    x"3EBE28F4",
    x"3EBE349F",
    x"3EBE404A",
    x"3EBE4BF5",
    x"3EBE579F",
    x"3EBE6349",
    x"3EBE6EF4",
    x"3EBE7A9E",
    x"3EBE8648",
    x"3EBE91F2",
    x"3EBE9D9C",
    x"3EBEA945",
    x"3EBEB4EF",
    x"3EBEC098",
    x"3EBECC42",
    x"3EBED7EB",
    x"3EBEE394",
    x"3EBEEF3D",
    x"3EBEFAE6",
    x"3EBF068F",
    x"3EBF1237",
    x"3EBF1DE0",
    x"3EBF2988",
    x"3EBF3530",
    x"3EBF40D9",
    x"3EBF4C81",
    x"3EBF5829",
    x"3EBF63D0",
    x"3EBF6F78",
    x"3EBF7B20",
    x"3EBF86C7",
    x"3EBF926F",
    x"3EBF9E16",
    x"3EBFA9BD",
    x"3EBFB564",
    x"3EBFC10B",
    x"3EBFCCB2",
    x"3EBFD858",
    x"3EBFE3FF",
    x"3EBFEFA5",
    x"3EBFFB4C",
    x"3EC006F2",
    x"3EC01298",
    x"3EC01E3E",
    x"3EC029E4",
    x"3EC0358A",
    x"3EC0412F",
    x"3EC04CD5",
    x"3EC0587A",
    x"3EC06420",
    x"3EC06FC5",
    x"3EC07B6A",
    x"3EC0870F",
    x"3EC092B4",
    x"3EC09E58",
    x"3EC0A9FD",
    x"3EC0B5A1",
    x"3EC0C146",
    x"3EC0CCEA",
    x"3EC0D88E",
    x"3EC0E432",
    x"3EC0EFD6",
    x"3EC0FB7A",
    x"3EC1071E",
    x"3EC112C1",
    x"3EC11E64",
    x"3EC12A08",
    x"3EC135AB",
    x"3EC1414E",
    x"3EC14CF1",
    x"3EC15894",
    x"3EC16437",
    x"3EC16FD9",
    x"3EC17B7C",
    x"3EC1871E",
    x"3EC192C0",
    x"3EC19E63",
    x"3EC1AA05",
    x"3EC1B5A7",
    x"3EC1C148",
    x"3EC1CCEA",
    x"3EC1D88C",
    x"3EC1E42D",
    x"3EC1EFCE",
    x"3EC1FB70",
    x"3EC20711",
    x"3EC212B2",
    x"3EC21E53",
    x"3EC229F3",
    x"3EC23594",
    x"3EC24135",
    x"3EC24CD5",
    x"3EC25875",
    x"3EC26415",
    x"3EC26FB5",
    x"3EC27B55",
    x"3EC286F5",
    x"3EC29295",
    x"3EC29E34",
    x"3EC2A9D4",
    x"3EC2B573",
    x"3EC2C112",
    x"3EC2CCB2",
    x"3EC2D851",
    x"3EC2E3EF",
    x"3EC2EF8E",
    x"3EC2FB2D",
    x"3EC306CB",
    x"3EC3126A",
    x"3EC31E08",
    x"3EC329A6",
    x"3EC33544",
    x"3EC340E2",
    x"3EC34C80",
    x"3EC3581E",
    x"3EC363BB",
    x"3EC36F59",
    x"3EC37AF6",
    x"3EC38693",
    x"3EC39231",
    x"3EC39DCE",
    x"3EC3A96A",
    x"3EC3B507",
    x"3EC3C0A4",
    x"3EC3CC40",
    x"3EC3D7DD",
    x"3EC3E379",
    x"3EC3EF15",
    x"3EC3FAB1",
    x"3EC4064D",
    x"3EC411E9",
    x"3EC41D85",
    x"3EC42920",
    x"3EC434BC",
    x"3EC44057",
    x"3EC44BF2",
    x"3EC4578D",
    x"3EC46328",
    x"3EC46EC3",
    x"3EC47A5E",
    x"3EC485F9",
    x"3EC49193",
    x"3EC49D2E",
    x"3EC4A8C8",
    x"3EC4B462",
    x"3EC4BFFC",
    x"3EC4CB96",
    x"3EC4D730",
    x"3EC4E2C9",
    x"3EC4EE63",
    x"3EC4F9FD",
    x"3EC50596",
    x"3EC5112F",
    x"3EC51CC8",
    x"3EC52861",
    x"3EC533FA",
    x"3EC53F93",
    x"3EC54B2B",
    x"3EC556C4",
    x"3EC5625C",
    x"3EC56DF4",
    x"3EC5798D",
    x"3EC58525",
    x"3EC590BD",
    x"3EC59C54",
    x"3EC5A7EC",
    x"3EC5B384",
    x"3EC5BF1B",
    x"3EC5CAB2",
    x"3EC5D649",
    x"3EC5E1E1",
    x"3EC5ED77",
    x"3EC5F90E",
    x"3EC604A5",
    x"3EC6103C",
    x"3EC61BD2",
    x"3EC62768",
    x"3EC632FF",
    x"3EC63E95",
    x"3EC64A2B",
    x"3EC655C1",
    x"3EC66156",
    x"3EC66CEC",
    x"3EC67882",
    x"3EC68417",
    x"3EC68FAC",
    x"3EC69B41",
    x"3EC6A6D6",
    x"3EC6B26B",
    x"3EC6BE00",
    x"3EC6C995",
    x"3EC6D529",
    x"3EC6E0BE",
    x"3EC6EC52",
    x"3EC6F7E6",
    x"3EC7037B",
    x"3EC70F0E",
    x"3EC71AA2",
    x"3EC72636",
    x"3EC731CA",
    x"3EC73D5D",
    x"3EC748F0",
    x"3EC75484",
    x"3EC76017",
    x"3EC76BAA",
    x"3EC7773D",
    x"3EC782D0",
    x"3EC78E62",
    x"3EC799F5",
    x"3EC7A587",
    x"3EC7B119",
    x"3EC7BCAC",
    x"3EC7C83E",
    x"3EC7D3CF",
    x"3EC7DF61",
    x"3EC7EAF3",
    x"3EC7F685",
    x"3EC80216",
    x"3EC80DA7",
    x"3EC81938",
    x"3EC824CA",
    x"3EC8305B",
    x"3EC83BEB",
    x"3EC8477C",
    x"3EC8530D",
    x"3EC85E9D",
    x"3EC86A2D",
    x"3EC875BE",
    x"3EC8814E",
    x"3EC88CDE",
    x"3EC8986E",
    x"3EC8A3FD",
    x"3EC8AF8D",
    x"3EC8BB1D",
    x"3EC8C6AC",
    x"3EC8D23B",
    x"3EC8DDCA",
    x"3EC8E959",
    x"3EC8F4E8",
    x"3EC90077",
    x"3EC90C06",
    x"3EC91794",
    x"3EC92323",
    x"3EC92EB1",
    x"3EC93A3F",
    x"3EC945CD",
    x"3EC9515B",
    x"3EC95CE9",
    x"3EC96877",
    x"3EC97404",
    x"3EC97F92",
    x"3EC98B1F",
    x"3EC996AC",
    x"3EC9A239",
    x"3EC9ADC6",
    x"3EC9B953",
    x"3EC9C4E0",
    x"3EC9D06C",
    x"3EC9DBF9",
    x"3EC9E785",
    x"3EC9F312",
    x"3EC9FE9E",
    x"3ECA0A2A",
    x"3ECA15B5",
    x"3ECA2141",
    x"3ECA2CCD",
    x"3ECA3858",
    x"3ECA43E4",
    x"3ECA4F6F",
    x"3ECA5AFA",
    x"3ECA6685",
    x"3ECA7210",
    x"3ECA7D9B",
    x"3ECA8925",
    x"3ECA94B0",
    x"3ECAA03A",
    x"3ECAABC5",
    x"3ECAB74F",
    x"3ECAC2D9",
    x"3ECACE63",
    x"3ECAD9ED",
    x"3ECAE576",
    x"3ECAF100",
    x"3ECAFC89",
    x"3ECB0813",
    x"3ECB139C",
    x"3ECB1F25",
    x"3ECB2AAE",
    x"3ECB3637",
    x"3ECB41BF",
    x"3ECB4D48",
    x"3ECB58D0",
    x"3ECB6459",
    x"3ECB6FE1",
    x"3ECB7B69",
    x"3ECB86F1",
    x"3ECB9279",
    x"3ECB9E00",
    x"3ECBA988",
    x"3ECBB50F",
    x"3ECBC097",
    x"3ECBCC1E",
    x"3ECBD7A5",
    x"3ECBE32C",
    x"3ECBEEB3",
    x"3ECBFA3A",
    x"3ECC05C0",
    x"3ECC1147",
    x"3ECC1CCD",
    x"3ECC2853",
    x"3ECC33DA",
    x"3ECC3F60",
    x"3ECC4AE5",
    x"3ECC566B",
    x"3ECC61F1",
    x"3ECC6D76",
    x"3ECC78FC",
    x"3ECC8481",
    x"3ECC9006",
    x"3ECC9B8B",
    x"3ECCA710",
    x"3ECCB295",
    x"3ECCBE19",
    x"3ECCC99E",
    x"3ECCD522",
    x"3ECCE0A7",
    x"3ECCEC2B",
    x"3ECCF7AF",
    x"3ECD0333",
    x"3ECD0EB6",
    x"3ECD1A3A",
    x"3ECD25BE",
    x"3ECD3141",
    x"3ECD3CC4",
    x"3ECD4847",
    x"3ECD53CA",
    x"3ECD5F4D",
    x"3ECD6AD0",
    x"3ECD7653",
    x"3ECD81D5",
    x"3ECD8D58",
    x"3ECD98DA",
    x"3ECDA45C",
    x"3ECDAFDE",
    x"3ECDBB60",
    x"3ECDC6E2",
    x"3ECDD264",
    x"3ECDDDE5",
    x"3ECDE967",
    x"3ECDF4E8",
    x"3ECE0069",
    x"3ECE0BEA",
    x"3ECE176B",
    x"3ECE22EC",
    x"3ECE2E6D",
    x"3ECE39ED",
    x"3ECE456E",
    x"3ECE50EE",
    x"3ECE5C6E",
    x"3ECE67EE",
    x"3ECE736E",
    x"3ECE7EEE",
    x"3ECE8A6E",
    x"3ECE95ED",
    x"3ECEA16D",
    x"3ECEACEC",
    x"3ECEB86B",
    x"3ECEC3EA",
    x"3ECECF69",
    x"3ECEDAE8",
    x"3ECEE667",
    x"3ECEF1E5",
    x"3ECEFD64",
    x"3ECF08E2",
    x"3ECF1460",
    x"3ECF1FDE",
    x"3ECF2B5C",
    x"3ECF36DA",
    x"3ECF4258",
    x"3ECF4DD5",
    x"3ECF5953",
    x"3ECF64D0",
    x"3ECF704D",
    x"3ECF7BCA",
    x"3ECF8747",
    x"3ECF92C4",
    x"3ECF9E41",
    x"3ECFA9BD",
    x"3ECFB53A",
    x"3ECFC0B6",
    x"3ECFCC32",
    x"3ECFD7AE",
    x"3ECFE32A",
    x"3ECFEEA6",
    x"3ECFFA22",
    x"3ED0059D",
    x"3ED01119",
    x"3ED01C94",
    x"3ED0280F",
    x"3ED0338A",
    x"3ED03F05",
    x"3ED04A80",
    x"3ED055FB",
    x"3ED06175",
    x"3ED06CF0",
    x"3ED0786A",
    x"3ED083E4",
    x"3ED08F5E",
    x"3ED09AD8",
    x"3ED0A652",
    x"3ED0B1CC",
    x"3ED0BD45",
    x"3ED0C8BF",
    x"3ED0D438",
    x"3ED0DFB1",
    x"3ED0EB2A",
    x"3ED0F6A3",
    x"3ED1021C",
    x"3ED10D95",
    x"3ED1190D",
    x"3ED12485",
    x"3ED12FFE",
    x"3ED13B76",
    x"3ED146EE",
    x"3ED15266",
    x"3ED15DDE",
    x"3ED16955",
    x"3ED174CD",
    x"3ED18044",
    x"3ED18BBC",
    x"3ED19733",
    x"3ED1A2AA",
    x"3ED1AE21",
    x"3ED1B998",
    x"3ED1C50E",
    x"3ED1D085",
    x"3ED1DBFB",
    x"3ED1E771",
    x"3ED1F2E8",
    x"3ED1FE5E",
    x"3ED209D3",
    x"3ED21549",
    x"3ED220BF",
    x"3ED22C34",
    x"3ED237AA",
    x"3ED2431F",
    x"3ED24E94",
    x"3ED25A09",
    x"3ED2657E",
    x"3ED270F3",
    x"3ED27C68",
    x"3ED287DC",
    x"3ED29350",
    x"3ED29EC5",
    x"3ED2AA39",
    x"3ED2B5AD",
    x"3ED2C121",
    x"3ED2CC94",
    x"3ED2D808",
    x"3ED2E37C",
    x"3ED2EEEF",
    x"3ED2FA62",
    x"3ED305D5",
    x"3ED31148",
    x"3ED31CBB",
    x"3ED3282E",
    x"3ED333A0",
    x"3ED33F13",
    x"3ED34A85",
    x"3ED355F7",
    x"3ED3616A",
    x"3ED36CDB",
    x"3ED3784D",
    x"3ED383BF",
    x"3ED38F31",
    x"3ED39AA2",
    x"3ED3A613",
    x"3ED3B185",
    x"3ED3BCF6",
    x"3ED3C867",
    x"3ED3D3D7",
    x"3ED3DF48",
    x"3ED3EAB9",
    x"3ED3F629",
    x"3ED40199",
    x"3ED40D0A",
    x"3ED4187A",
    x"3ED423EA",
    x"3ED42F59",
    x"3ED43AC9",
    x"3ED44639",
    x"3ED451A8",
    x"3ED45D17",
    x"3ED46886",
    x"3ED473F5",
    x"3ED47F64",
    x"3ED48AD3",
    x"3ED49642",
    x"3ED4A1B0",
    x"3ED4AD1F",
    x"3ED4B88D",
    x"3ED4C3FB",
    x"3ED4CF69",
    x"3ED4DAD7",
    x"3ED4E645",
    x"3ED4F1B2",
    x"3ED4FD20",
    x"3ED5088D",
    x"3ED513FA",
    x"3ED51F68",
    x"3ED52AD5",
    x"3ED53641",
    x"3ED541AE",
    x"3ED54D1B",
    x"3ED55887",
    x"3ED563F3",
    x"3ED56F60",
    x"3ED57ACC",
    x"3ED58638",
    x"3ED591A4",
    x"3ED59D0F",
    x"3ED5A87B",
    x"3ED5B3E6",
    x"3ED5BF52",
    x"3ED5CABD",
    x"3ED5D628",
    x"3ED5E193",
    x"3ED5ECFD",
    x"3ED5F868",
    x"3ED603D3",
    x"3ED60F3D",
    x"3ED61AA7",
    x"3ED62611",
    x"3ED6317B",
    x"3ED63CE5",
    x"3ED6484F",
    x"3ED653B9",
    x"3ED65F22",
    x"3ED66A8C",
    x"3ED675F5",
    x"3ED6815E",
    x"3ED68CC7",
    x"3ED69830",
    x"3ED6A399",
    x"3ED6AF01",
    x"3ED6BA6A",
    x"3ED6C5D2",
    x"3ED6D13A",
    x"3ED6DCA2",
    x"3ED6E80A",
    x"3ED6F372",
    x"3ED6FEDA",
    x"3ED70A41",
    x"3ED715A9",
    x"3ED72110",
    x"3ED72C77",
    x"3ED737DE",
    x"3ED74345",
    x"3ED74EAC",
    x"3ED75A13",
    x"3ED76579",
    x"3ED770E0",
    x"3ED77C46",
    x"3ED787AC",
    x"3ED79312",
    x"3ED79E78",
    x"3ED7A9DE",
    x"3ED7B543",
    x"3ED7C0A9",
    x"3ED7CC0E",
    x"3ED7D773",
    x"3ED7E2D8",
    x"3ED7EE3D",
    x"3ED7F9A2",
    x"3ED80507",
    x"3ED8106B",
    x"3ED81BD0",
    x"3ED82734",
    x"3ED83298",
    x"3ED83DFC",
    x"3ED84960",
    x"3ED854C4",
    x"3ED86028",
    x"3ED86B8B",
    x"3ED876EF",
    x"3ED88252",
    x"3ED88DB5",
    x"3ED89918",
    x"3ED8A47B",
    x"3ED8AFDE",
    x"3ED8BB40",
    x"3ED8C6A3",
    x"3ED8D205",
    x"3ED8DD67",
    x"3ED8E8CA",
    x"3ED8F42C",
    x"3ED8FF8D",
    x"3ED90AEF",
    x"3ED91651",
    x"3ED921B2",
    x"3ED92D13",
    x"3ED93875",
    x"3ED943D6",
    x"3ED94F37",
    x"3ED95A97",
    x"3ED965F8",
    x"3ED97159",
    x"3ED97CB9",
    x"3ED98819",
    x"3ED99379",
    x"3ED99ED9",
    x"3ED9AA39",
    x"3ED9B599",
    x"3ED9C0F9",
    x"3ED9CC58",
    x"3ED9D7B7",
    x"3ED9E317",
    x"3ED9EE76",
    x"3ED9F9D5",
    x"3EDA0533",
    x"3EDA1092",
    x"3EDA1BF1",
    x"3EDA274F",
    x"3EDA32AD",
    x"3EDA3E0C",
    x"3EDA496A",
    x"3EDA54C8",
    x"3EDA6025",
    x"3EDA6B83",
    x"3EDA76E0",
    x"3EDA823E",
    x"3EDA8D9B",
    x"3EDA98F8",
    x"3EDAA455",
    x"3EDAAFB2",
    x"3EDABB0F",
    x"3EDAC66B",
    x"3EDAD1C8",
    x"3EDADD24",
    x"3EDAE880",
    x"3EDAF3DC",
    x"3EDAFF38",
    x"3EDB0A94",
    x"3EDB15F0",
    x"3EDB214B",
    x"3EDB2CA7",
    x"3EDB3802",
    x"3EDB435D",
    x"3EDB4EB8",
    x"3EDB5A13",
    x"3EDB656E",
    x"3EDB70C8",
    x"3EDB7C23",
    x"3EDB877D",
    x"3EDB92D7",
    x"3EDB9E31",
    x"3EDBA98B",
    x"3EDBB4E5",
    x"3EDBC03F",
    x"3EDBCB98",
    x"3EDBD6F2",
    x"3EDBE24B",
    x"3EDBEDA4",
    x"3EDBF8FD",
    x"3EDC0456",
    x"3EDC0FAF",
    x"3EDC1B08",
    x"3EDC2660",
    x"3EDC31B8",
    x"3EDC3D11",
    x"3EDC4869",
    x"3EDC53C1",
    x"3EDC5F18",
    x"3EDC6A70",
    x"3EDC75C8",
    x"3EDC811F",
    x"3EDC8C76",
    x"3EDC97CE",
    x"3EDCA325",
    x"3EDCAE7C",
    x"3EDCB9D2",
    x"3EDCC529",
    x"3EDCD07F",
    x"3EDCDBD6",
    x"3EDCE72C",
    x"3EDCF282",
    x"3EDCFDD8",
    x"3EDD092E",
    x"3EDD1484",
    x"3EDD1FD9",
    x"3EDD2B2F",
    x"3EDD3684",
    x"3EDD41D9",
    x"3EDD4D2E",
    x"3EDD5883",
    x"3EDD63D8",
    x"3EDD6F2C",
    x"3EDD7A81",
    x"3EDD85D5",
    x"3EDD912A",
    x"3EDD9C7E",
    x"3EDDA7D2",
    x"3EDDB325",
    x"3EDDBE79",
    x"3EDDC9CD",
    x"3EDDD520",
    x"3EDDE073",
    x"3EDDEBC7",
    x"3EDDF71A",
    x"3EDE026C",
    x"3EDE0DBF",
    x"3EDE1912",
    x"3EDE2464",
    x"3EDE2FB7",
    x"3EDE3B09",
    x"3EDE465B",
    x"3EDE51AD",
    x"3EDE5CFF",
    x"3EDE6851",
    x"3EDE73A2",
    x"3EDE7EF3",
    x"3EDE8A45",
    x"3EDE9596",
    x"3EDEA0E7",
    x"3EDEAC38",
    x"3EDEB789",
    x"3EDEC2D9",
    x"3EDECE2A",
    x"3EDED97A",
    x"3EDEE4CA",
    x"3EDEF01A",
    x"3EDEFB6A",
    x"3EDF06BA",
    x"3EDF120A",
    x"3EDF1D59",
    x"3EDF28A9",
    x"3EDF33F8",
    x"3EDF3F47",
    x"3EDF4A96",
    x"3EDF55E5",
    x"3EDF6134",
    x"3EDF6C82",
    x"3EDF77D1",
    x"3EDF831F",
    x"3EDF8E6D",
    x"3EDF99BB",
    x"3EDFA509",
    x"3EDFB057",
    x"3EDFBBA5",
    x"3EDFC6F2",
    x"3EDFD240",
    x"3EDFDD8D",
    x"3EDFE8DA",
    x"3EDFF427",
    x"3EDFFF74",
    x"3EE00AC1",
    x"3EE0160D",
    x"3EE0215A",
    x"3EE02CA6",
    x"3EE037F2",
    x"3EE0433E",
    x"3EE04E8A",
    x"3EE059D6",
    x"3EE06522",
    x"3EE0706D",
    x"3EE07BB8",
    x"3EE08704",
    x"3EE0924F",
    x"3EE09D9A",
    x"3EE0A8E5",
    x"3EE0B42F",
    x"3EE0BF7A",
    x"3EE0CAC4",
    x"3EE0D60E",
    x"3EE0E159",
    x"3EE0ECA3",
    x"3EE0F7ED",
    x"3EE10336",
    x"3EE10E80",
    x"3EE119C9",
    x"3EE12513",
    x"3EE1305C",
    x"3EE13BA5",
    x"3EE146EE",
    x"3EE15237",
    x"3EE15D7F",
    x"3EE168C8",
    x"3EE17410",
    x"3EE17F58",
    x"3EE18AA1",
    x"3EE195E9",
    x"3EE1A130",
    x"3EE1AC78",
    x"3EE1B7C0",
    x"3EE1C307",
    x"3EE1CE4E",
    x"3EE1D996",
    x"3EE1E4DD",
    x"3EE1F023",
    x"3EE1FB6A",
    x"3EE206B1",
    x"3EE211F7",
    x"3EE21D3E",
    x"3EE22884",
    x"3EE233CA",
    x"3EE23F10",
    x"3EE24A56",
    x"3EE2559B",
    x"3EE260E1",
    x"3EE26C26",
    x"3EE2776C",
    x"3EE282B1",
    x"3EE28DF6",
    x"3EE2993A",
    x"3EE2A47F",
    x"3EE2AFC4",
    x"3EE2BB08",
    x"3EE2C64C",
    x"3EE2D191",
    x"3EE2DCD5",
    x"3EE2E819",
    x"3EE2F35C",
    x"3EE2FEA0",
    x"3EE309E3",
    x"3EE31527",
    x"3EE3206A",
    x"3EE32BAD",
    x"3EE336F0",
    x"3EE34233",
    x"3EE34D75",
    x"3EE358B8",
    x"3EE363FA",
    x"3EE36F3D",
    x"3EE37A7F",
    x"3EE385C1",
    x"3EE39102",
    x"3EE39C44",
    x"3EE3A786",
    x"3EE3B2C7",
    x"3EE3BE08",
    x"3EE3C94A",
    x"3EE3D48B",
    x"3EE3DFCB",
    x"3EE3EB0C",
    x"3EE3F64D",
    x"3EE4018D",
    x"3EE40CCE",
    x"3EE4180E",
    x"3EE4234E",
    x"3EE42E8E",
    x"3EE439CE",
    x"3EE4450D",
    x"3EE4504D",
    x"3EE45B8C",
    x"3EE466CB",
    x"3EE4720A",
    x"3EE47D49",
    x"3EE48888",
    x"3EE493C7",
    x"3EE49F05",
    x"3EE4AA44",
    x"3EE4B582",
    x"3EE4C0C0",
    x"3EE4CBFE",
    x"3EE4D73C",
    x"3EE4E27A",
    x"3EE4EDB7",
    x"3EE4F8F5",
    x"3EE50432",
    x"3EE50F6F",
    x"3EE51AAC",
    x"3EE525E9",
    x"3EE53126",
    x"3EE53C62",
    x"3EE5479F",
    x"3EE552DB",
    x"3EE55E17",
    x"3EE56953",
    x"3EE5748F",
    x"3EE57FCB",
    x"3EE58B07",
    x"3EE59642",
    x"3EE5A17E",
    x"3EE5ACB9",
    x"3EE5B7F4",
    x"3EE5C32F",
    x"3EE5CE6A",
    x"3EE5D9A4",
    x"3EE5E4DF",
    x"3EE5F019",
    x"3EE5FB54",
    x"3EE6068E",
    x"3EE611C8",
    x"3EE61D02",
    x"3EE6283B",
    x"3EE63375",
    x"3EE63EAE",
    x"3EE649E7",
    x"3EE65521",
    x"3EE6605A",
    x"3EE66B93",
    x"3EE676CB",
    x"3EE68204",
    x"3EE68D3C",
    x"3EE69875",
    x"3EE6A3AD",
    x"3EE6AEE5",
    x"3EE6BA1D",
    x"3EE6C554",
    x"3EE6D08C",
    x"3EE6DBC4",
    x"3EE6E6FB",
    x"3EE6F232",
    x"3EE6FD69",
    x"3EE708A0",
    x"3EE713D7",
    x"3EE71F0E",
    x"3EE72A44",
    x"3EE7357A",
    x"3EE740B1",
    x"3EE74BE7",
    x"3EE7571D",
    x"3EE76253",
    x"3EE76D88",
    x"3EE778BE",
    x"3EE783F3",
    x"3EE78F28",
    x"3EE79A5D",
    x"3EE7A592",
    x"3EE7B0C7",
    x"3EE7BBFC",
    x"3EE7C731",
    x"3EE7D265",
    x"3EE7DD99",
    x"3EE7E8CD",
    x"3EE7F401",
    x"3EE7FF35",
    x"3EE80A69",
    x"3EE8159C",
    x"3EE820D0",
    x"3EE82C03",
    x"3EE83736",
    x"3EE84269",
    x"3EE84D9C",
    x"3EE858CF",
    x"3EE86402",
    x"3EE86F34",
    x"3EE87A66",
    x"3EE88599",
    x"3EE890CB",
    x"3EE89BFD",
    x"3EE8A72E",
    x"3EE8B260",
    x"3EE8BD91",
    x"3EE8C8C3",
    x"3EE8D3F4",
    x"3EE8DF25",
    x"3EE8EA56",
    x"3EE8F587",
    x"3EE900B7",
    x"3EE90BE8",
    x"3EE91718",
    x"3EE92248",
    x"3EE92D78",
    x"3EE938A8",
    x"3EE943D8",
    x"3EE94F08",
    x"3EE95A37",
    x"3EE96567",
    x"3EE97096",
    x"3EE97BC5",
    x"3EE986F4",
    x"3EE99223",
    x"3EE99D51",
    x"3EE9A880",
    x"3EE9B3AE",
    x"3EE9BEDD",
    x"3EE9CA0B",
    x"3EE9D539",
    x"3EE9E066",
    x"3EE9EB94",
    x"3EE9F6C2",
    x"3EEA01EF",
    x"3EEA0D1C",
    x"3EEA1849",
    x"3EEA2376",
    x"3EEA2EA3",
    x"3EEA39D0",
    x"3EEA44FD",
    x"3EEA5029",
    x"3EEA5B55",
    x"3EEA6681",
    x"3EEA71AD",
    x"3EEA7CD9",
    x"3EEA8805",
    x"3EEA9330",
    x"3EEA9E5C",
    x"3EEAA987",
    x"3EEAB4B2",
    x"3EEABFDD",
    x"3EEACB08",
    x"3EEAD633",
    x"3EEAE15D",
    x"3EEAEC88",
    x"3EEAF7B2",
    x"3EEB02DC",
    x"3EEB0E06",
    x"3EEB1930",
    x"3EEB245A",
    x"3EEB2F84",
    x"3EEB3AAD",
    x"3EEB45D6",
    x"3EEB50FF",
    x"3EEB5C28",
    x"3EEB6751",
    x"3EEB727A",
    x"3EEB7DA3",
    x"3EEB88CB",
    x"3EEB93F3",
    x"3EEB9F1C",
    x"3EEBAA44",
    x"3EEBB56C",
    x"3EEBC093",
    x"3EEBCBBB",
    x"3EEBD6E2",
    x"3EEBE20A",
    x"3EEBED31",
    x"3EEBF858",
    x"3EEC037F",
    x"3EEC0EA5",
    x"3EEC19CC",
    x"3EEC24F3",
    x"3EEC3019",
    x"3EEC3B3F",
    x"3EEC4665",
    x"3EEC518B",
    x"3EEC5CB1",
    x"3EEC67D6",
    x"3EEC72FC",
    x"3EEC7E21",
    x"3EEC8946",
    x"3EEC946B",
    x"3EEC9F90",
    x"3EECAAB5",
    x"3EECB5DA",
    x"3EECC0FE",
    x"3EECCC22",
    x"3EECD747",
    x"3EECE26B",
    x"3EECED8F",
    x"3EECF8B2",
    x"3EED03D6",
    x"3EED0EF9",
    x"3EED1A1D",
    x"3EED2540",
    x"3EED3063",
    x"3EED3B86",
    x"3EED46A9",
    x"3EED51CB",
    x"3EED5CEE",
    x"3EED6810",
    x"3EED7332",
    x"3EED7E54",
    x"3EED8976",
    x"3EED9498",
    x"3EED9FB9",
    x"3EEDAADB",
    x"3EEDB5FC",
    x"3EEDC11D",
    x"3EEDCC3E",
    x"3EEDD75F",
    x"3EEDE280",
    x"3EEDEDA1",
    x"3EEDF8C1",
    x"3EEE03E2",
    x"3EEE0F02",
    x"3EEE1A22",
    x"3EEE2542",
    x"3EEE3061",
    x"3EEE3B81",
    x"3EEE46A0",
    x"3EEE51C0",
    x"3EEE5CDF",
    x"3EEE67FE",
    x"3EEE731D",
    x"3EEE7E3C",
    x"3EEE895A",
    x"3EEE9479",
    x"3EEE9F97",
    x"3EEEAAB5",
    x"3EEEB5D3",
    x"3EEEC0F1",
    x"3EEECC0F",
    x"3EEED72C",
    x"3EEEE24A",
    x"3EEEED67",
    x"3EEEF884",
    x"3EEF03A1",
    x"3EEF0EBE",
    x"3EEF19DB",
    x"3EEF24F7",
    x"3EEF3014",
    x"3EEF3B30",
    x"3EEF464C",
    x"3EEF5168",
    x"3EEF5C84",
    x"3EEF67A0",
    x"3EEF72BC",
    x"3EEF7DD7",
    x"3EEF88F2",
    x"3EEF940D",
    x"3EEF9F28",
    x"3EEFAA43",
    x"3EEFB55E",
    x"3EEFC079",
    x"3EEFCB93",
    x"3EEFD6AD",
    x"3EEFE1C7",
    x"3EEFECE1",
    x"3EEFF7FB",
    x"3EF00315",
    x"3EF00E2E",
    x"3EF01948",
    x"3EF02461",
    x"3EF02F7A",
    x"3EF03A93",
    x"3EF045AC",
    x"3EF050C5",
    x"3EF05BDD",
    x"3EF066F6",
    x"3EF0720E",
    x"3EF07D26",
    x"3EF0883E",
    x"3EF09356",
    x"3EF09E6E",
    x"3EF0A985",
    x"3EF0B49C",
    x"3EF0BFB4",
    x"3EF0CACB",
    x"3EF0D5E2",
    x"3EF0E0F9",
    x"3EF0EC0F",
    x"3EF0F726",
    x"3EF1023C",
    x"3EF10D52",
    x"3EF11868",
    x"3EF1237E",
    x"3EF12E94",
    x"3EF139AA",
    x"3EF144BF",
    x"3EF14FD5",
    x"3EF15AEA",
    x"3EF165FF",
    x"3EF17114",
    x"3EF17C28",
    x"3EF1873D",
    x"3EF19252",
    x"3EF19D66",
    x"3EF1A87A",
    x"3EF1B38E",
    x"3EF1BEA2",
    x"3EF1C9B6",
    x"3EF1D4C9",
    x"3EF1DFDD",
    x"3EF1EAF0",
    x"3EF1F603",
    x"3EF20116",
    x"3EF20C29",
    x"3EF2173C",
    x"3EF2224F",
    x"3EF22D61",
    x"3EF23873",
    x"3EF24385",
    x"3EF24E97",
    x"3EF259A9",
    x"3EF264BB",
    x"3EF26FCD",
    x"3EF27ADE",
    x"3EF285EF",
    x"3EF29100",
    x"3EF29C11",
    x"3EF2A722",
    x"3EF2B233",
    x"3EF2BD43",
    x"3EF2C854",
    x"3EF2D364",
    x"3EF2DE74",
    x"3EF2E984",
    x"3EF2F494",
    x"3EF2FFA4",
    x"3EF30AB3",
    x"3EF315C2",
    x"3EF320D2",
    x"3EF32BE1",
    x"3EF336F0",
    x"3EF341FE",
    x"3EF34D0D",
    x"3EF3581C",
    x"3EF3632A",
    x"3EF36E38",
    x"3EF37946",
    x"3EF38454",
    x"3EF38F62",
    x"3EF39A6F",
    x"3EF3A57D",
    x"3EF3B08A",
    x"3EF3BB97",
    x"3EF3C6A4",
    x"3EF3D1B1",
    x"3EF3DCBE",
    x"3EF3E7CB",
    x"3EF3F2D7",
    x"3EF3FDE3",
    x"3EF408F0",
    x"3EF413FB",
    x"3EF41F07",
    x"3EF42A13",
    x"3EF4351F",
    x"3EF4402A",
    x"3EF44B35",
    x"3EF45640",
    x"3EF4614B",
    x"3EF46C56",
    x"3EF47761",
    x"3EF4826B",
    x"3EF48D76",
    x"3EF49880",
    x"3EF4A38A",
    x"3EF4AE94",
    x"3EF4B99E",
    x"3EF4C4A7",
    x"3EF4CFB1",
    x"3EF4DABA",
    x"3EF4E5C3",
    x"3EF4F0CC",
    x"3EF4FBD5",
    x"3EF506DE",
    x"3EF511E7",
    x"3EF51CEF",
    x"3EF527F8",
    x"3EF53300",
    x"3EF53E08",
    x"3EF54910",
    x"3EF55417",
    x"3EF55F1F",
    x"3EF56A26",
    x"3EF5752E",
    x"3EF58035",
    x"3EF58B3C",
    x"3EF59643",
    x"3EF5A149",
    x"3EF5AC50",
    x"3EF5B756",
    x"3EF5C25C",
    x"3EF5CD62",
    x"3EF5D868",
    x"3EF5E36E",
    x"3EF5EE74",
    x"3EF5F979",
    x"3EF6047F",
    x"3EF60F84",
    x"3EF61A89",
    x"3EF6258E",
    x"3EF63093",
    x"3EF63B97",
    x"3EF6469C",
    x"3EF651A0",
    x"3EF65CA4",
    x"3EF667A8",
    x"3EF672AC",
    x"3EF67DB0",
    x"3EF688B3",
    x"3EF693B7",
    x"3EF69EBA",
    x"3EF6A9BD",
    x"3EF6B4C0",
    x"3EF6BFC3",
    x"3EF6CAC6",
    x"3EF6D5C8",
    x"3EF6E0CB",
    x"3EF6EBCD",
    x"3EF6F6CF",
    x"3EF701D1",
    x"3EF70CD3",
    x"3EF717D4",
    x"3EF722D6",
    x"3EF72DD7",
    x"3EF738D8",
    x"3EF743D9",
    x"3EF74EDA",
    x"3EF759DB",
    x"3EF764DC",
    x"3EF76FDC",
    x"3EF77ADC",
    x"3EF785DC",
    x"3EF790DC",
    x"3EF79BDC",
    x"3EF7A6DC",
    x"3EF7B1DC",
    x"3EF7BCDB",
    x"3EF7C7DA",
    x"3EF7D2D9",
    x"3EF7DDD8",
    x"3EF7E8D7",
    x"3EF7F3D6",
    x"3EF7FED4",
    x"3EF809D3",
    x"3EF814D1",
    x"3EF81FCF",
    x"3EF82ACD",
    x"3EF835CB",
    x"3EF840C8",
    x"3EF84BC6",
    x"3EF856C3",
    x"3EF861C0",
    x"3EF86CBD",
    x"3EF877BA",
    x"3EF882B7",
    x"3EF88DB3",
    x"3EF898B0",
    x"3EF8A3AC",
    x"3EF8AEA8",
    x"3EF8B9A4",
    x"3EF8C4A0",
    x"3EF8CF9C",
    x"3EF8DA97",
    x"3EF8E592",
    x"3EF8F08E",
    x"3EF8FB89",
    x"3EF90684",
    x"3EF9117E",
    x"3EF91C79",
    x"3EF92773",
    x"3EF9326E",
    x"3EF93D68",
    x"3EF94862",
    x"3EF9535C",
    x"3EF95E56",
    x"3EF9694F",
    x"3EF97449",
    x"3EF97F42",
    x"3EF98A3B",
    x"3EF99534",
    x"3EF9A02D",
    x"3EF9AB25",
    x"3EF9B61E",
    x"3EF9C116",
    x"3EF9CC0E",
    x"3EF9D707",
    x"3EF9E1FE",
    x"3EF9ECF6",
    x"3EF9F7EE",
    x"3EFA02E5",
    x"3EFA0DDD",
    x"3EFA18D4",
    x"3EFA23CB",
    x"3EFA2EC2",
    x"3EFA39B8",
    x"3EFA44AF",
    x"3EFA4FA5",
    x"3EFA5A9C",
    x"3EFA6592",
    x"3EFA7088",
    x"3EFA7B7D",
    x"3EFA8673",
    x"3EFA9169",
    x"3EFA9C5E",
    x"3EFAA753",
    x"3EFAB248",
    x"3EFABD3D",
    x"3EFAC832",
    x"3EFAD326",
    x"3EFADE1B",
    x"3EFAE90F",
    x"3EFAF403",
    x"3EFAFEF7",
    x"3EFB09EB",
    x"3EFB14DF",
    x"3EFB1FD2",
    x"3EFB2AC6",
    x"3EFB35B9",
    x"3EFB40AC",
    x"3EFB4B9F",
    x"3EFB5692",
    x"3EFB6184",
    x"3EFB6C77",
    x"3EFB7769",
    x"3EFB825B",
    x"3EFB8D4D",
    x"3EFB983F",
    x"3EFBA331",
    x"3EFBAE22",
    x"3EFBB914",
    x"3EFBC405",
    x"3EFBCEF6",
    x"3EFBD9E7",
    x"3EFBE4D8",
    x"3EFBEFC9",
    x"3EFBFAB9",
    x"3EFC05AA",
    x"3EFC109A",
    x"3EFC1B8A",
    x"3EFC267A",
    x"3EFC3169",
    x"3EFC3C59",
    x"3EFC4748",
    x"3EFC5238",
    x"3EFC5D27",
    x"3EFC6816",
    x"3EFC7305",
    x"3EFC7DF3",
    x"3EFC88E2",
    x"3EFC93D0",
    x"3EFC9EBF",
    x"3EFCA9AD",
    x"3EFCB49B",
    x"3EFCBF88",
    x"3EFCCA76",
    x"3EFCD563",
    x"3EFCE051",
    x"3EFCEB3E",
    x"3EFCF62B",
    x"3EFD0118",
    x"3EFD0C04",
    x"3EFD16F1",
    x"3EFD21DD",
    x"3EFD2CCA",
    x"3EFD37B6",
    x"3EFD42A2",
    x"3EFD4D8D",
    x"3EFD5879",
    x"3EFD6365",
    x"3EFD6E50",
    x"3EFD793B",
    x"3EFD8426",
    x"3EFD8F11",
    x"3EFD99FC",
    x"3EFDA4E6",
    x"3EFDAFD1",
    x"3EFDBABB",
    x"3EFDC5A5",
    x"3EFDD08F",
    x"3EFDDB79",
    x"3EFDE662",
    x"3EFDF14C",
    x"3EFDFC35",
    x"3EFE071E",
    x"3EFE1207",
    x"3EFE1CF0",
    x"3EFE27D9",
    x"3EFE32C2",
    x"3EFE3DAA",
    x"3EFE4892",
    x"3EFE537A",
    x"3EFE5E62",
    x"3EFE694A",
    x"3EFE7432",
    x"3EFE7F19",
    x"3EFE8A01",
    x"3EFE94E8",
    x"3EFE9FCF",
    x"3EFEAAB6",
    x"3EFEB59D",
    x"3EFEC083",
    x"3EFECB6A",
    x"3EFED650",
    x"3EFEE136",
    x"3EFEEC1C",
    x"3EFEF702",
    x"3EFF01E8",
    x"3EFF0CCD",
    x"3EFF17B2",
    x"3EFF2298",
    x"3EFF2D7D",
    x"3EFF3862",
    x"3EFF4346",
    x"3EFF4E2B",
    x"3EFF590F",
    x"3EFF63F4",
    x"3EFF6ED8",
    x"3EFF79BC",
    x"3EFF849F",
    x"3EFF8F83",
    x"3EFF9A67",
    x"3EFFA54A",
    x"3EFFB02D",
    x"3EFFBB10",
    x"3EFFC5F3",
    x"3EFFD0D6",
    x"3EFFDBB8",
    x"3EFFE69B",
    x"3EFFF17D",
    x"3EFFFC5F",
    x"3F0003A1",
    x"3F000912",
    x"3F000E82",
    x"3F0013F3",
    x"3F001964",
    x"3F001ED4",
    x"3F002445",
    x"3F0029B5",
    x"3F002F26",
    x"3F003496",
    x"3F003A06",
    x"3F003F76",
    x"3F0044E6",
    x"3F004A56",
    x"3F004FC6",
    x"3F005536",
    x"3F005AA6",
    x"3F006016",
    x"3F006585",
    x"3F006AF5",
    x"3F007064",
    x"3F0075D4",
    x"3F007B43",
    x"3F0080B2",
    x"3F008621",
    x"3F008B90",
    x"3F0090FF",
    x"3F00966E",
    x"3F009BDD",
    x"3F00A14C",
    x"3F00A6BA",
    x"3F00AC29",
    x"3F00B197",
    x"3F00B706",
    x"3F00BC74",
    x"3F00C1E2",
    x"3F00C751",
    x"3F00CCBF",
    x"3F00D22D",
    x"3F00D79B",
    x"3F00DD09",
    x"3F00E276",
    x"3F00E7E4",
    x"3F00ED52",
    x"3F00F2BF",
    x"3F00F82D",
    x"3F00FD9A",
    x"3F010308",
    x"3F010875",
    x"3F010DE2",
    x"3F01134F",
    x"3F0118BC",
    x"3F011E29",
    x"3F012396",
    x"3F012903",
    x"3F012E70",
    x"3F0133DC",
    x"3F013949",
    x"3F013EB5",
    x"3F014422",
    x"3F01498E",
    x"3F014EFA",
    x"3F015467",
    x"3F0159D3",
    x"3F015F3F",
    x"3F0164AB",
    x"3F016A17",
    x"3F016F82",
    x"3F0174EE",
    x"3F017A5A",
    x"3F017FC5",
    x"3F018531",
    x"3F018A9C",
    x"3F019007",
    x"3F019573",
    x"3F019ADE",
    x"3F01A049",
    x"3F01A5B4",
    x"3F01AB1F",
    x"3F01B08A",
    x"3F01B5F5",
    x"3F01BB5F",
    x"3F01C0CA",
    x"3F01C634",
    x"3F01CB9F",
    x"3F01D109",
    x"3F01D674",
    x"3F01DBDE",
    x"3F01E148",
    x"3F01E6B2",
    x"3F01EC1C",
    x"3F01F186",
    x"3F01F6F0",
    x"3F01FC59",
    x"3F0201C3",
    x"3F02072D",
    x"3F020C96",
    x"3F021200",
    x"3F021769",
    x"3F021CD2",
    x"3F02223C",
    x"3F0227A5",
    x"3F022D0E",
    x"3F023277",
    x"3F0237E0",
    x"3F023D48",
    x"3F0242B1",
    x"3F02481A",
    x"3F024D82",
    x"3F0252EB",
    x"3F025853",
    x"3F025DBC",
    x"3F026324",
    x"3F02688C",
    x"3F026DF4",
    x"3F02735C",
    x"3F0278C4",
    x"3F027E2C",
    x"3F028394",
    x"3F0288FC",
    x"3F028E63",
    x"3F0293CB",
    x"3F029932",
    x"3F029E9A",
    x"3F02A401",
    x"3F02A968",
    x"3F02AED0",
    x"3F02B437",
    x"3F02B99E",
    x"3F02BF05",
    x"3F02C46B",
    x"3F02C9D2",
    x"3F02CF39",
    x"3F02D49F",
    x"3F02DA06",
    x"3F02DF6C",
    x"3F02E4D3",
    x"3F02EA39",
    x"3F02EF9F",
    x"3F02F506",
    x"3F02FA6C",
    x"3F02FFD2",
    x"3F030537",
    x"3F030A9D",
    x"3F031003",
    x"3F031569",
    x"3F031ACE",
    x"3F032034",
    x"3F032599",
    x"3F032AFF",
    x"3F033064",
    x"3F0335C9",
    x"3F033B2E",
    x"3F034093",
    x"3F0345F8",
    x"3F034B5D",
    x"3F0350C2",
    x"3F035627",
    x"3F035B8B",
    x"3F0360F0",
    x"3F036654",
    x"3F036BB9",
    x"3F03711D",
    x"3F037681",
    x"3F037BE5",
    x"3F03814A",
    x"3F0386AE",
    x"3F038C11",
    x"3F039175",
    x"3F0396D9",
    x"3F039C3D",
    x"3F03A1A0",
    x"3F03A704",
    x"3F03AC67",
    x"3F03B1CB",
    x"3F03B72E",
    x"3F03BC91",
    x"3F03C1F4",
    x"3F03C757",
    x"3F03CCBA",
    x"3F03D21D",
    x"3F03D780",
    x"3F03DCE3",
    x"3F03E246",
    x"3F03E7A8",
    x"3F03ED0B",
    x"3F03F26D",
    x"3F03F7CF",
    x"3F03FD32",
    x"3F040294",
    x"3F0407F6",
    x"3F040D58",
    x"3F0412BA",
    x"3F04181C",
    x"3F041D7E",
    x"3F0422DF",
    x"3F042841",
    x"3F042DA2",
    x"3F043304",
    x"3F043865",
    x"3F043DC7",
    x"3F044328",
    x"3F044889",
    x"3F044DEA",
    x"3F04534B",
    x"3F0458AC",
    x"3F045E0D",
    x"3F04636E",
    x"3F0468CE",
    x"3F046E2F",
    x"3F04738F",
    x"3F0478F0",
    x"3F047E50",
    x"3F0483B0",
    x"3F048911",
    x"3F048E71",
    x"3F0493D1",
    x"3F049931",
    x"3F049E91",
    x"3F04A3F0",
    x"3F04A950",
    x"3F04AEB0",
    x"3F04B40F",
    x"3F04B96F",
    x"3F04BECE",
    x"3F04C42D",
    x"3F04C98D",
    x"3F04CEEC",
    x"3F04D44B",
    x"3F04D9AA",
    x"3F04DF09",
    x"3F04E468",
    x"3F04E9C6",
    x"3F04EF25",
    x"3F04F484",
    x"3F04F9E2",
    x"3F04FF41",
    x"3F05049F",
    x"3F0509FD",
    x"3F050F5B",
    x"3F0514BA",
    x"3F051A18",
    x"3F051F75",
    x"3F0524D3",
    x"3F052A31",
    x"3F052F8F",
    x"3F0534EC",
    x"3F053A4A",
    x"3F053FA8",
    x"3F054505",
    x"3F054A62",
    x"3F054FBF",
    x"3F05551D",
    x"3F055A7A",
    x"3F055FD7",
    x"3F056534",
    x"3F056A90",
    x"3F056FED",
    x"3F05754A",
    x"3F057AA6",
    x"3F058003",
    x"3F05855F",
    x"3F058ABC",
    x"3F059018",
    x"3F059574",
    x"3F059AD0",
    x"3F05A02C",
    x"3F05A588",
    x"3F05AAE4",
    x"3F05B040",
    x"3F05B59C",
    x"3F05BAF7",
    x"3F05C053",
    x"3F05C5AE",
    x"3F05CB0A",
    x"3F05D065",
    x"3F05D5C0",
    x"3F05DB1B",
    x"3F05E076",
    x"3F05E5D1",
    x"3F05EB2C",
    x"3F05F087",
    x"3F05F5E2",
    x"3F05FB3C",
    x"3F060097",
    x"3F0605F1",
    x"3F060B4C",
    x"3F0610A6",
    x"3F061600",
    x"3F061B5B",
    x"3F0620B5",
    x"3F06260F",
    x"3F062B69",
    x"3F0630C2",
    x"3F06361C",
    x"3F063B76",
    x"3F0640CF",
    x"3F064629",
    x"3F064B82",
    x"3F0650DC",
    x"3F065635",
    x"3F065B8E",
    x"3F0660E7",
    x"3F066640",
    x"3F066B99",
    x"3F0670F2",
    x"3F06764B",
    x"3F067BA4",
    x"3F0680FC",
    x"3F068655",
    x"3F068BAD",
    x"3F069106",
    x"3F06965E",
    x"3F069BB6",
    x"3F06A10E",
    x"3F06A667",
    x"3F06ABBF",
    x"3F06B116",
    x"3F06B66E",
    x"3F06BBC6",
    x"3F06C11E",
    x"3F06C675",
    x"3F06CBCD",
    x"3F06D124",
    x"3F06D67B",
    x"3F06DBD3",
    x"3F06E12A",
    x"3F06E681",
    x"3F06EBD8",
    x"3F06F12F",
    x"3F06F686",
    x"3F06FBDD",
    x"3F070133",
    x"3F07068A",
    x"3F070BE0",
    x"3F071137",
    x"3F07168D",
    x"3F071BE3",
    x"3F07213A",
    x"3F072690",
    x"3F072BE6",
    x"3F07313C",
    x"3F073692",
    x"3F073BE7",
    x"3F07413D",
    x"3F074693",
    x"3F074BE8",
    x"3F07513E",
    x"3F075693",
    x"3F075BE8",
    x"3F07613E",
    x"3F076693",
    x"3F076BE8",
    x"3F07713D",
    x"3F077692",
    x"3F077BE6",
    x"3F07813B",
    x"3F078690",
    x"3F078BE4",
    x"3F079139",
    x"3F07968D",
    x"3F079BE2",
    x"3F07A136",
    x"3F07A68A",
    x"3F07ABDE",
    x"3F07B132",
    x"3F07B686",
    x"3F07BBDA",
    x"3F07C12E",
    x"3F07C681",
    x"3F07CBD5",
    x"3F07D128",
    x"3F07D67C",
    x"3F07DBCF",
    x"3F07E122",
    x"3F07E676",
    x"3F07EBC9",
    x"3F07F11C",
    x"3F07F66F",
    x"3F07FBC1",
    x"3F080114",
    x"3F080667",
    x"3F080BB9",
    x"3F08110C",
    x"3F08165E",
    x"3F081BB1",
    x"3F082103",
    x"3F082655",
    x"3F082BA7",
    x"3F0830F9",
    x"3F08364B",
    x"3F083B9D",
    x"3F0840EF",
    x"3F084641",
    x"3F084B92",
    x"3F0850E4",
    x"3F085635",
    x"3F085B87",
    x"3F0860D8",
    x"3F086629",
    x"3F086B7A",
    x"3F0870CB",
    x"3F08761C",
    x"3F087B6D",
    x"3F0880BE",
    x"3F08860F",
    x"3F088B5F",
    x"3F0890B0",
    x"3F089600",
    x"3F089B51",
    x"3F08A0A1",
    x"3F08A5F1",
    x"3F08AB41",
    x"3F08B091",
    x"3F08B5E1",
    x"3F08BB31",
    x"3F08C081",
    x"3F08C5D1",
    x"3F08CB20",
    x"3F08D070",
    x"3F08D5BF",
    x"3F08DB0F",
    x"3F08E05E",
    x"3F08E5AD",
    x"3F08EAFD",
    x"3F08F04C",
    x"3F08F59B",
    x"3F08FAEA",
    x"3F090038",
    x"3F090587",
    x"3F090AD6",
    x"3F091024",
    x"3F091573",
    x"3F091AC1",
    x"3F092010",
    x"3F09255E",
    x"3F092AAC",
    x"3F092FFA",
    x"3F093548",
    x"3F093A96",
    x"3F093FE4",
    x"3F094531",
    x"3F094A7F",
    x"3F094FCD",
    x"3F09551A",
    x"3F095A68",
    x"3F095FB5",
    x"3F096502",
    x"3F096A4F",
    x"3F096F9C",
    x"3F0974E9",
    x"3F097A36",
    x"3F097F83",
    x"3F0984D0",
    x"3F098A1D",
    x"3F098F69",
    x"3F0994B6",
    x"3F099A02",
    x"3F099F4E",
    x"3F09A49B",
    x"3F09A9E7",
    x"3F09AF33",
    x"3F09B47F",
    x"3F09B9CB",
    x"3F09BF17",
    x"3F09C463",
    x"3F09C9AE",
    x"3F09CEFA",
    x"3F09D445",
    x"3F09D991",
    x"3F09DEDC",
    x"3F09E427",
    x"3F09E973",
    x"3F09EEBE",
    x"3F09F409",
    x"3F09F954",
    x"3F09FE9E",
    x"3F0A03E9",
    x"3F0A0934",
    x"3F0A0E7E",
    x"3F0A13C9",
    x"3F0A1913",
    x"3F0A1E5E",
    x"3F0A23A8",
    x"3F0A28F2",
    x"3F0A2E3C",
    x"3F0A3386",
    x"3F0A38D0",
    x"3F0A3E1A",
    x"3F0A4364",
    x"3F0A48AD",
    x"3F0A4DF7",
    x"3F0A5341",
    x"3F0A588A",
    x"3F0A5DD3",
    x"3F0A631D",
    x"3F0A6866",
    x"3F0A6DAF",
    x"3F0A72F8",
    x"3F0A7841",
    x"3F0A7D8A",
    x"3F0A82D2",
    x"3F0A881B",
    x"3F0A8D64",
    x"3F0A92AC",
    x"3F0A97F5",
    x"3F0A9D3D",
    x"3F0AA285",
    x"3F0AA7CD",
    x"3F0AAD16",
    x"3F0AB25E",
    x"3F0AB7A5",
    x"3F0ABCED",
    x"3F0AC235",
    x"3F0AC77D",
    x"3F0ACCC4",
    x"3F0AD20C",
    x"3F0AD753",
    x"3F0ADC9B",
    x"3F0AE1E2",
    x"3F0AE729",
    x"3F0AEC70",
    x"3F0AF1B7",
    x"3F0AF6FE",
    x"3F0AFC45",
    x"3F0B018C",
    x"3F0B06D2",
    x"3F0B0C19",
    x"3F0B115F",
    x"3F0B16A6",
    x"3F0B1BEC",
    x"3F0B2132",
    x"3F0B2679",
    x"3F0B2BBF",
    x"3F0B3105",
    x"3F0B364B",
    x"3F0B3B90",
    x"3F0B40D6",
    x"3F0B461C",
    x"3F0B4B61",
    x"3F0B50A7",
    x"3F0B55EC",
    x"3F0B5B32",
    x"3F0B6077",
    x"3F0B65BC",
    x"3F0B6B01",
    x"3F0B7046",
    x"3F0B758B",
    x"3F0B7AD0",
    x"3F0B8015",
    x"3F0B8559",
    x"3F0B8A9E",
    x"3F0B8FE2",
    x"3F0B9527",
    x"3F0B9A6B",
    x"3F0B9FAF",
    x"3F0BA4F4",
    x"3F0BAA38",
    x"3F0BAF7C",
    x"3F0BB4BF",
    x"3F0BBA03",
    x"3F0BBF47",
    x"3F0BC48B",
    x"3F0BC9CE",
    x"3F0BCF12",
    x"3F0BD455",
    x"3F0BD998",
    x"3F0BDEDC",
    x"3F0BE41F",
    x"3F0BE962",
    x"3F0BEEA5",
    x"3F0BF3E8",
    x"3F0BF92B",
    x"3F0BFE6D",
    x"3F0C03B0",
    x"3F0C08F2",
    x"3F0C0E35",
    x"3F0C1377",
    x"3F0C18BA",
    x"3F0C1DFC",
    x"3F0C233E",
    x"3F0C2880",
    x"3F0C2DC2",
    x"3F0C3304",
    x"3F0C3846",
    x"3F0C3D87",
    x"3F0C42C9",
    x"3F0C480B",
    x"3F0C4D4C",
    x"3F0C528D",
    x"3F0C57CF",
    x"3F0C5D10",
    x"3F0C6251",
    x"3F0C6792",
    x"3F0C6CD3",
    x"3F0C7214",
    x"3F0C7755",
    x"3F0C7C95",
    x"3F0C81D6",
    x"3F0C8716",
    x"3F0C8C57",
    x"3F0C9197",
    x"3F0C96D7",
    x"3F0C9C18",
    x"3F0CA158",
    x"3F0CA698",
    x"3F0CABD8",
    x"3F0CB118",
    x"3F0CB657",
    x"3F0CBB97",
    x"3F0CC0D7",
    x"3F0CC616",
    x"3F0CCB56",
    x"3F0CD095",
    x"3F0CD5D4",
    x"3F0CDB13",
    x"3F0CE052",
    x"3F0CE591",
    x"3F0CEAD0",
    x"3F0CF00F",
    x"3F0CF54E",
    x"3F0CFA8D",
    x"3F0CFFCB",
    x"3F0D050A",
    x"3F0D0A48",
    x"3F0D0F86",
    x"3F0D14C5",
    x"3F0D1A03",
    x"3F0D1F41",
    x"3F0D247F",
    x"3F0D29BD",
    x"3F0D2EFA",
    x"3F0D3438",
    x"3F0D3976",
    x"3F0D3EB3",
    x"3F0D43F1",
    x"3F0D492E",
    x"3F0D4E6C",
    x"3F0D53A9",
    x"3F0D58E6",
    x"3F0D5E23",
    x"3F0D6360",
    x"3F0D689D",
    x"3F0D6DDA",
    x"3F0D7316",
    x"3F0D7853",
    x"3F0D7D8F",
    x"3F0D82CC",
    x"3F0D8808",
    x"3F0D8D45",
    x"3F0D9281",
    x"3F0D97BD",
    x"3F0D9CF9",
    x"3F0DA235",
    x"3F0DA771",
    x"3F0DACAC",
    x"3F0DB1E8",
    x"3F0DB724",
    x"3F0DBC5F",
    x"3F0DC19B",
    x"3F0DC6D6",
    x"3F0DCC11",
    x"3F0DD14C",
    x"3F0DD687",
    x"3F0DDBC2",
    x"3F0DE0FD",
    x"3F0DE638",
    x"3F0DEB73",
    x"3F0DF0AE",
    x"3F0DF5E8",
    x"3F0DFB23",
    x"3F0E005D",
    x"3F0E0597",
    x"3F0E0AD2",
    x"3F0E100C",
    x"3F0E1546",
    x"3F0E1A80",
    x"3F0E1FBA",
    x"3F0E24F3",
    x"3F0E2A2D",
    x"3F0E2F67",
    x"3F0E34A0",
    x"3F0E39DA",
    x"3F0E3F13",
    x"3F0E444C",
    x"3F0E4986",
    x"3F0E4EBF",
    x"3F0E53F8",
    x"3F0E5931",
    x"3F0E5E6A",
    x"3F0E63A2",
    x"3F0E68DB",
    x"3F0E6E14",
    x"3F0E734C",
    x"3F0E7885",
    x"3F0E7DBD",
    x"3F0E82F5",
    x"3F0E882D",
    x"3F0E8D65",
    x"3F0E929D",
    x"3F0E97D5",
    x"3F0E9D0D",
    x"3F0EA245",
    x"3F0EA77D",
    x"3F0EACB4",
    x"3F0EB1EC",
    x"3F0EB723",
    x"3F0EBC5A",
    x"3F0EC192",
    x"3F0EC6C9",
    x"3F0ECC00",
    x"3F0ED137",
    x"3F0ED66E",
    x"3F0EDBA4",
    x"3F0EE0DB",
    x"3F0EE612",
    x"3F0EEB48",
    x"3F0EF07F",
    x"3F0EF5B5",
    x"3F0EFAEB",
    x"3F0F0022",
    x"3F0F0558",
    x"3F0F0A8E",
    x"3F0F0FC4",
    x"3F0F14FA",
    x"3F0F1A2F",
    x"3F0F1F65",
    x"3F0F249B",
    x"3F0F29D0",
    x"3F0F2F05",
    x"3F0F343B",
    x"3F0F3970",
    x"3F0F3EA5",
    x"3F0F43DA",
    x"3F0F490F",
    x"3F0F4E44",
    x"3F0F5379",
    x"3F0F58AE",
    x"3F0F5DE2",
    x"3F0F6317",
    x"3F0F684B",
    x"3F0F6D80",
    x"3F0F72B4",
    x"3F0F77E8",
    x"3F0F7D1C",
    x"3F0F8250",
    x"3F0F8784",
    x"3F0F8CB8",
    x"3F0F91EC",
    x"3F0F9720",
    x"3F0F9C53",
    x"3F0FA187",
    x"3F0FA6BA",
    x"3F0FABEE",
    x"3F0FB121",
    x"3F0FB654",
    x"3F0FBB87",
    x"3F0FC0BA",
    x"3F0FC5ED",
    x"3F0FCB20",
    x"3F0FD053",
    x"3F0FD585",
    x"3F0FDAB8",
    x"3F0FDFEA",
    x"3F0FE51D",
    x"3F0FEA4F",
    x"3F0FEF81",
    x"3F0FF4B3",
    x"3F0FF9E5",
    x"3F0FFF17",
    x"3F100449",
    x"3F10097B",
    x"3F100EAD",
    x"3F1013DE",
    x"3F101910",
    x"3F101E41",
    x"3F102373",
    x"3F1028A4",
    x"3F102DD5",
    x"3F103306",
    x"3F103837",
    x"3F103D68",
    x"3F104299",
    x"3F1047CA",
    x"3F104CFA",
    x"3F10522B",
    x"3F10575B",
    x"3F105C8C",
    x"3F1061BC",
    x"3F1066EC",
    x"3F106C1C",
    x"3F10714C",
    x"3F10767C",
    x"3F107BAC",
    x"3F1080DC",
    x"3F10860C",
    x"3F108B3B",
    x"3F10906B",
    x"3F10959A",
    x"3F109ACA",
    x"3F109FF9",
    x"3F10A528",
    x"3F10AA57",
    x"3F10AF86",
    x"3F10B4B5",
    x"3F10B9E4",
    x"3F10BF13",
    x"3F10C441",
    x"3F10C970",
    x"3F10CE9E",
    x"3F10D3CD",
    x"3F10D8FB",
    x"3F10DE29",
    x"3F10E357",
    x"3F10E885",
    x"3F10EDB3",
    x"3F10F2E1",
    x"3F10F80F",
    x"3F10FD3D",
    x"3F11026A",
    x"3F110798",
    x"3F110CC5",
    x"3F1111F3",
    x"3F111720",
    x"3F111C4D",
    x"3F11217A",
    x"3F1126A7",
    x"3F112BD4",
    x"3F113101",
    x"3F11362E",
    x"3F113B5A",
    x"3F114087",
    x"3F1145B3",
    x"3F114AE0",
    x"3F11500C",
    x"3F115538",
    x"3F115A64",
    x"3F115F90",
    x"3F1164BC",
    x"3F1169E8",
    x"3F116F14",
    x"3F117440",
    x"3F11796B",
    x"3F117E97",
    x"3F1183C2",
    x"3F1188ED",
    x"3F118E19",
    x"3F119344",
    x"3F11986F",
    x"3F119D9A",
    x"3F11A2C5",
    x"3F11A7F0",
    x"3F11AD1A",
    x"3F11B245",
    x"3F11B76F",
    x"3F11BC9A",
    x"3F11C1C4",
    x"3F11C6EF",
    x"3F11CC19",
    x"3F11D143",
    x"3F11D66D",
    x"3F11DB97",
    x"3F11E0C1",
    x"3F11E5EA",
    x"3F11EB14",
    x"3F11F03E",
    x"3F11F567",
    x"3F11FA91",
    x"3F11FFBA",
    x"3F1204E3",
    x"3F120A0C",
    x"3F120F35",
    x"3F12145E",
    x"3F121987",
    x"3F121EB0",
    x"3F1223D9",
    x"3F122901",
    x"3F122E2A",
    x"3F123352",
    x"3F12387A",
    x"3F123DA3",
    x"3F1242CB",
    x"3F1247F3",
    x"3F124D1B",
    x"3F125243",
    x"3F12576B",
    x"3F125C92",
    x"3F1261BA",
    x"3F1266E2",
    x"3F126C09",
    x"3F127130",
    x"3F127658",
    x"3F127B7F",
    x"3F1280A6",
    x"3F1285CD",
    x"3F128AF4",
    x"3F12901B",
    x"3F129542",
    x"3F129A68",
    x"3F129F8F",
    x"3F12A4B5",
    x"3F12A9DC",
    x"3F12AF02",
    x"3F12B428",
    x"3F12B94E",
    x"3F12BE74",
    x"3F12C39A",
    x"3F12C8C0",
    x"3F12CDE6",
    x"3F12D30C",
    x"3F12D831",
    x"3F12DD57",
    x"3F12E27C",
    x"3F12E7A2",
    x"3F12ECC7",
    x"3F12F1EC",
    x"3F12F711",
    x"3F12FC36",
    x"3F13015B",
    x"3F130680",
    x"3F130BA5",
    x"3F1310C9",
    x"3F1315EE",
    x"3F131B12",
    x"3F132037",
    x"3F13255B",
    x"3F132A7F",
    x"3F132FA3",
    x"3F1334C7",
    x"3F1339EB",
    x"3F133F0F",
    x"3F134433",
    x"3F134956",
    x"3F134E7A",
    x"3F13539D",
    x"3F1358C1",
    x"3F135DE4",
    x"3F136307",
    x"3F13682A",
    x"3F136D4D",
    x"3F137270",
    x"3F137793",
    x"3F137CB6",
    x"3F1381D9",
    x"3F1386FB",
    x"3F138C1E",
    x"3F139140",
    x"3F139663",
    x"3F139B85",
    x"3F13A0A7",
    x"3F13A5C9",
    x"3F13AAEB",
    x"3F13B00D",
    x"3F13B52F",
    x"3F13BA50",
    x"3F13BF72",
    x"3F13C493",
    x"3F13C9B5",
    x"3F13CED6",
    x"3F13D3F8",
    x"3F13D919",
    x"3F13DE3A",
    x"3F13E35B",
    x"3F13E87C",
    x"3F13ED9C",
    x"3F13F2BD",
    x"3F13F7DE",
    x"3F13FCFE",
    x"3F14021F",
    x"3F14073F",
    x"3F140C5F",
    x"3F141180",
    x"3F1416A0",
    x"3F141BC0",
    x"3F1420E0",
    x"3F142600",
    x"3F142B1F",
    x"3F14303F",
    x"3F14355E",
    x"3F143A7E",
    x"3F143F9D",
    x"3F1444BD",
    x"3F1449DC",
    x"3F144EFB",
    x"3F14541A",
    x"3F145939",
    x"3F145E58",
    x"3F146377",
    x"3F146895",
    x"3F146DB4",
    x"3F1472D2",
    x"3F1477F1",
    x"3F147D0F",
    x"3F14822D",
    x"3F14874B",
    x"3F148C69",
    x"3F149187",
    x"3F1496A5",
    x"3F149BC3",
    x"3F14A0E1",
    x"3F14A5FE",
    x"3F14AB1C",
    x"3F14B039",
    x"3F14B557",
    x"3F14BA74",
    x"3F14BF91",
    x"3F14C4AE",
    x"3F14C9CB",
    x"3F14CEE8",
    x"3F14D405",
    x"3F14D921",
    x"3F14DE3E",
    x"3F14E35A",
    x"3F14E877",
    x"3F14ED93",
    x"3F14F2B0",
    x"3F14F7CC",
    x"3F14FCE8",
    x"3F150204",
    x"3F150720",
    x"3F150C3B",
    x"3F151157",
    x"3F151673",
    x"3F151B8E",
    x"3F1520AA",
    x"3F1525C5",
    x"3F152AE0",
    x"3F152FFC",
    x"3F153517",
    x"3F153A32",
    x"3F153F4D",
    x"3F154467",
    x"3F154982",
    x"3F154E9D",
    x"3F1553B7",
    x"3F1558D2",
    x"3F155DEC",
    x"3F156306",
    x"3F156821",
    x"3F156D3B",
    x"3F157255",
    x"3F15776F",
    x"3F157C88",
    x"3F1581A2",
    x"3F1586BC",
    x"3F158BD5",
    x"3F1590EF",
    x"3F159608",
    x"3F159B21",
    x"3F15A03B",
    x"3F15A554",
    x"3F15AA6D",
    x"3F15AF86",
    x"3F15B49F",
    x"3F15B9B7",
    x"3F15BED0",
    x"3F15C3E9",
    x"3F15C901",
    x"3F15CE19",
    x"3F15D332",
    x"3F15D84A",
    x"3F15DD62",
    x"3F15E27A",
    x"3F15E792",
    x"3F15ECAA",
    x"3F15F1C2",
    x"3F15F6D9",
    x"3F15FBF1",
    x"3F160108",
    x"3F160620",
    x"3F160B37",
    x"3F16104E",
    x"3F161565",
    x"3F161A7C",
    x"3F161F93",
    x"3F1624AA",
    x"3F1629C1",
    x"3F162ED8",
    x"3F1633EE",
    x"3F163905",
    x"3F163E1B",
    x"3F164331",
    x"3F164847",
    x"3F164D5E",
    x"3F165274",
    x"3F16578A",
    x"3F165C9F",
    x"3F1661B5",
    x"3F1666CB",
    x"3F166BE0",
    x"3F1670F6",
    x"3F16760B",
    x"3F167B21",
    x"3F168036",
    x"3F16854B",
    x"3F168A60",
    x"3F168F75",
    x"3F16948A",
    x"3F16999F",
    x"3F169EB3",
    x"3F16A3C8",
    x"3F16A8DC",
    x"3F16ADF1",
    x"3F16B305",
    x"3F16B819",
    x"3F16BD2D",
    x"3F16C241",
    x"3F16C755",
    x"3F16CC69",
    x"3F16D17D",
    x"3F16D691",
    x"3F16DBA4",
    x"3F16E0B8",
    x"3F16E5CB",
    x"3F16EADE",
    x"3F16EFF2",
    x"3F16F505",
    x"3F16FA18",
    x"3F16FF2B",
    x"3F17043E",
    x"3F170950",
    x"3F170E63",
    x"3F171376",
    x"3F171888",
    x"3F171D9B",
    x"3F1722AD",
    x"3F1727BF",
    x"3F172CD1",
    x"3F1731E3",
    x"3F1736F5",
    x"3F173C07",
    x"3F174119",
    x"3F17462B",
    x"3F174B3C",
    x"3F17504E",
    x"3F17555F",
    x"3F175A70",
    x"3F175F82",
    x"3F176493",
    x"3F1769A4",
    x"3F176EB5",
    x"3F1773C6",
    x"3F1778D6",
    x"3F177DE7",
    x"3F1782F8",
    x"3F178808",
    x"3F178D18",
    x"3F179229",
    x"3F179739",
    x"3F179C49",
    x"3F17A159",
    x"3F17A669",
    x"3F17AB79",
    x"3F17B089",
    x"3F17B598",
    x"3F17BAA8",
    x"3F17BFB7",
    x"3F17C4C7",
    x"3F17C9D6",
    x"3F17CEE5",
    x"3F17D3F4",
    x"3F17D903",
    x"3F17DE12",
    x"3F17E321",
    x"3F17E830",
    x"3F17ED3F",
    x"3F17F24D",
    x"3F17F75C",
    x"3F17FC6A",
    x"3F180178",
    x"3F180687",
    x"3F180B95",
    x"3F1810A3",
    x"3F1815B1",
    x"3F181ABE",
    x"3F181FCC",
    x"3F1824DA",
    x"3F1829E7",
    x"3F182EF5",
    x"3F183402",
    x"3F183910",
    x"3F183E1D",
    x"3F18432A",
    x"3F184837",
    x"3F184D44",
    x"3F185251",
    x"3F18575D",
    x"3F185C6A",
    x"3F186177",
    x"3F186683",
    x"3F186B8F",
    x"3F18709C",
    x"3F1875A8",
    x"3F187AB4",
    x"3F187FC0",
    x"3F1884CC",
    x"3F1889D8",
    x"3F188EE3",
    x"3F1893EF",
    x"3F1898FB",
    x"3F189E06",
    x"3F18A311",
    x"3F18A81D",
    x"3F18AD28",
    x"3F18B233",
    x"3F18B73E",
    x"3F18BC49",
    x"3F18C154",
    x"3F18C65E",
    x"3F18CB69",
    x"3F18D073",
    x"3F18D57E",
    x"3F18DA88",
    x"3F18DF92",
    x"3F18E49D",
    x"3F18E9A7",
    x"3F18EEB1",
    x"3F18F3BB",
    x"3F18F8C4",
    x"3F18FDCE",
    x"3F1902D8",
    x"3F1907E1",
    x"3F190CEB",
    x"3F1911F4",
    x"3F1916FD",
    x"3F191C06",
    x"3F19210F",
    x"3F192618",
    x"3F192B21",
    x"3F19302A",
    x"3F193533",
    x"3F193A3B",
    x"3F193F44",
    x"3F19444C",
    x"3F194955",
    x"3F194E5D",
    x"3F195365",
    x"3F19586D",
    x"3F195D75",
    x"3F19627D",
    x"3F196784",
    x"3F196C8C",
    x"3F197194",
    x"3F19769B",
    x"3F197BA3",
    x"3F1980AA",
    x"3F1985B1",
    x"3F198AB8",
    x"3F198FBF",
    x"3F1994C6",
    x"3F1999CD",
    x"3F199ED4",
    x"3F19A3DA",
    x"3F19A8E1",
    x"3F19ADE7",
    x"3F19B2EE",
    x"3F19B7F4",
    x"3F19BCFA",
    x"3F19C200",
    x"3F19C706",
    x"3F19CC0C",
    x"3F19D112",
    x"3F19D618",
    x"3F19DB1E",
    x"3F19E023",
    x"3F19E529",
    x"3F19EA2E",
    x"3F19EF33",
    x"3F19F438",
    x"3F19F93D",
    x"3F19FE42",
    x"3F1A0347",
    x"3F1A084C",
    x"3F1A0D51",
    x"3F1A1255",
    x"3F1A175A",
    x"3F1A1C5E",
    x"3F1A2163",
    x"3F1A2667",
    x"3F1A2B6B",
    x"3F1A306F",
    x"3F1A3573",
    x"3F1A3A77",
    x"3F1A3F7B",
    x"3F1A447E",
    x"3F1A4982",
    x"3F1A4E86",
    x"3F1A5389",
    x"3F1A588C",
    x"3F1A5D8F",
    x"3F1A6293",
    x"3F1A6796",
    x"3F1A6C99",
    x"3F1A719B",
    x"3F1A769E",
    x"3F1A7BA1",
    x"3F1A80A3",
    x"3F1A85A6",
    x"3F1A8AA8",
    x"3F1A8FAB",
    x"3F1A94AD",
    x"3F1A99AF",
    x"3F1A9EB1",
    x"3F1AA3B3",
    x"3F1AA8B5",
    x"3F1AADB6",
    x"3F1AB2B8",
    x"3F1AB7BA",
    x"3F1ABCBB",
    x"3F1AC1BC",
    x"3F1AC6BE",
    x"3F1ACBBF",
    x"3F1AD0C0",
    x"3F1AD5C1",
    x"3F1ADAC2",
    x"3F1ADFC3",
    x"3F1AE4C3",
    x"3F1AE9C4",
    x"3F1AEEC4",
    x"3F1AF3C5",
    x"3F1AF8C5",
    x"3F1AFDC5",
    x"3F1B02C6",
    x"3F1B07C6",
    x"3F1B0CC6",
    x"3F1B11C5",
    x"3F1B16C5",
    x"3F1B1BC5",
    x"3F1B20C4",
    x"3F1B25C4",
    x"3F1B2AC3",
    x"3F1B2FC3",
    x"3F1B34C2",
    x"3F1B39C1",
    x"3F1B3EC0",
    x"3F1B43BF",
    x"3F1B48BE",
    x"3F1B4DBD",
    x"3F1B52BB",
    x"3F1B57BA",
    x"3F1B5CB8",
    x"3F1B61B7",
    x"3F1B66B5",
    x"3F1B6BB3",
    x"3F1B70B1",
    x"3F1B75AF",
    x"3F1B7AAD",
    x"3F1B7FAB",
    x"3F1B84A9",
    x"3F1B89A6",
    x"3F1B8EA4",
    x"3F1B93A1",
    x"3F1B989E",
    x"3F1B9D9C",
    x"3F1BA299",
    x"3F1BA796",
    x"3F1BAC93",
    x"3F1BB190",
    x"3F1BB68D",
    x"3F1BBB89",
    x"3F1BC086",
    x"3F1BC582",
    x"3F1BCA7F",
    x"3F1BCF7B",
    x"3F1BD477",
    x"3F1BD973",
    x"3F1BDE6F",
    x"3F1BE36B",
    x"3F1BE867",
    x"3F1BED63",
    x"3F1BF25F",
    x"3F1BF75A",
    x"3F1BFC56",
    x"3F1C0151",
    x"3F1C064C",
    x"3F1C0B47",
    x"3F1C1042",
    x"3F1C153D",
    x"3F1C1A38",
    x"3F1C1F33",
    x"3F1C242E",
    x"3F1C2929",
    x"3F1C2E23",
    x"3F1C331D",
    x"3F1C3818",
    x"3F1C3D12",
    x"3F1C420C",
    x"3F1C4706",
    x"3F1C4C00",
    x"3F1C50FA",
    x"3F1C55F4",
    x"3F1C5AEE",
    x"3F1C5FE7",
    x"3F1C64E1",
    x"3F1C69DA",
    x"3F1C6ED3",
    x"3F1C73CC",
    x"3F1C78C6",
    x"3F1C7DBF",
    x"3F1C82B8",
    x"3F1C87B0",
    x"3F1C8CA9",
    x"3F1C91A2",
    x"3F1C969A",
    x"3F1C9B93",
    x"3F1CA08B",
    x"3F1CA583",
    x"3F1CAA7C",
    x"3F1CAF74",
    x"3F1CB46C",
    x"3F1CB963",
    x"3F1CBE5B",
    x"3F1CC353",
    x"3F1CC84B",
    x"3F1CCD42",
    x"3F1CD239",
    x"3F1CD731",
    x"3F1CDC28",
    x"3F1CE11F",
    x"3F1CE616",
    x"3F1CEB0D",
    x"3F1CF004",
    x"3F1CF4FB",
    x"3F1CF9F1",
    x"3F1CFEE8",
    x"3F1D03DE",
    x"3F1D08D5",
    x"3F1D0DCB",
    x"3F1D12C1",
    x"3F1D17B7",
    x"3F1D1CAD",
    x"3F1D21A3",
    x"3F1D2699",
    x"3F1D2B8F",
    x"3F1D3084",
    x"3F1D357A",
    x"3F1D3A6F",
    x"3F1D3F65",
    x"3F1D445A",
    x"3F1D494F",
    x"3F1D4E44",
    x"3F1D5339",
    x"3F1D582E",
    x"3F1D5D23",
    x"3F1D6217",
    x"3F1D670C",
    x"3F1D6C00",
    x"3F1D70F5",
    x"3F1D75E9",
    x"3F1D7ADD",
    x"3F1D7FD1",
    x"3F1D84C5",
    x"3F1D89B9",
    x"3F1D8EAD",
    x"3F1D93A1",
    x"3F1D9894",
    x"3F1D9D88",
    x"3F1DA27B",
    x"3F1DA76F",
    x"3F1DAC62",
    x"3F1DB155",
    x"3F1DB648",
    x"3F1DBB3B",
    x"3F1DC02E",
    x"3F1DC521",
    x"3F1DCA13",
    x"3F1DCF06",
    x"3F1DD3F8",
    x"3F1DD8EB",
    x"3F1DDDDD",
    x"3F1DE2CF",
    x"3F1DE7C1",
    x"3F1DECB3",
    x"3F1DF1A5",
    x"3F1DF697",
    x"3F1DFB89",
    x"3F1E007B",
    x"3F1E056C",
    x"3F1E0A5D",
    x"3F1E0F4F",
    x"3F1E1440",
    x"3F1E1931",
    x"3F1E1E22",
    x"3F1E2313",
    x"3F1E2804",
    x"3F1E2CF5",
    x"3F1E31E6",
    x"3F1E36D6",
    x"3F1E3BC7",
    x"3F1E40B7",
    x"3F1E45A7",
    x"3F1E4A98",
    x"3F1E4F88",
    x"3F1E5478",
    x"3F1E5968",
    x"3F1E5E57",
    x"3F1E6347",
    x"3F1E6837",
    x"3F1E6D26",
    x"3F1E7216",
    x"3F1E7705",
    x"3F1E7BF4",
    x"3F1E80E3",
    x"3F1E85D2",
    x"3F1E8AC1",
    x"3F1E8FB0",
    x"3F1E949F",
    x"3F1E998E",
    x"3F1E9E7C",
    x"3F1EA36B",
    x"3F1EA859",
    x"3F1EAD47",
    x"3F1EB236",
    x"3F1EB724",
    x"3F1EBC12",
    x"3F1EC100",
    x"3F1EC5ED",
    x"3F1ECADB",
    x"3F1ECFC9",
    x"3F1ED4B6",
    x"3F1ED9A4",
    x"3F1EDE91",
    x"3F1EE37E",
    x"3F1EE86C",
    x"3F1EED59",
    x"3F1EF245",
    x"3F1EF732",
    x"3F1EFC1F",
    x"3F1F010C",
    x"3F1F05F8",
    x"3F1F0AE5",
    x"3F1F0FD1",
    x"3F1F14BD",
    x"3F1F19AA",
    x"3F1F1E96",
    x"3F1F2382",
    x"3F1F286E",
    x"3F1F2D59",
    x"3F1F3245",
    x"3F1F3731",
    x"3F1F3C1C",
    x"3F1F4108",
    x"3F1F45F3",
    x"3F1F4ADE",
    x"3F1F4FC9",
    x"3F1F54B4",
    x"3F1F599F",
    x"3F1F5E8A",
    x"3F1F6375",
    x"3F1F6860",
    x"3F1F6D4A",
    x"3F1F7235",
    x"3F1F771F",
    x"3F1F7C09",
    x"3F1F80F3",
    x"3F1F85DD",
    x"3F1F8AC7",
    x"3F1F8FB1",
    x"3F1F949B",
    x"3F1F9985",
    x"3F1F9E6E",
    x"3F1FA358",
    x"3F1FA841",
    x"3F1FAD2B",
    x"3F1FB214",
    x"3F1FB6FD",
    x"3F1FBBE6",
    x"3F1FC0CF",
    x"3F1FC5B8",
    x"3F1FCAA0",
    x"3F1FCF89",
    x"3F1FD472",
    x"3F1FD95A",
    x"3F1FDE42",
    x"3F1FE32B",
    x"3F1FE813",
    x"3F1FECFB",
    x"3F1FF1E3",
    x"3F1FF6CB",
    x"3F1FFBB2",
    x"3F20009A",
    x"3F200582",
    x"3F200A69",
    x"3F200F50",
    x"3F201438",
    x"3F20191F",
    x"3F201E06",
    x"3F2022ED",
    x"3F2027D4",
    x"3F202CBB",
    x"3F2031A1",
    x"3F203688",
    x"3F203B6F",
    x"3F204055",
    x"3F20453B",
    x"3F204A21",
    x"3F204F08",
    x"3F2053EE",
    x"3F2058D4",
    x"3F205DB9",
    x"3F20629F",
    x"3F206785",
    x"3F206C6A",
    x"3F207150",
    x"3F207635",
    x"3F207B1A",
    x"3F208000",
    x"3F2084E5",
    x"3F2089CA",
    x"3F208EAE",
    x"3F209393",
    x"3F209878",
    x"3F209D5C",
    x"3F20A241",
    x"3F20A725",
    x"3F20AC0A",
    x"3F20B0EE",
    x"3F20B5D2",
    x"3F20BAB6",
    x"3F20BF9A",
    x"3F20C47E",
    x"3F20C961",
    x"3F20CE45",
    x"3F20D328",
    x"3F20D80C",
    x"3F20DCEF",
    x"3F20E1D2",
    x"3F20E6B5",
    x"3F20EB99",
    x"3F20F07B",
    x"3F20F55E",
    x"3F20FA41",
    x"3F20FF24",
    x"3F210406",
    x"3F2108E9",
    x"3F210DCB",
    x"3F2112AD",
    x"3F21178F",
    x"3F211C71",
    x"3F212153",
    x"3F212635",
    x"3F212B17",
    x"3F212FF9",
    x"3F2134DA",
    x"3F2139BC",
    x"3F213E9D",
    x"3F21437E",
    x"3F214860",
    x"3F214D41",
    x"3F215222",
    x"3F215703",
    x"3F215BE3",
    x"3F2160C4",
    x"3F2165A5",
    x"3F216A85",
    x"3F216F66",
    x"3F217446",
    x"3F217926",
    x"3F217E06",
    x"3F2182E6",
    x"3F2187C6",
    x"3F218CA6",
    x"3F219186",
    x"3F219665",
    x"3F219B45",
    x"3F21A024",
    x"3F21A504",
    x"3F21A9E3",
    x"3F21AEC2",
    x"3F21B3A1",
    x"3F21B880",
    x"3F21BD5F",
    x"3F21C23E",
    x"3F21C71C",
    x"3F21CBFB",
    x"3F21D0D9",
    x"3F21D5B8",
    x"3F21DA96",
    x"3F21DF74",
    x"3F21E452",
    x"3F21E930",
    x"3F21EE0E",
    x"3F21F2EC",
    x"3F21F7C9",
    x"3F21FCA7",
    x"3F220185",
    x"3F220662",
    x"3F220B3F",
    x"3F22101C",
    x"3F2214FA",
    x"3F2219D7",
    x"3F221EB3",
    x"3F222390",
    x"3F22286D",
    x"3F222D4A",
    x"3F223226",
    x"3F223702",
    x"3F223BDF",
    x"3F2240BB",
    x"3F224597",
    x"3F224A73",
    x"3F224F4F",
    x"3F22542B",
    x"3F225907",
    x"3F225DE2",
    x"3F2262BE",
    x"3F226799",
    x"3F226C74",
    x"3F227150",
    x"3F22762B",
    x"3F227B06",
    x"3F227FE1",
    x"3F2284BC",
    x"3F228996",
    x"3F228E71",
    x"3F22934C",
    x"3F229826",
    x"3F229D00",
    x"3F22A1DB",
    x"3F22A6B5",
    x"3F22AB8F",
    x"3F22B069",
    x"3F22B543",
    x"3F22BA1D",
    x"3F22BEF6",
    x"3F22C3D0",
    x"3F22C8A9",
    x"3F22CD83",
    x"3F22D25C",
    x"3F22D735",
    x"3F22DC0E",
    x"3F22E0E7",
    x"3F22E5C0",
    x"3F22EA99",
    x"3F22EF72",
    x"3F22F44A",
    x"3F22F923",
    x"3F22FDFB",
    x"3F2302D3",
    x"3F2307AB",
    x"3F230C84",
    x"3F23115C",
    x"3F231633",
    x"3F231B0B",
    x"3F231FE3",
    x"3F2324BB",
    x"3F232992",
    x"3F232E6A",
    x"3F233341",
    x"3F233818",
    x"3F233CEF",
    x"3F2341C6",
    x"3F23469D",
    x"3F234B74",
    x"3F23504B",
    x"3F235521",
    x"3F2359F8",
    x"3F235ECE",
    x"3F2363A5",
    x"3F23687B",
    x"3F236D51",
    x"3F237227",
    x"3F2376FD",
    x"3F237BD3",
    x"3F2380A8",
    x"3F23857E",
    x"3F238A54",
    x"3F238F29",
    x"3F2393FE",
    x"3F2398D4",
    x"3F239DA9",
    x"3F23A27E",
    x"3F23A753",
    x"3F23AC28",
    x"3F23B0FC",
    x"3F23B5D1",
    x"3F23BAA6",
    x"3F23BF7A",
    x"3F23C44F",
    x"3F23C923",
    x"3F23CDF7",
    x"3F23D2CB",
    x"3F23D79F",
    x"3F23DC73",
    x"3F23E147",
    x"3F23E61A",
    x"3F23EAEE",
    x"3F23EFC1",
    x"3F23F495",
    x"3F23F968",
    x"3F23FE3B",
    x"3F24030E",
    x"3F2407E1",
    x"3F240CB4",
    x"3F241187",
    x"3F24165A",
    x"3F241B2C",
    x"3F241FFF",
    x"3F2424D1",
    x"3F2429A3",
    x"3F242E75",
    x"3F243348",
    x"3F24381A",
    x"3F243CEB",
    x"3F2441BD",
    x"3F24468F",
    x"3F244B60",
    x"3F245032",
    x"3F245503",
    x"3F2459D5",
    x"3F245EA6",
    x"3F246377",
    x"3F246848",
    x"3F246D19",
    x"3F2471EA",
    x"3F2476BA",
    x"3F247B8B",
    x"3F24805B",
    x"3F24852C",
    x"3F2489FC",
    x"3F248ECC",
    x"3F24939C",
    x"3F24986D",
    x"3F249D3C",
    x"3F24A20C",
    x"3F24A6DC",
    x"3F24ABAC",
    x"3F24B07B",
    x"3F24B54A",
    x"3F24BA1A",
    x"3F24BEE9",
    x"3F24C3B8",
    x"3F24C887",
    x"3F24CD56",
    x"3F24D225",
    x"3F24D6F4",
    x"3F24DBC2",
    x"3F24E091",
    x"3F24E55F",
    x"3F24EA2D",
    x"3F24EEFC",
    x"3F24F3CA",
    x"3F24F898",
    x"3F24FD66",
    x"3F250234",
    x"3F250701",
    x"3F250BCF",
    x"3F25109C",
    x"3F25156A",
    x"3F251A37",
    x"3F251F04",
    x"3F2523D2",
    x"3F25289F",
    x"3F252D6C",
    x"3F253238",
    x"3F253705",
    x"3F253BD2",
    x"3F25409E",
    x"3F25456B",
    x"3F254A37",
    x"3F254F03",
    x"3F2553CF",
    x"3F25589B",
    x"3F255D67",
    x"3F256233",
    x"3F2566FF",
    x"3F256BCB",
    x"3F257096",
    x"3F257562",
    x"3F257A2D",
    x"3F257EF8",
    x"3F2583C3",
    x"3F25888E",
    x"3F258D59",
    x"3F259224",
    x"3F2596EF",
    x"3F259BB9",
    x"3F25A084",
    x"3F25A54E",
    x"3F25AA19",
    x"3F25AEE3",
    x"3F25B3AD",
    x"3F25B877",
    x"3F25BD41",
    x"3F25C20B",
    x"3F25C6D5",
    x"3F25CB9E",
    x"3F25D068",
    x"3F25D531",
    x"3F25D9FB",
    x"3F25DEC4",
    x"3F25E38D",
    x"3F25E856",
    x"3F25ED1F",
    x"3F25F1E8",
    x"3F25F6B1",
    x"3F25FB79",
    x"3F260042",
    x"3F26050A",
    x"3F2609D3",
    x"3F260E9B",
    x"3F261363",
    x"3F26182B",
    x"3F261CF3",
    x"3F2621BB",
    x"3F262682",
    x"3F262B4A",
    x"3F263012",
    x"3F2634D9",
    x"3F2639A0",
    x"3F263E68",
    x"3F26432F",
    x"3F2647F6",
    x"3F264CBD",
    x"3F265184",
    x"3F26564A",
    x"3F265B11",
    x"3F265FD8",
    x"3F26649E",
    x"3F266964",
    x"3F266E2B",
    x"3F2672F1",
    x"3F2677B7",
    x"3F267C7D",
    x"3F268143",
    x"3F268608",
    x"3F268ACE",
    x"3F268F93",
    x"3F269459",
    x"3F26991E",
    x"3F269DE3",
    x"3F26A2A9",
    x"3F26A76E",
    x"3F26AC33",
    x"3F26B0F7",
    x"3F26B5BC",
    x"3F26BA81",
    x"3F26BF45",
    x"3F26C40A",
    x"3F26C8CE",
    x"3F26CD92",
    x"3F26D256",
    x"3F26D71A",
    x"3F26DBDE",
    x"3F26E0A2",
    x"3F26E566",
    x"3F26EA2A",
    x"3F26EEED",
    x"3F26F3B0",
    x"3F26F874",
    x"3F26FD37",
    x"3F2701FA",
    x"3F2706BD",
    x"3F270B80",
    x"3F271043",
    x"3F271506",
    x"3F2719C8",
    x"3F271E8B",
    x"3F27234D",
    x"3F272810",
    x"3F272CD2",
    x"3F273194",
    x"3F273656",
    x"3F273B18",
    x"3F273FDA",
    x"3F27449B",
    x"3F27495D",
    x"3F274E1E",
    x"3F2752E0",
    x"3F2757A1",
    x"3F275C62",
    x"3F276123",
    x"3F2765E5",
    x"3F276AA5",
    x"3F276F66",
    x"3F277427",
    x"3F2778E8",
    x"3F277DA8",
    x"3F278268",
    x"3F278729",
    x"3F278BE9",
    x"3F2790A9",
    x"3F279569",
    x"3F279A29",
    x"3F279EE9",
    x"3F27A3A8",
    x"3F27A868",
    x"3F27AD28",
    x"3F27B1E7",
    x"3F27B6A6",
    x"3F27BB65",
    x"3F27C025",
    x"3F27C4E4",
    x"3F27C9A2",
    x"3F27CE61",
    x"3F27D320",
    x"3F27D7DE",
    x"3F27DC9D",
    x"3F27E15B",
    x"3F27E61A",
    x"3F27EAD8",
    x"3F27EF96",
    x"3F27F454",
    x"3F27F912",
    x"3F27FDD0",
    x"3F28028D",
    x"3F28074B",
    x"3F280C08",
    x"3F2810C6",
    x"3F281583",
    x"3F281A40",
    x"3F281EFD",
    x"3F2823BA",
    x"3F282877",
    x"3F282D34",
    x"3F2831F0",
    x"3F2836AD",
    x"3F283B69",
    x"3F284026",
    x"3F2844E2",
    x"3F28499E",
    x"3F284E5A",
    x"3F285316",
    x"3F2857D2",
    x"3F285C8E",
    x"3F286149",
    x"3F286605",
    x"3F286AC0",
    x"3F286F7C",
    x"3F287437",
    x"3F2878F2",
    x"3F287DAD",
    x"3F288268",
    x"3F288723",
    x"3F288BDE",
    x"3F289098",
    x"3F289553",
    x"3F289A0D",
    x"3F289EC8",
    x"3F28A382",
    x"3F28A83C",
    x"3F28ACF6",
    x"3F28B1B0",
    x"3F28B66A",
    x"3F28BB23",
    x"3F28BFDD",
    x"3F28C497",
    x"3F28C950",
    x"3F28CE09",
    x"3F28D2C3",
    x"3F28D77C",
    x"3F28DC35",
    x"3F28E0EE",
    x"3F28E5A6",
    x"3F28EA5F",
    x"3F28EF18",
    x"3F28F3D0",
    x"3F28F889",
    x"3F28FD41",
    x"3F2901F9",
    x"3F2906B1",
    x"3F290B69",
    x"3F291021",
    x"3F2914D9",
    x"3F291991",
    x"3F291E48",
    x"3F292300",
    x"3F2927B7",
    x"3F292C6E",
    x"3F293125",
    x"3F2935DD",
    x"3F293A93",
    x"3F293F4A",
    x"3F294401",
    x"3F2948B8",
    x"3F294D6E",
    x"3F295225",
    x"3F2956DB",
    x"3F295B91",
    x"3F296048",
    x"3F2964FE",
    x"3F2969B4",
    x"3F296E69",
    x"3F29731F",
    x"3F2977D5",
    x"3F297C8A",
    x"3F298140",
    x"3F2985F5",
    x"3F298AAA",
    x"3F298F60",
    x"3F299415",
    x"3F2998CA",
    x"3F299D7E",
    x"3F29A233",
    x"3F29A6E8",
    x"3F29AB9C",
    x"3F29B051",
    x"3F29B505",
    x"3F29B9B9",
    x"3F29BE6D",
    x"3F29C321",
    x"3F29C7D5",
    x"3F29CC89",
    x"3F29D13D",
    x"3F29D5F0",
    x"3F29DAA4",
    x"3F29DF57",
    x"3F29E40B",
    x"3F29E8BE",
    x"3F29ED71",
    x"3F29F224",
    x"3F29F6D7",
    x"3F29FB89",
    x"3F2A003C",
    x"3F2A04EF",
    x"3F2A09A1",
    x"3F2A0E54",
    x"3F2A1306",
    x"3F2A17B8",
    x"3F2A1C6A",
    x"3F2A211C",
    x"3F2A25CE",
    x"3F2A2A80",
    x"3F2A2F31",
    x"3F2A33E3",
    x"3F2A3894",
    x"3F2A3D46",
    x"3F2A41F7",
    x"3F2A46A8",
    x"3F2A4B59",
    x"3F2A500A",
    x"3F2A54BB",
    x"3F2A596C",
    x"3F2A5E1C",
    x"3F2A62CD",
    x"3F2A677D",
    x"3F2A6C2E",
    x"3F2A70DE",
    x"3F2A758E",
    x"3F2A7A3E",
    x"3F2A7EEE",
    x"3F2A839E",
    x"3F2A884D",
    x"3F2A8CFD",
    x"3F2A91AC",
    x"3F2A965C",
    x"3F2A9B0B",
    x"3F2A9FBA",
    x"3F2AA469",
    x"3F2AA918",
    x"3F2AADC7",
    x"3F2AB276",
    x"3F2AB725",
    x"3F2ABBD3",
    x"3F2AC082",
    x"3F2AC530",
    x"3F2AC9DE",
    x"3F2ACE8D",
    x"3F2AD33B",
    x"3F2AD7E9",
    x"3F2ADC96",
    x"3F2AE144",
    x"3F2AE5F2",
    x"3F2AEA9F",
    x"3F2AEF4D",
    x"3F2AF3FA",
    x"3F2AF8A7",
    x"3F2AFD55",
    x"3F2B0202",
    x"3F2B06AF",
    x"3F2B0B5B",
    x"3F2B1008",
    x"3F2B14B5",
    x"3F2B1961",
    x"3F2B1E0E",
    x"3F2B22BA",
    x"3F2B2766",
    x"3F2B2C12",
    x"3F2B30BE",
    x"3F2B356A",
    x"3F2B3A16",
    x"3F2B3EC2",
    x"3F2B436D",
    x"3F2B4819",
    x"3F2B4CC4",
    x"3F2B516F",
    x"3F2B561B",
    x"3F2B5AC6",
    x"3F2B5F71",
    x"3F2B641B",
    x"3F2B68C6",
    x"3F2B6D71",
    x"3F2B721B",
    x"3F2B76C6",
    x"3F2B7B70",
    x"3F2B801A",
    x"3F2B84C5",
    x"3F2B896F",
    x"3F2B8E19",
    x"3F2B92C2",
    x"3F2B976C",
    x"3F2B9C16",
    x"3F2BA0BF",
    x"3F2BA569",
    x"3F2BAA12",
    x"3F2BAEBB",
    x"3F2BB364",
    x"3F2BB80D",
    x"3F2BBCB6",
    x"3F2BC15F",
    x"3F2BC608",
    x"3F2BCAB0",
    x"3F2BCF59",
    x"3F2BD401",
    x"3F2BD8AA",
    x"3F2BDD52",
    x"3F2BE1FA",
    x"3F2BE6A2",
    x"3F2BEB4A",
    x"3F2BEFF1",
    x"3F2BF499",
    x"3F2BF941",
    x"3F2BFDE8",
    x"3F2C028F",
    x"3F2C0737",
    x"3F2C0BDE",
    x"3F2C1085",
    x"3F2C152C",
    x"3F2C19D3",
    x"3F2C1E79",
    x"3F2C2320",
    x"3F2C27C7",
    x"3F2C2C6D",
    x"3F2C3113",
    x"3F2C35B9",
    x"3F2C3A60",
    x"3F2C3F06",
    x"3F2C43AB",
    x"3F2C4851",
    x"3F2C4CF7",
    x"3F2C519D",
    x"3F2C5642",
    x"3F2C5AE7",
    x"3F2C5F8D",
    x"3F2C6432",
    x"3F2C68D7",
    x"3F2C6D7C",
    x"3F2C7221",
    x"3F2C76C5",
    x"3F2C7B6A",
    x"3F2C800F",
    x"3F2C84B3",
    x"3F2C8957",
    x"3F2C8DFC",
    x"3F2C92A0",
    x"3F2C9744",
    x"3F2C9BE8",
    x"3F2CA08C",
    x"3F2CA52F",
    x"3F2CA9D3",
    x"3F2CAE76",
    x"3F2CB31A",
    x"3F2CB7BD",
    x"3F2CBC60",
    x"3F2CC103",
    x"3F2CC5A6",
    x"3F2CCA49",
    x"3F2CCEEC",
    x"3F2CD38F",
    x"3F2CD831",
    x"3F2CDCD4",
    x"3F2CE176",
    x"3F2CE618",
    x"3F2CEABB",
    x"3F2CEF5D",
    x"3F2CF3FF",
    x"3F2CF8A0",
    x"3F2CFD42",
    x"3F2D01E4",
    x"3F2D0685",
    x"3F2D0B27",
    x"3F2D0FC8",
    x"3F2D1469",
    x"3F2D190A",
    x"3F2D1DAB",
    x"3F2D224C",
    x"3F2D26ED",
    x"3F2D2B8E",
    x"3F2D302E",
    x"3F2D34CF",
    x"3F2D396F",
    x"3F2D3E10",
    x"3F2D42B0",
    x"3F2D4750",
    x"3F2D4BF0",
    x"3F2D5090",
    x"3F2D552F",
    x"3F2D59CF",
    x"3F2D5E6F",
    x"3F2D630E",
    x"3F2D67AD",
    x"3F2D6C4D",
    x"3F2D70EC",
    x"3F2D758B",
    x"3F2D7A2A",
    x"3F2D7EC9",
    x"3F2D8367",
    x"3F2D8806",
    x"3F2D8CA4",
    x"3F2D9143",
    x"3F2D95E1",
    x"3F2D9A7F",
    x"3F2D9F1D",
    x"3F2DA3BB",
    x"3F2DA859",
    x"3F2DACF7",
    x"3F2DB195",
    x"3F2DB632",
    x"3F2DBAD0",
    x"3F2DBF6D",
    x"3F2DC40A",
    x"3F2DC8A7",
    x"3F2DCD44",
    x"3F2DD1E1",
    x"3F2DD67E",
    x"3F2DDB1B",
    x"3F2DDFB8",
    x"3F2DE454",
    x"3F2DE8F0",
    x"3F2DED8D",
    x"3F2DF229",
    x"3F2DF6C5",
    x"3F2DFB61",
    x"3F2DFFFD",
    x"3F2E0499",
    x"3F2E0934",
    x"3F2E0DD0",
    x"3F2E126B",
    x"3F2E1707",
    x"3F2E1BA2",
    x"3F2E203D",
    x"3F2E24D8",
    x"3F2E2973",
    x"3F2E2E0E",
    x"3F2E32A9",
    x"3F2E3743",
    x"3F2E3BDE",
    x"3F2E4078",
    x"3F2E4513",
    x"3F2E49AD",
    x"3F2E4E47",
    x"3F2E52E1",
    x"3F2E577B",
    x"3F2E5C15",
    x"3F2E60AE",
    x"3F2E6548",
    x"3F2E69E1",
    x"3F2E6E7B",
    x"3F2E7314",
    x"3F2E77AD",
    x"3F2E7C46",
    x"3F2E80DF",
    x"3F2E8578",
    x"3F2E8A11",
    x"3F2E8EA9",
    x"3F2E9342",
    x"3F2E97DA",
    x"3F2E9C73",
    x"3F2EA10B",
    x"3F2EA5A3",
    x"3F2EAA3B",
    x"3F2EAED3",
    x"3F2EB36B",
    x"3F2EB802",
    x"3F2EBC9A",
    x"3F2EC131",
    x"3F2EC5C9",
    x"3F2ECA60",
    x"3F2ECEF7",
    x"3F2ED38E",
    x"3F2ED825",
    x"3F2EDCBC",
    x"3F2EE153",
    x"3F2EE5E9",
    x"3F2EEA80",
    x"3F2EEF16",
    x"3F2EF3AD",
    x"3F2EF843",
    x"3F2EFCD9",
    x"3F2F016F",
    x"3F2F0605",
    x"3F2F0A9B",
    x"3F2F0F30",
    x"3F2F13C6",
    x"3F2F185B",
    x"3F2F1CF1",
    x"3F2F2186",
    x"3F2F261B",
    x"3F2F2AB0",
    x"3F2F2F45",
    x"3F2F33DA",
    x"3F2F386F",
    x"3F2F3D03",
    x"3F2F4198",
    x"3F2F462C",
    x"3F2F4AC1",
    x"3F2F4F55",
    x"3F2F53E9",
    x"3F2F587D",
    x"3F2F5D11",
    x"3F2F61A5",
    x"3F2F6638",
    x"3F2F6ACC",
    x"3F2F6F5F",
    x"3F2F73F3",
    x"3F2F7886",
    x"3F2F7D19",
    x"3F2F81AC",
    x"3F2F863F",
    x"3F2F8AD2",
    x"3F2F8F65",
    x"3F2F93F7",
    x"3F2F988A",
    x"3F2F9D1C",
    x"3F2FA1AF",
    x"3F2FA641",
    x"3F2FAAD3",
    x"3F2FAF65",
    x"3F2FB3F7",
    x"3F2FB888",
    x"3F2FBD1A",
    x"3F2FC1AC",
    x"3F2FC63D",
    x"3F2FCACF",
    x"3F2FCF60",
    x"3F2FD3F1",
    x"3F2FD882",
    x"3F2FDD13",
    x"3F2FE1A4",
    x"3F2FE634",
    x"3F2FEAC5",
    x"3F2FEF56",
    x"3F2FF3E6",
    x"3F2FF876",
    x"3F2FFD06",
    x"3F300196",
    x"3F300626",
    x"3F300AB6",
    x"3F300F46",
    x"3F3013D6",
    x"3F301865",
    x"3F301CF5",
    x"3F302184",
    x"3F302613",
    x"3F302AA2",
    x"3F302F31",
    x"3F3033C0",
    x"3F30384F",
    x"3F303CDE",
    x"3F30416C",
    x"3F3045FB",
    x"3F304A89",
    x"3F304F18",
    x"3F3053A6",
    x"3F305834",
    x"3F305CC2",
    x"3F306150",
    x"3F3065DD",
    x"3F306A6B",
    x"3F306EF9",
    x"3F307386",
    x"3F307813",
    x"3F307CA1",
    x"3F30812E",
    x"3F3085BB",
    x"3F308A48",
    x"3F308ED4",
    x"3F309361",
    x"3F3097EE",
    x"3F309C7A",
    x"3F30A106",
    x"3F30A593",
    x"3F30AA1F",
    x"3F30AEAB",
    x"3F30B337",
    x"3F30B7C3",
    x"3F30BC4E",
    x"3F30C0DA",
    x"3F30C566",
    x"3F30C9F1",
    x"3F30CE7C",
    x"3F30D307",
    x"3F30D792",
    x"3F30DC1D",
    x"3F30E0A8",
    x"3F30E533",
    x"3F30E9BE",
    x"3F30EE48",
    x"3F30F2D3",
    x"3F30F75D",
    x"3F30FBE7",
    x"3F310071",
    x"3F3104FB",
    x"3F310985",
    x"3F310E0F",
    x"3F311299",
    x"3F311722",
    x"3F311BAC",
    x"3F312035",
    x"3F3124BF",
    x"3F312948",
    x"3F312DD1",
    x"3F31325A",
    x"3F3136E3",
    x"3F313B6B",
    x"3F313FF4",
    x"3F31447D",
    x"3F314905",
    x"3F314D8D",
    x"3F315215",
    x"3F31569E",
    x"3F315B26",
    x"3F315FAD",
    x"3F316435",
    x"3F3168BD",
    x"3F316D44",
    x"3F3171CC",
    x"3F317653",
    x"3F317ADB",
    x"3F317F62",
    x"3F3183E9",
    x"3F318870",
    x"3F318CF6",
    x"3F31917D",
    x"3F319604",
    x"3F319A8A",
    x"3F319F11",
    x"3F31A397",
    x"3F31A81D",
    x"3F31ACA3",
    x"3F31B129",
    x"3F31B5AF",
    x"3F31BA35",
    x"3F31BEBA",
    x"3F31C340",
    x"3F31C7C5",
    x"3F31CC4B",
    x"3F31D0D0",
    x"3F31D555",
    x"3F31D9DA",
    x"3F31DE5F",
    x"3F31E2E4",
    x"3F31E768",
    x"3F31EBED",
    x"3F31F071",
    x"3F31F4F6",
    x"3F31F97A",
    x"3F31FDFE",
    x"3F320282",
    x"3F320706",
    x"3F320B8A",
    x"3F32100E",
    x"3F321491",
    x"3F321915",
    x"3F321D98",
    x"3F32221B",
    x"3F32269E",
    x"3F322B22",
    x"3F322FA5",
    x"3F323427",
    x"3F3238AA",
    x"3F323D2D",
    x"3F3241AF",
    x"3F324632",
    x"3F324AB4",
    x"3F324F36",
    x"3F3253B8",
    x"3F32583A",
    x"3F325CBC",
    x"3F32613E",
    x"3F3265C0",
    x"3F326A41",
    x"3F326EC3",
    x"3F327344",
    x"3F3277C5",
    x"3F327C46",
    x"3F3280C7",
    x"3F328548",
    x"3F3289C9",
    x"3F328E4A",
    x"3F3292CA",
    x"3F32974B",
    x"3F329BCB",
    x"3F32A04C",
    x"3F32A4CC",
    x"3F32A94C",
    x"3F32ADCC",
    x"3F32B24C",
    x"3F32B6CB",
    x"3F32BB4B",
    x"3F32BFCA",
    x"3F32C44A",
    x"3F32C8C9",
    x"3F32CD48",
    x"3F32D1C7",
    x"3F32D646",
    x"3F32DAC5",
    x"3F32DF44",
    x"3F32E3C3",
    x"3F32E841",
    x"3F32ECC0",
    x"3F32F13E",
    x"3F32F5BC",
    x"3F32FA3A",
    x"3F32FEB8",
    x"3F330336",
    x"3F3307B4",
    x"3F330C32",
    x"3F3310AF",
    x"3F33152D",
    x"3F3319AA",
    x"3F331E27",
    x"3F3322A5",
    x"3F332722",
    x"3F332B9F",
    x"3F33301B",
    x"3F333498",
    x"3F333915",
    x"3F333D91",
    x"3F33420E",
    x"3F33468A",
    x"3F334B06",
    x"3F334F82",
    x"3F3353FE",
    x"3F33587A",
    x"3F335CF6",
    x"3F336171",
    x"3F3365ED",
    x"3F336A68",
    x"3F336EE4",
    x"3F33735F",
    x"3F3377DA",
    x"3F337C55",
    x"3F3380D0",
    x"3F33854B",
    x"3F3389C5",
    x"3F338E40",
    x"3F3392BA",
    x"3F339735",
    x"3F339BAF",
    x"3F33A029",
    x"3F33A4A3",
    x"3F33A91D",
    x"3F33AD97",
    x"3F33B210",
    x"3F33B68A",
    x"3F33BB03",
    x"3F33BF7D",
    x"3F33C3F6",
    x"3F33C86F",
    x"3F33CCE8",
    x"3F33D161",
    x"3F33D5DA",
    x"3F33DA53",
    x"3F33DECB",
    x"3F33E344",
    x"3F33E7BC",
    x"3F33EC34",
    x"3F33F0AD",
    x"3F33F525",
    x"3F33F99D",
    x"3F33FE14",
    x"3F34028C",
    x"3F340704",
    x"3F340B7B",
    x"3F340FF3",
    x"3F34146A",
    x"3F3418E1",
    x"3F341D58",
    x"3F3421CF",
    x"3F342646",
    x"3F342ABD",
    x"3F342F34",
    x"3F3433AA",
    x"3F343821",
    x"3F343C97",
    x"3F34410D",
    x"3F344583",
    x"3F3449F9",
    x"3F344E6F",
    x"3F3452E5",
    x"3F34575B",
    x"3F345BD0",
    x"3F346046",
    x"3F3464BB",
    x"3F346930",
    x"3F346DA5",
    x"3F34721A",
    x"3F34768F",
    x"3F347B04",
    x"3F347F79",
    x"3F3483ED",
    x"3F348862",
    x"3F348CD6",
    x"3F34914B",
    x"3F3495BF",
    x"3F349A33",
    x"3F349EA7",
    x"3F34A31B",
    x"3F34A78E",
    x"3F34AC02",
    x"3F34B075",
    x"3F34B4E9",
    x"3F34B95C",
    x"3F34BDCF",
    x"3F34C242",
    x"3F34C6B5",
    x"3F34CB28",
    x"3F34CF9B",
    x"3F34D40D",
    x"3F34D880",
    x"3F34DCF2",
    x"3F34E165",
    x"3F34E5D7",
    x"3F34EA49",
    x"3F34EEBB",
    x"3F34F32D",
    x"3F34F79F",
    x"3F34FC10",
    x"3F350082",
    x"3F3504F3",
    x"3F350965",
    x"3F350DD6",
    x"3F351247",
    x"3F3516B8",
    x"3F351B29",
    x"3F351F9A",
    x"3F35240A",
    x"3F35287B",
    x"3F352CEB",
    x"3F35315C",
    x"3F3535CC",
    x"3F353A3C",
    x"3F353EAC",
    x"3F35431C",
    x"3F35478C",
    x"3F354BFB",
    x"3F35506B",
    x"3F3554DA",
    x"3F35594A",
    x"3F355DB9",
    x"3F356228",
    x"3F356697",
    x"3F356B06",
    x"3F356F75",
    x"3F3573E4",
    x"3F357852",
    x"3F357CC1",
    x"3F35812F",
    x"3F35859D",
    x"3F358A0B",
    x"3F358E79",
    x"3F3592E7",
    x"3F359755",
    x"3F359BC3",
    x"3F35A031",
    x"3F35A49E",
    x"3F35A90B",
    x"3F35AD79",
    x"3F35B1E6",
    x"3F35B653",
    x"3F35BAC0",
    x"3F35BF2D",
    x"3F35C39A",
    x"3F35C806",
    x"3F35CC73",
    x"3F35D0DF",
    x"3F35D54B",
    x"3F35D9B8",
    x"3F35DE24",
    x"3F35E290",
    x"3F35E6FB",
    x"3F35EB67",
    x"3F35EFD3",
    x"3F35F43E",
    x"3F35F8AA",
    x"3F35FD15",
    x"3F360180",
    x"3F3605EB",
    x"3F360A56",
    x"3F360EC1",
    x"3F36132C",
    x"3F361797",
    x"3F361C01",
    x"3F36206C",
    x"3F3624D6",
    x"3F362940",
    x"3F362DAA",
    x"3F363214",
    x"3F36367E",
    x"3F363AE8",
    x"3F363F52",
    x"3F3643BB",
    x"3F364825",
    x"3F364C8E",
    x"3F3650F7",
    x"3F365560",
    x"3F3659C9",
    x"3F365E32",
    x"3F36629B",
    x"3F366704",
    x"3F366B6C",
    x"3F366FD5",
    x"3F36743D",
    x"3F3678A5",
    x"3F367D0D",
    x"3F368175",
    x"3F3685DD",
    x"3F368A45",
    x"3F368EAD",
    x"3F369314",
    x"3F36977C",
    x"3F369BE3",
    x"3F36A04A",
    x"3F36A4B2",
    x"3F36A919",
    x"3F36AD7F",
    x"3F36B1E6",
    x"3F36B64D",
    x"3F36BAB4",
    x"3F36BF1A",
    x"3F36C380",
    x"3F36C7E7",
    x"3F36CC4D",
    x"3F36D0B3",
    x"3F36D519",
    x"3F36D97F",
    x"3F36DDE4",
    x"3F36E24A",
    x"3F36E6AF",
    x"3F36EB15",
    x"3F36EF7A",
    x"3F36F3DF",
    x"3F36F844",
    x"3F36FCA9",
    x"3F37010E",
    x"3F370573",
    x"3F3709D7",
    x"3F370E3C",
    x"3F3712A0",
    x"3F371704",
    x"3F371B69",
    x"3F371FCD",
    x"3F372431",
    x"3F372894",
    x"3F372CF8",
    x"3F37315C",
    x"3F3735BF",
    x"3F373A23",
    x"3F373E86",
    x"3F3742E9",
    x"3F37474C",
    x"3F374BAF",
    x"3F375012",
    x"3F375475",
    x"3F3758D7",
    x"3F375D3A",
    x"3F37619C",
    x"3F3765FE",
    x"3F376A61",
    x"3F376EC3",
    x"3F377325",
    x"3F377787",
    x"3F377BE8",
    x"3F37804A",
    x"3F3784AB",
    x"3F37890D",
    x"3F378D6E",
    x"3F3791CF",
    x"3F379630",
    x"3F379A91",
    x"3F379EF2",
    x"3F37A353",
    x"3F37A7B4",
    x"3F37AC14",
    x"3F37B074",
    x"3F37B4D5",
    x"3F37B935",
    x"3F37BD95",
    x"3F37C1F5",
    x"3F37C655",
    x"3F37CAB5",
    x"3F37CF14",
    x"3F37D374",
    x"3F37D7D3",
    x"3F37DC32",
    x"3F37E092",
    x"3F37E4F1",
    x"3F37E950",
    x"3F37EDAF",
    x"3F37F20D",
    x"3F37F66C",
    x"3F37FACA",
    x"3F37FF29",
    x"3F380387",
    x"3F3807E5",
    x"3F380C43",
    x"3F3810A1",
    x"3F3814FF",
    x"3F38195D",
    x"3F381DBB",
    x"3F382218",
    x"3F382676",
    x"3F382AD3",
    x"3F382F30",
    x"3F38338D",
    x"3F3837EA",
    x"3F383C47",
    x"3F3840A4",
    x"3F384500",
    x"3F38495D",
    x"3F384DB9",
    x"3F385216",
    x"3F385672",
    x"3F385ACE",
    x"3F385F2A",
    x"3F386386",
    x"3F3867E1",
    x"3F386C3D",
    x"3F387099",
    x"3F3874F4",
    x"3F38794F",
    x"3F387DAB",
    x"3F388206",
    x"3F388661",
    x"3F388ABB",
    x"3F388F16",
    x"3F389371",
    x"3F3897CB",
    x"3F389C26",
    x"3F38A080",
    x"3F38A4DA",
    x"3F38A934",
    x"3F38AD8E",
    x"3F38B1E8",
    x"3F38B642",
    x"3F38BA9C",
    x"3F38BEF5",
    x"3F38C34F",
    x"3F38C7A8",
    x"3F38CC01",
    x"3F38D05A",
    x"3F38D4B3",
    x"3F38D90C",
    x"3F38DD65",
    x"3F38E1BD",
    x"3F38E616",
    x"3F38EA6E",
    x"3F38EEC7",
    x"3F38F31F",
    x"3F38F777",
    x"3F38FBCF",
    x"3F390027",
    x"3F39047E",
    x"3F3908D6",
    x"3F390D2E",
    x"3F391185",
    x"3F3915DC",
    x"3F391A33",
    x"3F391E8B",
    x"3F3922E1",
    x"3F392738",
    x"3F392B8F",
    x"3F392FE6",
    x"3F39343C",
    x"3F393893",
    x"3F393CE9",
    x"3F39413F",
    x"3F394595",
    x"3F3949EB",
    x"3F394E41",
    x"3F395297",
    x"3F3956EC",
    x"3F395B42",
    x"3F395F97",
    x"3F3963ED",
    x"3F396842",
    x"3F396C97",
    x"3F3970EC",
    x"3F397541",
    x"3F397995",
    x"3F397DEA",
    x"3F39823E",
    x"3F398693",
    x"3F398AE7",
    x"3F398F3B",
    x"3F39938F",
    x"3F3997E3",
    x"3F399C37",
    x"3F39A08B",
    x"3F39A4DF",
    x"3F39A932",
    x"3F39AD85",
    x"3F39B1D9",
    x"3F39B62C",
    x"3F39BA7F",
    x"3F39BED2",
    x"3F39C325",
    x"3F39C777",
    x"3F39CBCA",
    x"3F39D01D",
    x"3F39D46F",
    x"3F39D8C1",
    x"3F39DD13",
    x"3F39E165",
    x"3F39E5B7",
    x"3F39EA09",
    x"3F39EE5B",
    x"3F39F2AC",
    x"3F39F6FE",
    x"3F39FB4F",
    x"3F39FFA1",
    x"3F3A03F2",
    x"3F3A0843",
    x"3F3A0C94",
    x"3F3A10E4",
    x"3F3A1535",
    x"3F3A1986",
    x"3F3A1DD6",
    x"3F3A2227",
    x"3F3A2677",
    x"3F3A2AC7",
    x"3F3A2F17",
    x"3F3A3367",
    x"3F3A37B7",
    x"3F3A3C06",
    x"3F3A4056",
    x"3F3A44A6",
    x"3F3A48F5",
    x"3F3A4D44",
    x"3F3A5193",
    x"3F3A55E2",
    x"3F3A5A31",
    x"3F3A5E80",
    x"3F3A62CF",
    x"3F3A671D",
    x"3F3A6B6C",
    x"3F3A6FBA",
    x"3F3A7408",
    x"3F3A7856",
    x"3F3A7CA4",
    x"3F3A80F2",
    x"3F3A8540",
    x"3F3A898E",
    x"3F3A8DDB",
    x"3F3A9229",
    x"3F3A9676",
    x"3F3A9AC3",
    x"3F3A9F10",
    x"3F3AA35D",
    x"3F3AA7AA",
    x"3F3AABF7",
    x"3F3AB044",
    x"3F3AB490",
    x"3F3AB8DD",
    x"3F3ABD29",
    x"3F3AC175",
    x"3F3AC5C1",
    x"3F3ACA0D",
    x"3F3ACE59",
    x"3F3AD2A5",
    x"3F3AD6F1",
    x"3F3ADB3C",
    x"3F3ADF88",
    x"3F3AE3D3",
    x"3F3AE81E",
    x"3F3AEC69",
    x"3F3AF0B4",
    x"3F3AF4FF",
    x"3F3AF94A",
    x"3F3AFD94",
    x"3F3B01DF",
    x"3F3B0629",
    x"3F3B0A74",
    x"3F3B0EBE",
    x"3F3B1308",
    x"3F3B1752",
    x"3F3B1B9C",
    x"3F3B1FE5",
    x"3F3B242F",
    x"3F3B2879",
    x"3F3B2CC2",
    x"3F3B310B",
    x"3F3B3554",
    x"3F3B399E",
    x"3F3B3DE6",
    x"3F3B422F",
    x"3F3B4678",
    x"3F3B4AC1",
    x"3F3B4F09",
    x"3F3B5351",
    x"3F3B579A",
    x"3F3B5BE2",
    x"3F3B602A",
    x"3F3B6472",
    x"3F3B68BA",
    x"3F3B6D01",
    x"3F3B7149",
    x"3F3B7590",
    x"3F3B79D8",
    x"3F3B7E1F",
    x"3F3B8266",
    x"3F3B86AD",
    x"3F3B8AF4",
    x"3F3B8F3B",
    x"3F3B9382",
    x"3F3B97C8",
    x"3F3B9C0F",
    x"3F3BA055",
    x"3F3BA49B",
    x"3F3BA8E1",
    x"3F3BAD27",
    x"3F3BB16D",
    x"3F3BB5B3",
    x"3F3BB9F9",
    x"3F3BBE3E",
    x"3F3BC284",
    x"3F3BC6C9",
    x"3F3BCB0E",
    x"3F3BCF53",
    x"3F3BD398",
    x"3F3BD7DD",
    x"3F3BDC22",
    x"3F3BE067",
    x"3F3BE4AB",
    x"3F3BE8F0",
    x"3F3BED34",
    x"3F3BF178",
    x"3F3BF5BC",
    x"3F3BFA00",
    x"3F3BFE44",
    x"3F3C0288",
    x"3F3C06CB",
    x"3F3C0B0F",
    x"3F3C0F52",
    x"3F3C1396",
    x"3F3C17D9",
    x"3F3C1C1C",
    x"3F3C205F",
    x"3F3C24A2",
    x"3F3C28E4",
    x"3F3C2D27",
    x"3F3C316A",
    x"3F3C35AC",
    x"3F3C39EE",
    x"3F3C3E30",
    x"3F3C4272",
    x"3F3C46B4",
    x"3F3C4AF6",
    x"3F3C4F38",
    x"3F3C5379",
    x"3F3C57BB",
    x"3F3C5BFC",
    x"3F3C603E",
    x"3F3C647F",
    x"3F3C68C0",
    x"3F3C6D01",
    x"3F3C7141",
    x"3F3C7582",
    x"3F3C79C3",
    x"3F3C7E03",
    x"3F3C8244",
    x"3F3C8684",
    x"3F3C8AC4",
    x"3F3C8F04",
    x"3F3C9344",
    x"3F3C9784",
    x"3F3C9BC3",
    x"3F3CA003",
    x"3F3CA442",
    x"3F3CA881",
    x"3F3CACC1",
    x"3F3CB100",
    x"3F3CB53F",
    x"3F3CB97E",
    x"3F3CBDBC",
    x"3F3CC1FB",
    x"3F3CC63A",
    x"3F3CCA78",
    x"3F3CCEB6",
    x"3F3CD2F4",
    x"3F3CD733",
    x"3F3CDB70",
    x"3F3CDFAE",
    x"3F3CE3EC",
    x"3F3CE82A",
    x"3F3CEC67",
    x"3F3CF0A5",
    x"3F3CF4E2",
    x"3F3CF91F",
    x"3F3CFD5C",
    x"3F3D0199",
    x"3F3D05D6",
    x"3F3D0A12",
    x"3F3D0E4F",
    x"3F3D128C",
    x"3F3D16C8",
    x"3F3D1B04",
    x"3F3D1F40",
    x"3F3D237C",
    x"3F3D27B8",
    x"3F3D2BF4",
    x"3F3D3030",
    x"3F3D346B",
    x"3F3D38A7",
    x"3F3D3CE2",
    x"3F3D411D",
    x"3F3D4558",
    x"3F3D4993",
    x"3F3D4DCE",
    x"3F3D5209",
    x"3F3D5644",
    x"3F3D5A7E",
    x"3F3D5EB9",
    x"3F3D62F3",
    x"3F3D672D",
    x"3F3D6B67",
    x"3F3D6FA1",
    x"3F3D73DB",
    x"3F3D7815",
    x"3F3D7C4E",
    x"3F3D8088",
    x"3F3D84C1",
    x"3F3D88FB",
    x"3F3D8D34",
    x"3F3D916D",
    x"3F3D95A6",
    x"3F3D99DF",
    x"3F3D9E17",
    x"3F3DA250",
    x"3F3DA688",
    x"3F3DAAC1",
    x"3F3DAEF9",
    x"3F3DB331",
    x"3F3DB769",
    x"3F3DBBA1",
    x"3F3DBFD9",
    x"3F3DC411",
    x"3F3DC848",
    x"3F3DCC80",
    x"3F3DD0B7",
    x"3F3DD4EE",
    x"3F3DD925",
    x"3F3DDD5C",
    x"3F3DE193",
    x"3F3DE5CA",
    x"3F3DEA01",
    x"3F3DEE37",
    x"3F3DF26E",
    x"3F3DF6A4",
    x"3F3DFADA",
    x"3F3DFF10",
    x"3F3E0346",
    x"3F3E077C",
    x"3F3E0BB2",
    x"3F3E0FE7",
    x"3F3E141D",
    x"3F3E1852",
    x"3F3E1C88",
    x"3F3E20BD",
    x"3F3E24F2",
    x"3F3E2927",
    x"3F3E2D5C",
    x"3F3E3190",
    x"3F3E35C5",
    x"3F3E39F9",
    x"3F3E3E2E",
    x"3F3E4262",
    x"3F3E4696",
    x"3F3E4ACA",
    x"3F3E4EFE",
    x"3F3E5332",
    x"3F3E5766",
    x"3F3E5B99",
    x"3F3E5FCD",
    x"3F3E6400",
    x"3F3E6833",
    x"3F3E6C66",
    x"3F3E7099",
    x"3F3E74CC",
    x"3F3E78FF",
    x"3F3E7D31",
    x"3F3E8164",
    x"3F3E8596",
    x"3F3E89C9",
    x"3F3E8DFB",
    x"3F3E922D",
    x"3F3E965F",
    x"3F3E9A91",
    x"3F3E9EC3",
    x"3F3EA2F4",
    x"3F3EA726",
    x"3F3EAB57",
    x"3F3EAF88",
    x"3F3EB3B9",
    x"3F3EB7EA",
    x"3F3EBC1B",
    x"3F3EC04C",
    x"3F3EC47D",
    x"3F3EC8AD",
    x"3F3ECCDE",
    x"3F3ED10E",
    x"3F3ED53F",
    x"3F3ED96F",
    x"3F3EDD9F",
    x"3F3EE1CF",
    x"3F3EE5FE",
    x"3F3EEA2E",
    x"3F3EEE5E",
    x"3F3EF28D",
    x"3F3EF6BC",
    x"3F3EFAEB",
    x"3F3EFF1B",
    x"3F3F034A",
    x"3F3F0778",
    x"3F3F0BA7",
    x"3F3F0FD6",
    x"3F3F1404",
    x"3F3F1833",
    x"3F3F1C61",
    x"3F3F208F",
    x"3F3F24BD",
    x"3F3F28EB",
    x"3F3F2D19",
    x"3F3F3147",
    x"3F3F3574",
    x"3F3F39A2",
    x"3F3F3DCF",
    x"3F3F41FC",
    x"3F3F4629",
    x"3F3F4A56",
    x"3F3F4E83",
    x"3F3F52B0",
    x"3F3F56DD",
    x"3F3F5B09",
    x"3F3F5F36",
    x"3F3F6362",
    x"3F3F678E",
    x"3F3F6BBA",
    x"3F3F6FE6",
    x"3F3F7412",
    x"3F3F783E",
    x"3F3F7C6A",
    x"3F3F8095",
    x"3F3F84C0",
    x"3F3F88EC",
    x"3F3F8D17",
    x"3F3F9142",
    x"3F3F956D",
    x"3F3F9998",
    x"3F3F9DC2",
    x"3F3FA1ED",
    x"3F3FA617",
    x"3F3FAA42",
    x"3F3FAE6C",
    x"3F3FB296",
    x"3F3FB6C0",
    x"3F3FBAEA",
    x"3F3FBF14",
    x"3F3FC33E",
    x"3F3FC767",
    x"3F3FCB91",
    x"3F3FCFBA",
    x"3F3FD3E3",
    x"3F3FD80C",
    x"3F3FDC35",
    x"3F3FE05E",
    x"3F3FE487",
    x"3F3FE8AF",
    x"3F3FECD8",
    x"3F3FF100",
    x"3F3FF529",
    x"3F3FF951",
    x"3F3FFD79",
    x"3F4001A1",
    x"3F4005C8",
    x"3F4009F0",
    x"3F400E18",
    x"3F40123F",
    x"3F401667",
    x"3F401A8E",
    x"3F401EB5",
    x"3F4022DC",
    x"3F402703",
    x"3F402B2A",
    x"3F402F50",
    x"3F403377",
    x"3F40379D",
    x"3F403BC4",
    x"3F403FEA",
    x"3F404410",
    x"3F404836",
    x"3F404C5C",
    x"3F405081",
    x"3F4054A7",
    x"3F4058CD",
    x"3F405CF2",
    x"3F406117",
    x"3F40653C",
    x"3F406961",
    x"3F406D86",
    x"3F4071AB",
    x"3F4075D0",
    x"3F4079F4",
    x"3F407E19",
    x"3F40823D",
    x"3F408661",
    x"3F408A85",
    x"3F408EA9",
    x"3F4092CD",
    x"3F4096F1",
    x"3F409B15",
    x"3F409F38",
    x"3F40A35C",
    x"3F40A77F",
    x"3F40ABA2",
    x"3F40AFC5",
    x"3F40B3E8",
    x"3F40B80B",
    x"3F40BC2E",
    x"3F40C050",
    x"3F40C473",
    x"3F40C895",
    x"3F40CCB7",
    x"3F40D0DA",
    x"3F40D4FC",
    x"3F40D91E",
    x"3F40DD3F",
    x"3F40E161",
    x"3F40E583",
    x"3F40E9A4",
    x"3F40EDC5",
    x"3F40F1E7",
    x"3F40F608",
    x"3F40FA29",
    x"3F40FE49",
    x"3F41026A",
    x"3F41068B",
    x"3F410AAB",
    x"3F410ECC",
    x"3F4112EC",
    x"3F41170C",
    x"3F411B2C",
    x"3F411F4C",
    x"3F41236C",
    x"3F41278C",
    x"3F412BAB",
    x"3F412FCB",
    x"3F4133EA",
    x"3F413809",
    x"3F413C28",
    x"3F414047",
    x"3F414466",
    x"3F414885",
    x"3F414CA4",
    x"3F4150C2",
    x"3F4154E1",
    x"3F4158FF",
    x"3F415D1D",
    x"3F41613B",
    x"3F416559",
    x"3F416977",
    x"3F416D95",
    x"3F4171B2",
    x"3F4175D0",
    x"3F4179ED",
    x"3F417E0A",
    x"3F418228",
    x"3F418645",
    x"3F418A61",
    x"3F418E7E",
    x"3F41929B",
    x"3F4196B7",
    x"3F419AD4",
    x"3F419EF0",
    x"3F41A30C",
    x"3F41A728",
    x"3F41AB44",
    x"3F41AF60",
    x"3F41B37C",
    x"3F41B798",
    x"3F41BBB3",
    x"3F41BFCF",
    x"3F41C3EA",
    x"3F41C805",
    x"3F41CC20",
    x"3F41D03B",
    x"3F41D456",
    x"3F41D870",
    x"3F41DC8B",
    x"3F41E0A5",
    x"3F41E4C0",
    x"3F41E8DA",
    x"3F41ECF4",
    x"3F41F10E",
    x"3F41F528",
    x"3F41F942",
    x"3F41FD5B",
    x"3F420175",
    x"3F42058E",
    x"3F4209A7",
    x"3F420DC1",
    x"3F4211DA",
    x"3F4215F3",
    x"3F421A0B",
    x"3F421E24",
    x"3F42223D",
    x"3F422655",
    x"3F422A6E",
    x"3F422E86",
    x"3F42329E",
    x"3F4236B6",
    x"3F423ACE",
    x"3F423EE5",
    x"3F4242FD",
    x"3F424715",
    x"3F424B2C",
    x"3F424F43",
    x"3F42535B",
    x"3F425772",
    x"3F425B89",
    x"3F425F9F",
    x"3F4263B6",
    x"3F4267CD",
    x"3F426BE3",
    x"3F426FFA",
    x"3F427410",
    x"3F427826",
    x"3F427C3C",
    x"3F428052",
    x"3F428468",
    x"3F42887D",
    x"3F428C93",
    x"3F4290A8",
    x"3F4294BD",
    x"3F4298D3",
    x"3F429CE8",
    x"3F42A0FD",
    x"3F42A511",
    x"3F42A926",
    x"3F42AD3B",
    x"3F42B14F",
    x"3F42B564",
    x"3F42B978",
    x"3F42BD8C",
    x"3F42C1A0",
    x"3F42C5B4",
    x"3F42C9C8",
    x"3F42CDDB",
    x"3F42D1EF",
    x"3F42D602",
    x"3F42DA16",
    x"3F42DE29",
    x"3F42E23C",
    x"3F42E64F",
    x"3F42EA62",
    x"3F42EE74",
    x"3F42F287",
    x"3F42F69A",
    x"3F42FAAC",
    x"3F42FEBE",
    x"3F4302D0",
    x"3F4306E2",
    x"3F430AF4",
    x"3F430F06",
    x"3F431318",
    x"3F431729",
    x"3F431B3B",
    x"3F431F4C",
    x"3F43235D",
    x"3F43276E",
    x"3F432B7F",
    x"3F432F90",
    x"3F4333A1",
    x"3F4337B1",
    x"3F433BC2",
    x"3F433FD2",
    x"3F4343E2",
    x"3F4347F3",
    x"3F434C03",
    x"3F435012",
    x"3F435422",
    x"3F435832",
    x"3F435C41",
    x"3F436051",
    x"3F436460",
    x"3F43686F",
    x"3F436C7F",
    x"3F43708D",
    x"3F43749C",
    x"3F4378AB",
    x"3F437CBA",
    x"3F4380C8",
    x"3F4384D6",
    x"3F4388E5",
    x"3F438CF3",
    x"3F439101",
    x"3F43950F",
    x"3F43991D",
    x"3F439D2A",
    x"3F43A138",
    x"3F43A545",
    x"3F43A953",
    x"3F43AD60",
    x"3F43B16D",
    x"3F43B57A",
    x"3F43B987",
    x"3F43BD93",
    x"3F43C1A0",
    x"3F43C5AC",
    x"3F43C9B9",
    x"3F43CDC5",
    x"3F43D1D1",
    x"3F43D5DD",
    x"3F43D9E9",
    x"3F43DDF5",
    x"3F43E200",
    x"3F43E60C",
    x"3F43EA17",
    x"3F43EE23",
    x"3F43F22E",
    x"3F43F639",
    x"3F43FA44",
    x"3F43FE4F",
    x"3F44025A",
    x"3F440664",
    x"3F440A6F",
    x"3F440E79",
    x"3F441283",
    x"3F44168D",
    x"3F441A97",
    x"3F441EA1",
    x"3F4422AB",
    x"3F4426B5",
    x"3F442ABE",
    x"3F442EC8",
    x"3F4432D1",
    x"3F4436DA",
    x"3F443AE3",
    x"3F443EEC",
    x"3F4442F5",
    x"3F4446FE",
    x"3F444B06",
    x"3F444F0F",
    x"3F445317",
    x"3F44571F",
    x"3F445B27",
    x"3F445F2F",
    x"3F446337",
    x"3F44673F",
    x"3F446B47",
    x"3F446F4E",
    x"3F447356",
    x"3F44775D",
    x"3F447B64",
    x"3F447F6B",
    x"3F448372",
    x"3F448779",
    x"3F448B80",
    x"3F448F86",
    x"3F44938D",
    x"3F449793",
    x"3F449B99",
    x"3F449F9F",
    x"3F44A3A5",
    x"3F44A7AB",
    x"3F44ABB1",
    x"3F44AFB6",
    x"3F44B3BC",
    x"3F44B7C1",
    x"3F44BBC7",
    x"3F44BFCC",
    x"3F44C3D1",
    x"3F44C7D6",
    x"3F44CBDB",
    x"3F44CFDF",
    x"3F44D3E4",
    x"3F44D7E8",
    x"3F44DBED",
    x"3F44DFF1",
    x"3F44E3F5",
    x"3F44E7F9",
    x"3F44EBFD",
    x"3F44F000",
    x"3F44F404",
    x"3F44F807",
    x"3F44FC0B",
    x"3F45000E",
    x"3F450411",
    x"3F450814",
    x"3F450C17",
    x"3F45101A",
    x"3F45141D",
    x"3F45181F",
    x"3F451C22",
    x"3F452024",
    x"3F452426",
    x"3F452828",
    x"3F452C2A",
    x"3F45302C",
    x"3F45342E",
    x"3F45382F",
    x"3F453C31",
    x"3F454032",
    x"3F454433",
    x"3F454834",
    x"3F454C35",
    x"3F455036",
    x"3F455437",
    x"3F455838",
    x"3F455C38",
    x"3F456039",
    x"3F456439",
    x"3F456839",
    x"3F456C39",
    x"3F457039",
    x"3F457439",
    x"3F457839",
    x"3F457C38",
    x"3F458038",
    x"3F458437",
    x"3F458836",
    x"3F458C35",
    x"3F459034",
    x"3F459433",
    x"3F459832",
    x"3F459C31",
    x"3F45A02F",
    x"3F45A42D",
    x"3F45A82C",
    x"3F45AC2A",
    x"3F45B028",
    x"3F45B426",
    x"3F45B824",
    x"3F45BC21",
    x"3F45C01F",
    x"3F45C41C",
    x"3F45C819",
    x"3F45CC17",
    x"3F45D014",
    x"3F45D411",
    x"3F45D80E",
    x"3F45DC0A",
    x"3F45E007",
    x"3F45E403",
    x"3F45E800",
    x"3F45EBFC",
    x"3F45EFF8",
    x"3F45F3F4",
    x"3F45F7F0",
    x"3F45FBEC",
    x"3F45FFE7",
    x"3F4603E3",
    x"3F4607DE",
    x"3F460BDA",
    x"3F460FD5",
    x"3F4613D0",
    x"3F4617CB",
    x"3F461BC6",
    x"3F461FC0",
    x"3F4623BB",
    x"3F4627B5",
    x"3F462BB0",
    x"3F462FAA",
    x"3F4633A4",
    x"3F46379E",
    x"3F463B98",
    x"3F463F91",
    x"3F46438B",
    x"3F464785",
    x"3F464B7E",
    x"3F464F77",
    x"3F465370",
    x"3F465769",
    x"3F465B62",
    x"3F465F5B",
    x"3F466354",
    x"3F46674C",
    x"3F466B45",
    x"3F466F3D",
    x"3F467335",
    x"3F46772D",
    x"3F467B25",
    x"3F467F1D",
    x"3F468315",
    x"3F46870C",
    x"3F468B04",
    x"3F468EFB",
    x"3F4692F2",
    x"3F4696E9",
    x"3F469AE0",
    x"3F469ED7",
    x"3F46A2CE",
    x"3F46A6C5",
    x"3F46AABB",
    x"3F46AEB1",
    x"3F46B2A8",
    x"3F46B69E",
    x"3F46BA94",
    x"3F46BE8A",
    x"3F46C280",
    x"3F46C675",
    x"3F46CA6B",
    x"3F46CE60",
    x"3F46D256",
    x"3F46D64B",
    x"3F46DA40",
    x"3F46DE35",
    x"3F46E22A",
    x"3F46E61E",
    x"3F46EA13",
    x"3F46EE07",
    x"3F46F1FC",
    x"3F46F5F0",
    x"3F46F9E4",
    x"3F46FDD8",
    x"3F4701CC",
    x"3F4705C0",
    x"3F4709B3",
    x"3F470DA7",
    x"3F47119A",
    x"3F47158D",
    x"3F471981",
    x"3F471D74",
    x"3F472167",
    x"3F472559",
    x"3F47294C",
    x"3F472D3F",
    x"3F473131",
    x"3F473523",
    x"3F473916",
    x"3F473D08",
    x"3F4740FA",
    x"3F4744EB",
    x"3F4748DD",
    x"3F474CCF",
    x"3F4750C0",
    x"3F4754B2",
    x"3F4758A3",
    x"3F475C94",
    x"3F476085",
    x"3F476476",
    x"3F476866",
    x"3F476C57",
    x"3F477048",
    x"3F477438",
    x"3F477828",
    x"3F477C18",
    x"3F478008",
    x"3F4783F8",
    x"3F4787E8",
    x"3F478BD8",
    x"3F478FC7",
    x"3F4793B7",
    x"3F4797A6",
    x"3F479B95",
    x"3F479F84",
    x"3F47A373",
    x"3F47A762",
    x"3F47AB51",
    x"3F47AF3F",
    x"3F47B32E",
    x"3F47B71C",
    x"3F47BB0A",
    x"3F47BEF9",
    x"3F47C2E7",
    x"3F47C6D4",
    x"3F47CAC2",
    x"3F47CEB0",
    x"3F47D29D",
    x"3F47D68B",
    x"3F47DA78",
    x"3F47DE65",
    x"3F47E252",
    x"3F47E63F",
    x"3F47EA2C",
    x"3F47EE18",
    x"3F47F205",
    x"3F47F5F1",
    x"3F47F9DE",
    x"3F47FDCA",
    x"3F4801B6",
    x"3F4805A2",
    x"3F48098E",
    x"3F480D79",
    x"3F481165",
    x"3F481550",
    x"3F48193C",
    x"3F481D27",
    x"3F482112",
    x"3F4824FD",
    x"3F4828E8",
    x"3F482CD3",
    x"3F4830BD",
    x"3F4834A8",
    x"3F483892",
    x"3F483C7C",
    x"3F484067",
    x"3F484451",
    x"3F48483A",
    x"3F484C24",
    x"3F48500E",
    x"3F4853F7",
    x"3F4857E1",
    x"3F485BCA",
    x"3F485FB3",
    x"3F48639C",
    x"3F486785",
    x"3F486B6E",
    x"3F486F57",
    x"3F48733F",
    x"3F487728",
    x"3F487B10",
    x"3F487EF8",
    x"3F4882E0",
    x"3F4886C8",
    x"3F488AB0",
    x"3F488E98",
    x"3F48927F",
    x"3F489667",
    x"3F489A4E",
    x"3F489E36",
    x"3F48A21D",
    x"3F48A604",
    x"3F48A9EA",
    x"3F48ADD1",
    x"3F48B1B8",
    x"3F48B59E",
    x"3F48B985",
    x"3F48BD6B",
    x"3F48C151",
    x"3F48C537",
    x"3F48C91D",
    x"3F48CD03",
    x"3F48D0E9",
    x"3F48D4CE",
    x"3F48D8B3",
    x"3F48DC99",
    x"3F48E07E",
    x"3F48E463",
    x"3F48E848",
    x"3F48EC2D",
    x"3F48F011",
    x"3F48F3F6",
    x"3F48F7DA",
    x"3F48FBBF",
    x"3F48FFA3",
    x"3F490387",
    x"3F49076B",
    x"3F490B4F",
    x"3F490F33",
    x"3F491316",
    x"3F4916FA",
    x"3F491ADD",
    x"3F491EC0",
    x"3F4922A3",
    x"3F492686",
    x"3F492A69",
    x"3F492E4C",
    x"3F49322F",
    x"3F493611",
    x"3F4939F4",
    x"3F493DD6",
    x"3F4941B8",
    x"3F49459A",
    x"3F49497C",
    x"3F494D5E",
    x"3F49513F",
    x"3F495521",
    x"3F495902",
    x"3F495CE4",
    x"3F4960C5",
    x"3F4964A6",
    x"3F496887",
    x"3F496C68",
    x"3F497048",
    x"3F497429",
    x"3F497809",
    x"3F497BEA",
    x"3F497FCA",
    x"3F4983AA",
    x"3F49878A",
    x"3F498B6A",
    x"3F498F4A",
    x"3F499329",
    x"3F499709",
    x"3F499AE8",
    x"3F499EC7",
    x"3F49A2A6",
    x"3F49A685",
    x"3F49AA64",
    x"3F49AE43",
    x"3F49B222",
    x"3F49B600",
    x"3F49B9DF",
    x"3F49BDBD",
    x"3F49C19B",
    x"3F49C579",
    x"3F49C957",
    x"3F49CD35",
    x"3F49D112",
    x"3F49D4F0",
    x"3F49D8CD",
    x"3F49DCAB",
    x"3F49E088",
    x"3F49E465",
    x"3F49E842",
    x"3F49EC1F",
    x"3F49EFFB",
    x"3F49F3D8",
    x"3F49F7B4",
    x"3F49FB91",
    x"3F49FF6D",
    x"3F4A0349",
    x"3F4A0725",
    x"3F4A0B01",
    x"3F4A0EDC",
    x"3F4A12B8",
    x"3F4A1693",
    x"3F4A1A6F",
    x"3F4A1E4A",
    x"3F4A2225",
    x"3F4A2600",
    x"3F4A29DB",
    x"3F4A2DB6",
    x"3F4A3190",
    x"3F4A356B",
    x"3F4A3945",
    x"3F4A3D1F",
    x"3F4A40F9",
    x"3F4A44D3",
    x"3F4A48AD",
    x"3F4A4C87",
    x"3F4A5061",
    x"3F4A543A",
    x"3F4A5814",
    x"3F4A5BED",
    x"3F4A5FC6",
    x"3F4A639F",
    x"3F4A6778",
    x"3F4A6B51",
    x"3F4A6F29",
    x"3F4A7302",
    x"3F4A76DA",
    x"3F4A7AB3",
    x"3F4A7E8B",
    x"3F4A8263",
    x"3F4A863B",
    x"3F4A8A13",
    x"3F4A8DEA",
    x"3F4A91C2",
    x"3F4A9599",
    x"3F4A9971",
    x"3F4A9D48",
    x"3F4AA11F",
    x"3F4AA4F6",
    x"3F4AA8CD",
    x"3F4AACA4",
    x"3F4AB07A",
    x"3F4AB451",
    x"3F4AB827",
    x"3F4ABBFD",
    x"3F4ABFD3",
    x"3F4AC3A9",
    x"3F4AC77F",
    x"3F4ACB55",
    x"3F4ACF2A",
    x"3F4AD300",
    x"3F4AD6D5",
    x"3F4ADAAB",
    x"3F4ADE80",
    x"3F4AE255",
    x"3F4AE62A",
    x"3F4AE9FE",
    x"3F4AEDD3",
    x"3F4AF1A8",
    x"3F4AF57C",
    x"3F4AF950",
    x"3F4AFD24",
    x"3F4B00F8",
    x"3F4B04CC",
    x"3F4B08A0",
    x"3F4B0C74",
    x"3F4B1047",
    x"3F4B141B",
    x"3F4B17EE",
    x"3F4B1BC1",
    x"3F4B1F94",
    x"3F4B2367",
    x"3F4B273A",
    x"3F4B2B0D",
    x"3F4B2EDF",
    x"3F4B32B2",
    x"3F4B3684",
    x"3F4B3A56",
    x"3F4B3E28",
    x"3F4B41FA",
    x"3F4B45CC",
    x"3F4B499E",
    x"3F4B4D6F",
    x"3F4B5141",
    x"3F4B5512",
    x"3F4B58E3",
    x"3F4B5CB4",
    x"3F4B6085",
    x"3F4B6456",
    x"3F4B6827",
    x"3F4B6BF7",
    x"3F4B6FC8",
    x"3F4B7398",
    x"3F4B7768",
    x"3F4B7B39",
    x"3F4B7F09",
    x"3F4B82D8",
    x"3F4B86A8",
    x"3F4B8A78",
    x"3F4B8E47",
    x"3F4B9217",
    x"3F4B95E6",
    x"3F4B99B5",
    x"3F4B9D84",
    x"3F4BA153",
    x"3F4BA522",
    x"3F4BA8F0",
    x"3F4BACBF",
    x"3F4BB08D",
    x"3F4BB45B",
    x"3F4BB82A",
    x"3F4BBBF8",
    x"3F4BBFC6",
    x"3F4BC393",
    x"3F4BC761",
    x"3F4BCB2F",
    x"3F4BCEFC",
    x"3F4BD2C9",
    x"3F4BD696",
    x"3F4BDA63",
    x"3F4BDE30",
    x"3F4BE1FD",
    x"3F4BE5CA",
    x"3F4BE996",
    x"3F4BED63",
    x"3F4BF12F",
    x"3F4BF4FB",
    x"3F4BF8C7",
    x"3F4BFC93",
    x"3F4C005F",
    x"3F4C042B",
    x"3F4C07F6",
    x"3F4C0BC2",
    x"3F4C0F8D",
    x"3F4C1358",
    x"3F4C1723",
    x"3F4C1AEE",
    x"3F4C1EB9",
    x"3F4C2284",
    x"3F4C264E",
    x"3F4C2A19",
    x"3F4C2DE3",
    x"3F4C31AD",
    x"3F4C3578",
    x"3F4C3942",
    x"3F4C3D0B",
    x"3F4C40D5",
    x"3F4C449F",
    x"3F4C4868",
    x"3F4C4C32",
    x"3F4C4FFB",
    x"3F4C53C4",
    x"3F4C578D",
    x"3F4C5B56",
    x"3F4C5F1E",
    x"3F4C62E7",
    x"3F4C66B0",
    x"3F4C6A78",
    x"3F4C6E40",
    x"3F4C7208",
    x"3F4C75D0",
    x"3F4C7998",
    x"3F4C7D60",
    x"3F4C8128",
    x"3F4C84EF",
    x"3F4C88B6",
    x"3F4C8C7E",
    x"3F4C9045",
    x"3F4C940C",
    x"3F4C97D3",
    x"3F4C9B99",
    x"3F4C9F60",
    x"3F4CA327",
    x"3F4CA6ED",
    x"3F4CAAB3",
    x"3F4CAE79",
    x"3F4CB23F",
    x"3F4CB605",
    x"3F4CB9CB",
    x"3F4CBD91",
    x"3F4CC156",
    x"3F4CC51C",
    x"3F4CC8E1",
    x"3F4CCCA6",
    x"3F4CD06B",
    x"3F4CD430",
    x"3F4CD7F5",
    x"3F4CDBBA",
    x"3F4CDF7E",
    x"3F4CE343",
    x"3F4CE707",
    x"3F4CEACB",
    x"3F4CEE8F",
    x"3F4CF253",
    x"3F4CF617",
    x"3F4CF9DB",
    x"3F4CFD9E",
    x"3F4D0162",
    x"3F4D0525",
    x"3F4D08E8",
    x"3F4D0CAB",
    x"3F4D106E",
    x"3F4D1431",
    x"3F4D17F4",
    x"3F4D1BB6",
    x"3F4D1F79",
    x"3F4D233B",
    x"3F4D26FD",
    x"3F4D2ABF",
    x"3F4D2E81",
    x"3F4D3243",
    x"3F4D3605",
    x"3F4D39C6",
    x"3F4D3D88",
    x"3F4D4149",
    x"3F4D450A",
    x"3F4D48CB",
    x"3F4D4C8C",
    x"3F4D504D",
    x"3F4D540E",
    x"3F4D57CE",
    x"3F4D5B8F",
    x"3F4D5F4F",
    x"3F4D6310",
    x"3F4D66D0",
    x"3F4D6A90",
    x"3F4D6E4F",
    x"3F4D720F",
    x"3F4D75CF",
    x"3F4D798E",
    x"3F4D7D4E",
    x"3F4D810D",
    x"3F4D84CC",
    x"3F4D888B",
    x"3F4D8C4A",
    x"3F4D9009",
    x"3F4D93C7",
    x"3F4D9786",
    x"3F4D9B44",
    x"3F4D9F02",
    x"3F4DA2C0",
    x"3F4DA67E",
    x"3F4DAA3C",
    x"3F4DADFA",
    x"3F4DB1B8",
    x"3F4DB575",
    x"3F4DB932",
    x"3F4DBCF0",
    x"3F4DC0AD",
    x"3F4DC46A",
    x"3F4DC827",
    x"3F4DCBE3",
    x"3F4DCFA0",
    x"3F4DD35D",
    x"3F4DD719",
    x"3F4DDAD5",
    x"3F4DDE91",
    x"3F4DE24D",
    x"3F4DE609",
    x"3F4DE9C5",
    x"3F4DED81",
    x"3F4DF13C",
    x"3F4DF4F8",
    x"3F4DF8B3",
    x"3F4DFC6E",
    x"3F4E0029",
    x"3F4E03E4",
    x"3F4E079F",
    x"3F4E0B59",
    x"3F4E0F14",
    x"3F4E12CE",
    x"3F4E1689",
    x"3F4E1A43",
    x"3F4E1DFD",
    x"3F4E21B7",
    x"3F4E2570",
    x"3F4E292A",
    x"3F4E2CE4",
    x"3F4E309D",
    x"3F4E3456",
    x"3F4E380F",
    x"3F4E3BC8",
    x"3F4E3F81",
    x"3F4E433A",
    x"3F4E46F3",
    x"3F4E4AAB",
    x"3F4E4E64",
    x"3F4E521C",
    x"3F4E55D4",
    x"3F4E598C",
    x"3F4E5D44",
    x"3F4E60FC",
    x"3F4E64B4",
    x"3F4E686B",
    x"3F4E6C23",
    x"3F4E6FDA",
    x"3F4E7391",
    x"3F4E7748",
    x"3F4E7AFF",
    x"3F4E7EB6",
    x"3F4E826C",
    x"3F4E8623",
    x"3F4E89D9",
    x"3F4E8D90",
    x"3F4E9146",
    x"3F4E94FC",
    x"3F4E98B2",
    x"3F4E9C68",
    x"3F4EA01D",
    x"3F4EA3D3",
    x"3F4EA788",
    x"3F4EAB3E",
    x"3F4EAEF3",
    x"3F4EB2A8",
    x"3F4EB65D",
    x"3F4EBA12",
    x"3F4EBDC6",
    x"3F4EC17B",
    x"3F4EC52F",
    x"3F4EC8E4",
    x"3F4ECC98",
    x"3F4ED04C",
    x"3F4ED400",
    x"3F4ED7B3",
    x"3F4EDB67",
    x"3F4EDF1B",
    x"3F4EE2CE",
    x"3F4EE681",
    x"3F4EEA35",
    x"3F4EEDE8",
    x"3F4EF19B",
    x"3F4EF54D",
    x"3F4EF900",
    x"3F4EFCB3",
    x"3F4F0065",
    x"3F4F0417",
    x"3F4F07CA",
    x"3F4F0B7C",
    x"3F4F0F2E",
    x"3F4F12DF",
    x"3F4F1691",
    x"3F4F1A43",
    x"3F4F1DF4",
    x"3F4F21A5",
    x"3F4F2557",
    x"3F4F2908",
    x"3F4F2CB9",
    x"3F4F3069",
    x"3F4F341A",
    x"3F4F37CB",
    x"3F4F3B7B",
    x"3F4F3F2B",
    x"3F4F42DC",
    x"3F4F468C",
    x"3F4F4A3C",
    x"3F4F4DEB",
    x"3F4F519B",
    x"3F4F554B",
    x"3F4F58FA",
    x"3F4F5CA9",
    x"3F4F6059",
    x"3F4F6408",
    x"3F4F67B7",
    x"3F4F6B65",
    x"3F4F6F14",
    x"3F4F72C3",
    x"3F4F7671",
    x"3F4F7A1F",
    x"3F4F7DCE",
    x"3F4F817C",
    x"3F4F852A",
    x"3F4F88D7",
    x"3F4F8C85",
    x"3F4F9033",
    x"3F4F93E0",
    x"3F4F978D",
    x"3F4F9B3B",
    x"3F4F9EE8",
    x"3F4FA295",
    x"3F4FA642",
    x"3F4FA9EE",
    x"3F4FAD9B",
    x"3F4FB147",
    x"3F4FB4F4",
    x"3F4FB8A0",
    x"3F4FBC4C",
    x"3F4FBFF8",
    x"3F4FC3A4",
    x"3F4FC74F",
    x"3F4FCAFB",
    x"3F4FCEA6",
    x"3F4FD252",
    x"3F4FD5FD",
    x"3F4FD9A8",
    x"3F4FDD53",
    x"3F4FE0FE",
    x"3F4FE4A8",
    x"3F4FE853",
    x"3F4FEBFD",
    x"3F4FEFA8",
    x"3F4FF352",
    x"3F4FF6FC",
    x"3F4FFAA6",
    x"3F4FFE50",
    x"3F5001F9",
    x"3F5005A3",
    x"3F50094C",
    x"3F500CF6",
    x"3F50109F",
    x"3F501448",
    x"3F5017F1",
    x"3F501B9A",
    x"3F501F42",
    x"3F5022EB",
    x"3F502693",
    x"3F502A3B",
    x"3F502DE4",
    x"3F50318C",
    x"3F503534",
    x"3F5038DB",
    x"3F503C83",
    x"3F50402B",
    x"3F5043D2",
    x"3F504779",
    x"3F504B21",
    x"3F504EC8",
    x"3F50526F",
    x"3F505615",
    x"3F5059BC",
    x"3F505D63",
    x"3F506109",
    x"3F5064AF",
    x"3F506856",
    x"3F506BFC",
    x"3F506FA1",
    x"3F507347",
    x"3F5076ED",
    x"3F507A92",
    x"3F507E38",
    x"3F5081DD",
    x"3F508582",
    x"3F508927",
    x"3F508CCC",
    x"3F509071",
    x"3F509416",
    x"3F5097BA",
    x"3F509B5F",
    x"3F509F03",
    x"3F50A2A7",
    x"3F50A64B",
    x"3F50A9EF",
    x"3F50AD93",
    x"3F50B137",
    x"3F50B4DA",
    x"3F50B87E",
    x"3F50BC21",
    x"3F50BFC4",
    x"3F50C367",
    x"3F50C70A",
    x"3F50CAAD",
    x"3F50CE4F",
    x"3F50D1F2",
    x"3F50D594",
    x"3F50D937",
    x"3F50DCD9",
    x"3F50E07B",
    x"3F50E41D",
    x"3F50E7BE",
    x"3F50EB60",
    x"3F50EF02",
    x"3F50F2A3",
    x"3F50F644",
    x"3F50F9E5",
    x"3F50FD86",
    x"3F510127",
    x"3F5104C8",
    x"3F510869",
    x"3F510C09",
    x"3F510FAA",
    x"3F51134A",
    x"3F5116EA",
    x"3F511A8A",
    x"3F511E2A",
    x"3F5121CA",
    x"3F512569",
    x"3F512909",
    x"3F512CA8",
    x"3F513047",
    x"3F5133E7",
    x"3F513786",
    x"3F513B25",
    x"3F513EC3",
    x"3F514262",
    x"3F514600",
    x"3F51499F",
    x"3F514D3D",
    x"3F5150DB",
    x"3F515479",
    x"3F515817",
    x"3F515BB5",
    x"3F515F52",
    x"3F5162F0",
    x"3F51668D",
    x"3F516A2A",
    x"3F516DC8",
    x"3F517165",
    x"3F517501",
    x"3F51789E",
    x"3F517C3B",
    x"3F517FD7",
    x"3F518374",
    x"3F518710",
    x"3F518AAC",
    x"3F518E48",
    x"3F5191E4",
    x"3F51957F",
    x"3F51991B",
    x"3F519CB7",
    x"3F51A052",
    x"3F51A3ED",
    x"3F51A788",
    x"3F51AB23",
    x"3F51AEBE",
    x"3F51B259",
    x"3F51B5F3",
    x"3F51B98E",
    x"3F51BD28",
    x"3F51C0C2",
    x"3F51C45C",
    x"3F51C7F6",
    x"3F51CB90",
    x"3F51CF2A",
    x"3F51D2C3",
    x"3F51D65D",
    x"3F51D9F6",
    x"3F51DD8F",
    x"3F51E129",
    x"3F51E4C1",
    x"3F51E85A",
    x"3F51EBF3",
    x"3F51EF8C",
    x"3F51F324",
    x"3F51F6BC",
    x"3F51FA54",
    x"3F51FDED",
    x"3F520184",
    x"3F52051C",
    x"3F5208B4",
    x"3F520C4C",
    x"3F520FE3",
    x"3F52137A",
    x"3F521711",
    x"3F521AA8",
    x"3F521E3F",
    x"3F5221D6",
    x"3F52256D",
    x"3F522903",
    x"3F522C9A",
    x"3F523030",
    x"3F5233C6",
    x"3F52375C",
    x"3F523AF2",
    x"3F523E88",
    x"3F52421E",
    x"3F5245B3",
    x"3F524949",
    x"3F524CDE",
    x"3F525073",
    x"3F525408",
    x"3F52579D",
    x"3F525B32",
    x"3F525EC6",
    x"3F52625B",
    x"3F5265EF",
    x"3F526983",
    x"3F526D18",
    x"3F5270AC",
    x"3F52743F",
    x"3F5277D3",
    x"3F527B67",
    x"3F527EFA",
    x"3F52828E",
    x"3F528621",
    x"3F5289B4",
    x"3F528D47",
    x"3F5290DA",
    x"3F52946D",
    x"3F5297FF",
    x"3F529B92",
    x"3F529F24",
    x"3F52A2B6",
    x"3F52A649",
    x"3F52A9DA",
    x"3F52AD6C",
    x"3F52B0FE",
    x"3F52B490",
    x"3F52B821",
    x"3F52BBB2",
    x"3F52BF44",
    x"3F52C2D5",
    x"3F52C666",
    x"3F52C9F7",
    x"3F52CD87",
    x"3F52D118",
    x"3F52D4A8",
    x"3F52D839",
    x"3F52DBC9",
    x"3F52DF59",
    x"3F52E2E9",
    x"3F52E679",
    x"3F52EA08",
    x"3F52ED98",
    x"3F52F127",
    x"3F52F4B7",
    x"3F52F846",
    x"3F52FBD5",
    x"3F52FF64",
    x"3F5302F3",
    x"3F530681",
    x"3F530A10",
    x"3F530D9E",
    x"3F53112D",
    x"3F5314BB",
    x"3F531849",
    x"3F531BD7",
    x"3F531F65",
    x"3F5322F2",
    x"3F532680",
    x"3F532A0D",
    x"3F532D9A",
    x"3F533128",
    x"3F5334B5",
    x"3F533841",
    x"3F533BCE",
    x"3F533F5B",
    x"3F5342E7",
    x"3F534674",
    x"3F534A00",
    x"3F534D8C",
    x"3F535118",
    x"3F5354A4",
    x"3F535830",
    x"3F535BBB",
    x"3F535F47",
    x"3F5362D2",
    x"3F53665E",
    x"3F5369E9",
    x"3F536D74",
    x"3F5370FF",
    x"3F537489",
    x"3F537814",
    x"3F537B9E",
    x"3F537F29",
    x"3F5382B3",
    x"3F53863D",
    x"3F5389C7",
    x"3F538D51",
    x"3F5390DB",
    x"3F539464",
    x"3F5397EE",
    x"3F539B77",
    x"3F539F00",
    x"3F53A289",
    x"3F53A612",
    x"3F53A99B",
    x"3F53AD24",
    x"3F53B0AC",
    x"3F53B435",
    x"3F53B7BD",
    x"3F53BB45",
    x"3F53BECD",
    x"3F53C255",
    x"3F53C5DD",
    x"3F53C965",
    x"3F53CCEC",
    x"3F53D074",
    x"3F53D3FB",
    x"3F53D782",
    x"3F53DB09",
    x"3F53DE90",
    x"3F53E217",
    x"3F53E59D",
    x"3F53E924",
    x"3F53ECAA",
    x"3F53F031",
    x"3F53F3B7",
    x"3F53F73D",
    x"3F53FAC3",
    x"3F53FE48",
    x"3F5401CE",
    x"3F540553",
    x"3F5408D9",
    x"3F540C5E",
    x"3F540FE3",
    x"3F541368",
    x"3F5416ED",
    x"3F541A72",
    x"3F541DF6",
    x"3F54217B",
    x"3F5424FF",
    x"3F542883",
    x"3F542C08",
    x"3F542F8C",
    x"3F54330F",
    x"3F543693",
    x"3F543A17",
    x"3F543D9A",
    x"3F54411D",
    x"3F5444A1",
    x"3F544824",
    x"3F544BA7",
    x"3F544F2A",
    x"3F5452AC",
    x"3F54562F",
    x"3F5459B1",
    x"3F545D33",
    x"3F5460B6",
    x"3F546438",
    x"3F5467BA",
    x"3F546B3B",
    x"3F546EBD",
    x"3F54723F",
    x"3F5475C0",
    x"3F547941",
    x"3F547CC3",
    x"3F548044",
    x"3F5483C4",
    x"3F548745",
    x"3F548AC6",
    x"3F548E46",
    x"3F5491C7",
    x"3F549547",
    x"3F5498C7",
    x"3F549C47",
    x"3F549FC7",
    x"3F54A347",
    x"3F54A6C6",
    x"3F54AA46",
    x"3F54ADC5",
    x"3F54B144",
    x"3F54B4C4",
    x"3F54B843",
    x"3F54BBC1",
    x"3F54BF40",
    x"3F54C2BF",
    x"3F54C63D",
    x"3F54C9BC",
    x"3F54CD3A",
    x"3F54D0B8",
    x"3F54D436",
    x"3F54D7B4",
    x"3F54DB31",
    x"3F54DEAF",
    x"3F54E22C",
    x"3F54E5AA",
    x"3F54E927",
    x"3F54ECA4",
    x"3F54F021",
    x"3F54F39E",
    x"3F54F71A",
    x"3F54FA97",
    x"3F54FE13",
    x"3F55018F",
    x"3F55050C",
    x"3F550888",
    x"3F550C04",
    x"3F550F7F",
    x"3F5512FB",
    x"3F551676",
    x"3F5519F2",
    x"3F551D6D",
    x"3F5520E8",
    x"3F552463",
    x"3F5527DE",
    x"3F552B59",
    x"3F552ED4",
    x"3F55324E",
    x"3F5535C8",
    x"3F553943",
    x"3F553CBD",
    x"3F554037",
    x"3F5543B1",
    x"3F55472A",
    x"3F554AA4",
    x"3F554E1D",
    x"3F555197",
    x"3F555510",
    x"3F555889",
    x"3F555C02",
    x"3F555F7B",
    x"3F5562F3",
    x"3F55666C",
    x"3F5569E4",
    x"3F556D5D",
    x"3F5570D5",
    x"3F55744D",
    x"3F5577C5",
    x"3F557B3D",
    x"3F557EB4",
    x"3F55822C",
    x"3F5585A3",
    x"3F55891A",
    x"3F558C92",
    x"3F559009",
    x"3F55937F",
    x"3F5596F6",
    x"3F559A6D",
    x"3F559DE3",
    x"3F55A15A",
    x"3F55A4D0",
    x"3F55A846",
    x"3F55ABBC",
    x"3F55AF32",
    x"3F55B2A8",
    x"3F55B61D",
    x"3F55B993",
    x"3F55BD08",
    x"3F55C07D",
    x"3F55C3F2",
    x"3F55C767",
    x"3F55CADC",
    x"3F55CE51",
    x"3F55D1C5",
    x"3F55D53A",
    x"3F55D8AE",
    x"3F55DC22",
    x"3F55DF96",
    x"3F55E30A",
    x"3F55E67E",
    x"3F55E9F2",
    x"3F55ED65",
    x"3F55F0D9",
    x"3F55F44C",
    x"3F55F7BF",
    x"3F55FB32",
    x"3F55FEA5",
    x"3F560218",
    x"3F56058B",
    x"3F5608FD",
    x"3F560C70",
    x"3F560FE2",
    x"3F561354",
    x"3F5616C6",
    x"3F561A38",
    x"3F561DA9",
    x"3F56211B",
    x"3F56248D",
    x"3F5627FE",
    x"3F562B6F",
    x"3F562EE0",
    x"3F563251",
    x"3F5635C2",
    x"3F563933",
    x"3F563CA3",
    x"3F564014",
    x"3F564384",
    x"3F5646F4",
    x"3F564A64",
    x"3F564DD4",
    x"3F565144",
    x"3F5654B4",
    x"3F565823",
    x"3F565B93",
    x"3F565F02",
    x"3F566271",
    x"3F5665E0",
    x"3F56694F",
    x"3F566CBE",
    x"3F56702C",
    x"3F56739B",
    x"3F567709",
    x"3F567A78",
    x"3F567DE6",
    x"3F568154",
    x"3F5684C2",
    x"3F56882F",
    x"3F568B9D",
    x"3F568F0A",
    x"3F569278",
    x"3F5695E5",
    x"3F569952",
    x"3F569CBF",
    x"3F56A02C",
    x"3F56A399",
    x"3F56A705",
    x"3F56AA72",
    x"3F56ADDE",
    x"3F56B14A",
    x"3F56B4B6",
    x"3F56B822",
    x"3F56BB8E",
    x"3F56BEF9",
    x"3F56C265",
    x"3F56C5D0",
    x"3F56C93C",
    x"3F56CCA7",
    x"3F56D012",
    x"3F56D37D",
    x"3F56D6E8",
    x"3F56DA52",
    x"3F56DDBD",
    x"3F56E127",
    x"3F56E491",
    x"3F56E7FB",
    x"3F56EB65",
    x"3F56EECF",
    x"3F56F239",
    x"3F56F5A3",
    x"3F56F90C",
    x"3F56FC75",
    x"3F56FFDF",
    x"3F570348",
    x"3F5706B1",
    x"3F570A19",
    x"3F570D82",
    x"3F5710EB",
    x"3F571453",
    x"3F5717BB",
    x"3F571B24",
    x"3F571E8C",
    x"3F5721F3",
    x"3F57255B",
    x"3F5728C3",
    x"3F572C2A",
    x"3F572F92",
    x"3F5732F9",
    x"3F573660",
    x"3F5739C7",
    x"3F573D2E",
    x"3F574095",
    x"3F5743FB",
    x"3F574762",
    x"3F574AC8",
    x"3F574E2F",
    x"3F575195",
    x"3F5754FB",
    x"3F575860",
    x"3F575BC6",
    x"3F575F2C",
    x"3F576291",
    x"3F5765F6",
    x"3F57695C",
    x"3F576CC1",
    x"3F577026",
    x"3F57738A",
    x"3F5776EF",
    x"3F577A54",
    x"3F577DB8",
    x"3F57811C",
    x"3F578480",
    x"3F5787E4",
    x"3F578B48",
    x"3F578EAC",
    x"3F579210",
    x"3F579573",
    x"3F5798D7",
    x"3F579C3A",
    x"3F579F9D",
    x"3F57A300",
    x"3F57A663",
    x"3F57A9C6",
    x"3F57AD28",
    x"3F57B08B",
    x"3F57B3ED",
    x"3F57B74F",
    x"3F57BAB1",
    x"3F57BE13",
    x"3F57C175",
    x"3F57C4D7",
    x"3F57C838",
    x"3F57CB9A",
    x"3F57CEFB",
    x"3F57D25C",
    x"3F57D5BD",
    x"3F57D91E",
    x"3F57DC7F",
    x"3F57DFDF",
    x"3F57E340",
    x"3F57E6A0",
    x"3F57EA01",
    x"3F57ED61",
    x"3F57F0C1",
    x"3F57F421",
    x"3F57F780",
    x"3F57FAE0",
    x"3F57FE3F",
    x"3F58019F",
    x"3F5804FE",
    x"3F58085D",
    x"3F580BBC",
    x"3F580F1B",
    x"3F581279",
    x"3F5815D8",
    x"3F581936",
    x"3F581C95",
    x"3F581FF3",
    x"3F582351",
    x"3F5826AF",
    x"3F582A0D",
    x"3F582D6A",
    x"3F5830C8",
    x"3F583425",
    x"3F583782",
    x"3F583AE0",
    x"3F583E3D",
    x"3F584199",
    x"3F5844F6",
    x"3F584853",
    x"3F584BAF",
    x"3F584F0C",
    x"3F585268",
    x"3F5855C4",
    x"3F585920",
    x"3F585C7C",
    x"3F585FD7",
    x"3F586333",
    x"3F58668E",
    x"3F5869EA",
    x"3F586D45",
    x"3F5870A0",
    x"3F5873FB",
    x"3F587756",
    x"3F587AB0",
    x"3F587E0B",
    x"3F588165",
    x"3F5884BF",
    x"3F58881A",
    x"3F588B74",
    x"3F588ECD",
    x"3F589227",
    x"3F589581",
    x"3F5898DA",
    x"3F589C34",
    x"3F589F8D",
    x"3F58A2E6",
    x"3F58A63F",
    x"3F58A998",
    x"3F58ACF0",
    x"3F58B049",
    x"3F58B3A1",
    x"3F58B6FA",
    x"3F58BA52",
    x"3F58BDAA",
    x"3F58C102",
    x"3F58C45A",
    x"3F58C7B1",
    x"3F58CB09",
    x"3F58CE60",
    x"3F58D1B7",
    x"3F58D50E",
    x"3F58D865",
    x"3F58DBBC",
    x"3F58DF13",
    x"3F58E26A",
    x"3F58E5C0",
    x"3F58E916",
    x"3F58EC6D",
    x"3F58EFC3",
    x"3F58F319",
    x"3F58F66F",
    x"3F58F9C4",
    x"3F58FD1A",
    x"3F59006F",
    x"3F5903C5",
    x"3F59071A",
    x"3F590A6F",
    x"3F590DC4",
    x"3F591118",
    x"3F59146D",
    x"3F5917C2",
    x"3F591B16",
    x"3F591E6A",
    x"3F5921BE",
    x"3F592512",
    x"3F592866",
    x"3F592BBA",
    x"3F592F0E",
    x"3F593261",
    x"3F5935B4",
    x"3F593908",
    x"3F593C5B",
    x"3F593FAE",
    x"3F594300",
    x"3F594653",
    x"3F5949A6",
    x"3F594CF8",
    x"3F59504A",
    x"3F59539C",
    x"3F5956EE",
    x"3F595A40",
    x"3F595D92",
    x"3F5960E4",
    x"3F596435",
    x"3F596787",
    x"3F596AD8",
    x"3F596E29",
    x"3F59717A",
    x"3F5974CB",
    x"3F59781C",
    x"3F597B6C",
    x"3F597EBD",
    x"3F59820D",
    x"3F59855D",
    x"3F5988AD",
    x"3F598BFD",
    x"3F598F4D",
    x"3F59929D",
    x"3F5995EC",
    x"3F59993C",
    x"3F599C8B",
    x"3F599FDA",
    x"3F59A329",
    x"3F59A678",
    x"3F59A9C7",
    x"3F59AD15",
    x"3F59B064",
    x"3F59B3B2",
    x"3F59B700",
    x"3F59BA4E",
    x"3F59BD9C",
    x"3F59C0EA",
    x"3F59C438",
    x"3F59C785",
    x"3F59CAD3",
    x"3F59CE20",
    x"3F59D16D",
    x"3F59D4BA",
    x"3F59D807",
    x"3F59DB54",
    x"3F59DEA1",
    x"3F59E1ED",
    x"3F59E53A",
    x"3F59E886",
    x"3F59EBD2",
    x"3F59EF1E",
    x"3F59F26A",
    x"3F59F5B6",
    x"3F59F901",
    x"3F59FC4D",
    x"3F59FF98",
    x"3F5A02E3",
    x"3F5A062E",
    x"3F5A0979",
    x"3F5A0CC4",
    x"3F5A100F",
    x"3F5A1359",
    x"3F5A16A4",
    x"3F5A19EE",
    x"3F5A1D38",
    x"3F5A2082",
    x"3F5A23CC",
    x"3F5A2716",
    x"3F5A2A60",
    x"3F5A2DA9",
    x"3F5A30F2",
    x"3F5A343C",
    x"3F5A3785",
    x"3F5A3ACE",
    x"3F5A3E17",
    x"3F5A415F",
    x"3F5A44A8",
    x"3F5A47F0",
    x"3F5A4B39",
    x"3F5A4E81",
    x"3F5A51C9",
    x"3F5A5511",
    x"3F5A5859",
    x"3F5A5BA0",
    x"3F5A5EE8",
    x"3F5A622F",
    x"3F5A6577",
    x"3F5A68BE",
    x"3F5A6C05",
    x"3F5A6F4C",
    x"3F5A7292",
    x"3F5A75D9",
    x"3F5A791F",
    x"3F5A7C66",
    x"3F5A7FAC",
    x"3F5A82F2",
    x"3F5A8638",
    x"3F5A897E",
    x"3F5A8CC3",
    x"3F5A9009",
    x"3F5A934E",
    x"3F5A9694",
    x"3F5A99D9",
    x"3F5A9D1E",
    x"3F5AA063",
    x"3F5AA3A8",
    x"3F5AA6EC",
    x"3F5AAA31",
    x"3F5AAD75",
    x"3F5AB0B9",
    x"3F5AB3FD",
    x"3F5AB741",
    x"3F5ABA85",
    x"3F5ABDC9",
    x"3F5AC10D",
    x"3F5AC450",
    x"3F5AC793",
    x"3F5ACAD6",
    x"3F5ACE1A",
    x"3F5AD15C",
    x"3F5AD49F",
    x"3F5AD7E2",
    x"3F5ADB24",
    x"3F5ADE67",
    x"3F5AE1A9",
    x"3F5AE4EB",
    x"3F5AE82D",
    x"3F5AEB6F",
    x"3F5AEEB1",
    x"3F5AF1F2",
    x"3F5AF534",
    x"3F5AF875",
    x"3F5AFBB6",
    x"3F5AFEF7",
    x"3F5B0238",
    x"3F5B0579",
    x"3F5B08BA",
    x"3F5B0BFA",
    x"3F5B0F3B",
    x"3F5B127B",
    x"3F5B15BB",
    x"3F5B18FB",
    x"3F5B1C3B",
    x"3F5B1F7B",
    x"3F5B22BB",
    x"3F5B25FA",
    x"3F5B2939",
    x"3F5B2C79",
    x"3F5B2FB8",
    x"3F5B32F7",
    x"3F5B3636",
    x"3F5B3974",
    x"3F5B3CB3",
    x"3F5B3FF1",
    x"3F5B4330",
    x"3F5B466E",
    x"3F5B49AC",
    x"3F5B4CEA",
    x"3F5B5027",
    x"3F5B5365",
    x"3F5B56A3",
    x"3F5B59E0",
    x"3F5B5D1D",
    x"3F5B605A",
    x"3F5B6397",
    x"3F5B66D4",
    x"3F5B6A11",
    x"3F5B6D4D",
    x"3F5B708A",
    x"3F5B73C6",
    x"3F5B7702",
    x"3F5B7A3E",
    x"3F5B7D7A",
    x"3F5B80B6",
    x"3F5B83F2",
    x"3F5B872D",
    x"3F5B8A69",
    x"3F5B8DA4",
    x"3F5B90DF",
    x"3F5B941A",
    x"3F5B9755",
    x"3F5B9A90",
    x"3F5B9DCA",
    x"3F5BA105",
    x"3F5BA43F",
    x"3F5BA779",
    x"3F5BAAB3",
    x"3F5BADED",
    x"3F5BB127",
    x"3F5BB461",
    x"3F5BB79A",
    x"3F5BBAD4",
    x"3F5BBE0D",
    x"3F5BC146",
    x"3F5BC47F",
    x"3F5BC7B8",
    x"3F5BCAF1",
    x"3F5BCE29",
    x"3F5BD162",
    x"3F5BD49A",
    x"3F5BD7D3",
    x"3F5BDB0B",
    x"3F5BDE43",
    x"3F5BE17A",
    x"3F5BE4B2",
    x"3F5BE7EA",
    x"3F5BEB21",
    x"3F5BEE58",
    x"3F5BF190",
    x"3F5BF4C7",
    x"3F5BF7FD",
    x"3F5BFB34",
    x"3F5BFE6B",
    x"3F5C01A1",
    x"3F5C04D8",
    x"3F5C080E",
    x"3F5C0B44",
    x"3F5C0E7A",
    x"3F5C11B0",
    x"3F5C14E6",
    x"3F5C181B",
    x"3F5C1B51",
    x"3F5C1E86",
    x"3F5C21BB",
    x"3F5C24F0",
    x"3F5C2825",
    x"3F5C2B5A",
    x"3F5C2E8E",
    x"3F5C31C3",
    x"3F5C34F7",
    x"3F5C382B",
    x"3F5C3B60",
    x"3F5C3E94",
    x"3F5C41C7",
    x"3F5C44FB",
    x"3F5C482F",
    x"3F5C4B62",
    x"3F5C4E95",
    x"3F5C51C9",
    x"3F5C54FC",
    x"3F5C582F",
    x"3F5C5B61",
    x"3F5C5E94",
    x"3F5C61C7",
    x"3F5C64F9",
    x"3F5C682B",
    x"3F5C6B5D",
    x"3F5C6E8F",
    x"3F5C71C1",
    x"3F5C74F3",
    x"3F5C7824",
    x"3F5C7B56",
    x"3F5C7E87",
    x"3F5C81B8",
    x"3F5C84EA",
    x"3F5C881A",
    x"3F5C8B4B",
    x"3F5C8E7C",
    x"3F5C91AC",
    x"3F5C94DD",
    x"3F5C980D",
    x"3F5C9B3D",
    x"3F5C9E6D",
    x"3F5CA19D",
    x"3F5CA4CD",
    x"3F5CA7FC",
    x"3F5CAB2C",
    x"3F5CAE5B",
    x"3F5CB18A",
    x"3F5CB4B9",
    x"3F5CB7E8",
    x"3F5CBB17",
    x"3F5CBE46",
    x"3F5CC174",
    x"3F5CC4A3",
    x"3F5CC7D1",
    x"3F5CCAFF",
    x"3F5CCE2D",
    x"3F5CD15B",
    x"3F5CD489",
    x"3F5CD7B6",
    x"3F5CDAE4",
    x"3F5CDE11",
    x"3F5CE13E",
    x"3F5CE46B",
    x"3F5CE798",
    x"3F5CEAC5",
    x"3F5CEDF2",
    x"3F5CF11E",
    x"3F5CF44B",
    x"3F5CF777",
    x"3F5CFAA3",
    x"3F5CFDCF",
    x"3F5D00FB",
    x"3F5D0427",
    x"3F5D0752",
    x"3F5D0A7E",
    x"3F5D0DA9",
    x"3F5D10D4",
    x"3F5D13FF",
    x"3F5D172A",
    x"3F5D1A55",
    x"3F5D1D80",
    x"3F5D20AA",
    x"3F5D23D5",
    x"3F5D26FF",
    x"3F5D2A29",
    x"3F5D2D53",
    x"3F5D307D",
    x"3F5D33A7",
    x"3F5D36D0",
    x"3F5D39FA",
    x"3F5D3D23",
    x"3F5D404C",
    x"3F5D4376",
    x"3F5D469E",
    x"3F5D49C7",
    x"3F5D4CF0",
    x"3F5D5018",
    x"3F5D5341",
    x"3F5D5669",
    x"3F5D5991",
    x"3F5D5CB9",
    x"3F5D5FE1",
    x"3F5D6309",
    x"3F5D6631",
    x"3F5D6958",
    x"3F5D6C7F",
    x"3F5D6FA7",
    x"3F5D72CE",
    x"3F5D75F5",
    x"3F5D791B",
    x"3F5D7C42",
    x"3F5D7F69",
    x"3F5D828F",
    x"3F5D85B5",
    x"3F5D88DB",
    x"3F5D8C01",
    x"3F5D8F27",
    x"3F5D924D",
    x"3F5D9573",
    x"3F5D9898",
    x"3F5D9BBD",
    x"3F5D9EE3",
    x"3F5DA208",
    x"3F5DA52D",
    x"3F5DA851",
    x"3F5DAB76",
    x"3F5DAE9B",
    x"3F5DB1BF",
    x"3F5DB4E3",
    x"3F5DB807",
    x"3F5DBB2B",
    x"3F5DBE4F",
    x"3F5DC173",
    x"3F5DC497",
    x"3F5DC7BA",
    x"3F5DCADD",
    x"3F5DCE01",
    x"3F5DD124",
    x"3F5DD447",
    x"3F5DD769",
    x"3F5DDA8C",
    x"3F5DDDAF",
    x"3F5DE0D1",
    x"3F5DE3F3",
    x"3F5DE715",
    x"3F5DEA37",
    x"3F5DED59",
    x"3F5DF07B",
    x"3F5DF39D",
    x"3F5DF6BE",
    x"3F5DF9DF",
    x"3F5DFD01",
    x"3F5E0022",
    x"3F5E0343",
    x"3F5E0663",
    x"3F5E0984",
    x"3F5E0CA5",
    x"3F5E0FC5",
    x"3F5E12E5",
    x"3F5E1605",
    x"3F5E1925",
    x"3F5E1C45",
    x"3F5E1F65",
    x"3F5E2285",
    x"3F5E25A4",
    x"3F5E28C3",
    x"3F5E2BE3",
    x"3F5E2F02",
    x"3F5E3221",
    x"3F5E353F",
    x"3F5E385E",
    x"3F5E3B7D",
    x"3F5E3E9B",
    x"3F5E41B9",
    x"3F5E44D7",
    x"3F5E47F5",
    x"3F5E4B13",
    x"3F5E4E31",
    x"3F5E514E",
    x"3F5E546C",
    x"3F5E5789",
    x"3F5E5AA6",
    x"3F5E5DC3",
    x"3F5E60E0",
    x"3F5E63FD",
    x"3F5E671A",
    x"3F5E6A36",
    x"3F5E6D53",
    x"3F5E706F",
    x"3F5E738B",
    x"3F5E76A7",
    x"3F5E79C3",
    x"3F5E7CDE",
    x"3F5E7FFA",
    x"3F5E8316",
    x"3F5E8631",
    x"3F5E894C",
    x"3F5E8C67",
    x"3F5E8F82",
    x"3F5E929D",
    x"3F5E95B7",
    x"3F5E98D2",
    x"3F5E9BEC",
    x"3F5E9F06",
    x"3F5EA221",
    x"3F5EA53A",
    x"3F5EA854",
    x"3F5EAB6E",
    x"3F5EAE88",
    x"3F5EB1A1",
    x"3F5EB4BA",
    x"3F5EB7D3",
    x"3F5EBAEC",
    x"3F5EBE05",
    x"3F5EC11E",
    x"3F5EC437",
    x"3F5EC74F",
    x"3F5ECA68",
    x"3F5ECD80",
    x"3F5ED098",
    x"3F5ED3B0",
    x"3F5ED6C8",
    x"3F5ED9DF",
    x"3F5EDCF7",
    x"3F5EE00E",
    x"3F5EE326",
    x"3F5EE63D",
    x"3F5EE954",
    x"3F5EEC6B",
    x"3F5EEF81",
    x"3F5EF298",
    x"3F5EF5AE",
    x"3F5EF8C5",
    x"3F5EFBDB",
    x"3F5EFEF1",
    x"3F5F0207",
    x"3F5F051D",
    x"3F5F0833",
    x"3F5F0B48",
    x"3F5F0E5D",
    x"3F5F1173",
    x"3F5F1488",
    x"3F5F179D",
    x"3F5F1AB2",
    x"3F5F1DC6",
    x"3F5F20DB",
    x"3F5F23EF",
    x"3F5F2704",
    x"3F5F2A18",
    x"3F5F2D2C",
    x"3F5F3040",
    x"3F5F3354",
    x"3F5F3667",
    x"3F5F397B",
    x"3F5F3C8E",
    x"3F5F3FA2",
    x"3F5F42B5",
    x"3F5F45C8",
    x"3F5F48DB",
    x"3F5F4BED",
    x"3F5F4F00",
    x"3F5F5212",
    x"3F5F5525",
    x"3F5F5837",
    x"3F5F5B49",
    x"3F5F5E5B",
    x"3F5F616C",
    x"3F5F647E",
    x"3F5F6790",
    x"3F5F6AA1",
    x"3F5F6DB2",
    x"3F5F70C3",
    x"3F5F73D4",
    x"3F5F76E5",
    x"3F5F79F6",
    x"3F5F7D06",
    x"3F5F8017",
    x"3F5F8327",
    x"3F5F8637",
    x"3F5F8947",
    x"3F5F8C57",
    x"3F5F8F67",
    x"3F5F9276",
    x"3F5F9586",
    x"3F5F9895",
    x"3F5F9BA5",
    x"3F5F9EB4",
    x"3F5FA1C3",
    x"3F5FA4D1",
    x"3F5FA7E0",
    x"3F5FAAEF",
    x"3F5FADFD",
    x"3F5FB10B",
    x"3F5FB419",
    x"3F5FB727",
    x"3F5FBA35",
    x"3F5FBD43",
    x"3F5FC051",
    x"3F5FC35E",
    x"3F5FC66B",
    x"3F5FC979",
    x"3F5FCC86",
    x"3F5FCF93",
    x"3F5FD29F",
    x"3F5FD5AC",
    x"3F5FD8B8",
    x"3F5FDBC5",
    x"3F5FDED1",
    x"3F5FE1DD",
    x"3F5FE4E9",
    x"3F5FE7F5",
    x"3F5FEB01",
    x"3F5FEE0C",
    x"3F5FF118",
    x"3F5FF423",
    x"3F5FF72E",
    x"3F5FFA39",
    x"3F5FFD44",
    x"3F60004F",
    x"3F60035A",
    x"3F600664",
    x"3F60096E",
    x"3F600C79",
    x"3F600F83",
    x"3F60128D",
    x"3F601596",
    x"3F6018A0",
    x"3F601BAA",
    x"3F601EB3",
    x"3F6021BC",
    x"3F6024C6",
    x"3F6027CF",
    x"3F602AD7",
    x"3F602DE0",
    x"3F6030E9",
    x"3F6033F1",
    x"3F6036FA",
    x"3F603A02",
    x"3F603D0A",
    x"3F604012",
    x"3F60431A",
    x"3F604621",
    x"3F604929",
    x"3F604C30",
    x"3F604F37",
    x"3F60523E",
    x"3F605545",
    x"3F60584C",
    x"3F605B53",
    x"3F605E5A",
    x"3F606160",
    x"3F606466",
    x"3F60676D",
    x"3F606A73",
    x"3F606D78",
    x"3F60707E",
    x"3F607384",
    x"3F607689",
    x"3F60798F",
    x"3F607C94",
    x"3F607F99",
    x"3F60829E",
    x"3F6085A3",
    x"3F6088A7",
    x"3F608BAC",
    x"3F608EB0",
    x"3F6091B5",
    x"3F6094B9",
    x"3F6097BD",
    x"3F609AC1",
    x"3F609DC4",
    x"3F60A0C8",
    x"3F60A3CC",
    x"3F60A6CF",
    x"3F60A9D2",
    x"3F60ACD5",
    x"3F60AFD8",
    x"3F60B2DB",
    x"3F60B5DE",
    x"3F60B8E0",
    x"3F60BBE2",
    x"3F60BEE5",
    x"3F60C1E7",
    x"3F60C4E9",
    x"3F60C7EB",
    x"3F60CAEC",
    x"3F60CDEE",
    x"3F60D0EF",
    x"3F60D3F1",
    x"3F60D6F2",
    x"3F60D9F3",
    x"3F60DCF4",
    x"3F60DFF4",
    x"3F60E2F5",
    x"3F60E5F6",
    x"3F60E8F6",
    x"3F60EBF6",
    x"3F60EEF6",
    x"3F60F1F6",
    x"3F60F4F6",
    x"3F60F7F6",
    x"3F60FAF5",
    x"3F60FDF5",
    x"3F6100F4",
    x"3F6103F3",
    x"3F6106F2",
    x"3F6109F1",
    x"3F610CF0",
    x"3F610FEE",
    x"3F6112ED",
    x"3F6115EB",
    x"3F6118E9",
    x"3F611BE7",
    x"3F611EE5",
    x"3F6121E3",
    x"3F6124E1",
    x"3F6127DE",
    x"3F612ADB",
    x"3F612DD9",
    x"3F6130D6",
    x"3F6133D3",
    x"3F6136D0",
    x"3F6139CC",
    x"3F613CC9",
    x"3F613FC5",
    x"3F6142C1",
    x"3F6145BE",
    x"3F6148BA",
    x"3F614BB5",
    x"3F614EB1",
    x"3F6151AD",
    x"3F6154A8",
    x"3F6157A4",
    x"3F615A9F",
    x"3F615D9A",
    x"3F616095",
    x"3F616390",
    x"3F61668A",
    x"3F616985",
    x"3F616C7F",
    x"3F616F79",
    x"3F617274",
    x"3F61756E",
    x"3F617867",
    x"3F617B61",
    x"3F617E5B",
    x"3F618154",
    x"3F61844D",
    x"3F618747",
    x"3F618A40",
    x"3F618D38",
    x"3F619031",
    x"3F61932A",
    x"3F619622",
    x"3F61991B",
    x"3F619C13",
    x"3F619F0B",
    x"3F61A203",
    x"3F61A4FB",
    x"3F61A7F2",
    x"3F61AAEA",
    x"3F61ADE1",
    x"3F61B0D9",
    x"3F61B3D0",
    x"3F61B6C7",
    x"3F61B9BE",
    x"3F61BCB4",
    x"3F61BFAB",
    x"3F61C2A1",
    x"3F61C598",
    x"3F61C88E",
    x"3F61CB84",
    x"3F61CE7A",
    x"3F61D16F",
    x"3F61D465",
    x"3F61D75B",
    x"3F61DA50",
    x"3F61DD45",
    x"3F61E03A",
    x"3F61E32F",
    x"3F61E624",
    x"3F61E919",
    x"3F61EC0D",
    x"3F61EF02",
    x"3F61F1F6",
    x"3F61F4EA",
    x"3F61F7DE",
    x"3F61FAD2",
    x"3F61FDC6",
    x"3F6200B9",
    x"3F6203AD",
    x"3F6206A0",
    x"3F620993",
    x"3F620C86",
    x"3F620F79",
    x"3F62126C",
    x"3F62155E",
    x"3F621851",
    x"3F621B43",
    x"3F621E35",
    x"3F622128",
    x"3F62241A",
    x"3F62270B",
    x"3F6229FD",
    x"3F622CEF",
    x"3F622FE0",
    x"3F6232D1",
    x"3F6235C2",
    x"3F6238B3",
    x"3F623BA4",
    x"3F623E95",
    x"3F624186",
    x"3F624476",
    x"3F624766",
    x"3F624A57",
    x"3F624D47",
    x"3F625036",
    x"3F625326",
    x"3F625616",
    x"3F625905",
    x"3F625BF5",
    x"3F625EE4",
    x"3F6261D3",
    x"3F6264C2",
    x"3F6267B1",
    x"3F626AA0",
    x"3F626D8E",
    x"3F62707C",
    x"3F62736B",
    x"3F627659",
    x"3F627947",
    x"3F627C35",
    x"3F627F22",
    x"3F628210",
    x"3F6284FD",
    x"3F6287EB",
    x"3F628AD8",
    x"3F628DC5",
    x"3F6290B2",
    x"3F62939F",
    x"3F62968B",
    x"3F629978",
    x"3F629C64",
    x"3F629F50",
    x"3F62A23D",
    x"3F62A528",
    x"3F62A814",
    x"3F62AB00",
    x"3F62ADEB",
    x"3F62B0D7",
    x"3F62B3C2",
    x"3F62B6AD",
    x"3F62B998",
    x"3F62BC83",
    x"3F62BF6E",
    x"3F62C258",
    x"3F62C543",
    x"3F62C82D",
    x"3F62CB17",
    x"3F62CE01",
    x"3F62D0EB",
    x"3F62D3D5",
    x"3F62D6BF",
    x"3F62D9A8",
    x"3F62DC92",
    x"3F62DF7B",
    x"3F62E264",
    x"3F62E54D",
    x"3F62E836",
    x"3F62EB1E",
    x"3F62EE07",
    x"3F62F0EF",
    x"3F62F3D8",
    x"3F62F6C0",
    x"3F62F9A8",
    x"3F62FC8F",
    x"3F62FF77",
    x"3F63025F",
    x"3F630546",
    x"3F63082E",
    x"3F630B15",
    x"3F630DFC",
    x"3F6310E3",
    x"3F6313C9",
    x"3F6316B0",
    x"3F631996",
    x"3F631C7D",
    x"3F631F63",
    x"3F632249",
    x"3F63252F",
    x"3F632815",
    x"3F632AFB",
    x"3F632DE0",
    x"3F6330C5",
    x"3F6333AB",
    x"3F633690",
    x"3F633975",
    x"3F633C5A",
    x"3F633F3E",
    x"3F634223",
    x"3F634507",
    x"3F6347EC",
    x"3F634AD0",
    x"3F634DB4",
    x"3F635098",
    x"3F63537B",
    x"3F63565F",
    x"3F635943",
    x"3F635C26",
    x"3F635F09",
    x"3F6361EC",
    x"3F6364CF",
    x"3F6367B2",
    x"3F636A95",
    x"3F636D77",
    x"3F637059",
    x"3F63733C",
    x"3F63761E",
    x"3F637900",
    x"3F637BE2",
    x"3F637EC3",
    x"3F6381A5",
    x"3F638486",
    x"3F638767",
    x"3F638A49",
    x"3F638D2A",
    x"3F63900B",
    x"3F6392EB",
    x"3F6395CC",
    x"3F6398AC",
    x"3F639B8D",
    x"3F639E6D",
    x"3F63A14D",
    x"3F63A42D",
    x"3F63A70D",
    x"3F63A9EC",
    x"3F63ACCC",
    x"3F63AFAB",
    x"3F63B28A",
    x"3F63B569",
    x"3F63B848",
    x"3F63BB27",
    x"3F63BE06",
    x"3F63C0E4",
    x"3F63C3C3",
    x"3F63C6A1",
    x"3F63C97F",
    x"3F63CC5D",
    x"3F63CF3B",
    x"3F63D219",
    x"3F63D4F6",
    x"3F63D7D4",
    x"3F63DAB1",
    x"3F63DD8E",
    x"3F63E06B",
    x"3F63E348",
    x"3F63E625",
    x"3F63E901",
    x"3F63EBDE",
    x"3F63EEBA",
    x"3F63F196",
    x"3F63F473",
    x"3F63F74E",
    x"3F63FA2A",
    x"3F63FD06",
    x"3F63FFE1",
    x"3F6402BD",
    x"3F640598",
    x"3F640873",
    x"3F640B4E",
    x"3F640E29",
    x"3F641104",
    x"3F6413DE",
    x"3F6416B9",
    x"3F641993",
    x"3F641C6D",
    x"3F641F47",
    x"3F642221",
    x"3F6424FB",
    x"3F6427D4",
    x"3F642AAE",
    x"3F642D87",
    x"3F643060",
    x"3F643339",
    x"3F643612",
    x"3F6438EB",
    x"3F643BC4",
    x"3F643E9C",
    x"3F644174",
    x"3F64444D",
    x"3F644725",
    x"3F6449FD",
    x"3F644CD5",
    x"3F644FAC",
    x"3F645284",
    x"3F64555B",
    x"3F645832",
    x"3F645B0A",
    x"3F645DE1",
    x"3F6460B7",
    x"3F64638E",
    x"3F646665",
    x"3F64693B",
    x"3F646C11",
    x"3F646EE8",
    x"3F6471BE",
    x"3F647493",
    x"3F647769",
    x"3F647A3F",
    x"3F647D14",
    x"3F647FEA",
    x"3F6482BF",
    x"3F648594",
    x"3F648869",
    x"3F648B3E",
    x"3F648E12",
    x"3F6490E7",
    x"3F6493BB",
    x"3F64968F",
    x"3F649963",
    x"3F649C37",
    x"3F649F0B",
    x"3F64A1DF",
    x"3F64A4B2",
    x"3F64A786",
    x"3F64AA59",
    x"3F64AD2C",
    x"3F64AFFF",
    x"3F64B2D2",
    x"3F64B5A5",
    x"3F64B877",
    x"3F64BB4A",
    x"3F64BE1C",
    x"3F64C0EE",
    x"3F64C3C0",
    x"3F64C692",
    x"3F64C964",
    x"3F64CC35",
    x"3F64CF07",
    x"3F64D1D8",
    x"3F64D4AA",
    x"3F64D77B",
    x"3F64DA4B",
    x"3F64DD1C",
    x"3F64DFED",
    x"3F64E2BD",
    x"3F64E58E",
    x"3F64E85E",
    x"3F64EB2E",
    x"3F64EDFE",
    x"3F64F0CE",
    x"3F64F39E",
    x"3F64F66D",
    x"3F64F93D",
    x"3F64FC0C",
    x"3F64FEDB",
    x"3F6501AA",
    x"3F650479",
    x"3F650748",
    x"3F650A16",
    x"3F650CE5",
    x"3F650FB3",
    x"3F651281",
    x"3F65154F",
    x"3F65181D",
    x"3F651AEB",
    x"3F651DB8",
    x"3F652086",
    x"3F652353",
    x"3F652620",
    x"3F6528ED",
    x"3F652BBA",
    x"3F652E87",
    x"3F653154",
    x"3F653420",
    x"3F6536ED",
    x"3F6539B9",
    x"3F653C85",
    x"3F653F51",
    x"3F65421D",
    x"3F6544E8",
    x"3F6547B4",
    x"3F654A7F",
    x"3F654D4B",
    x"3F655016",
    x"3F6552E1",
    x"3F6555AC",
    x"3F655876",
    x"3F655B41",
    x"3F655E0B",
    x"3F6560D6",
    x"3F6563A0",
    x"3F65666A",
    x"3F656934",
    x"3F656BFD",
    x"3F656EC7",
    x"3F657190",
    x"3F65745A",
    x"3F657723",
    x"3F6579EC",
    x"3F657CB5",
    x"3F657F7E",
    x"3F658246",
    x"3F65850F",
    x"3F6587D7",
    x"3F658AA0",
    x"3F658D68",
    x"3F659030",
    x"3F6592F7",
    x"3F6595BF",
    x"3F659887",
    x"3F659B4E",
    x"3F659E15",
    x"3F65A0DC",
    x"3F65A3A3",
    x"3F65A66A",
    x"3F65A931",
    x"3F65ABF7",
    x"3F65AEBE",
    x"3F65B184",
    x"3F65B44A",
    x"3F65B710",
    x"3F65B9D6",
    x"3F65BC9C",
    x"3F65BF62",
    x"3F65C227",
    x"3F65C4EC",
    x"3F65C7B1",
    x"3F65CA77",
    x"3F65CD3B",
    x"3F65D000",
    x"3F65D2C5",
    x"3F65D589",
    x"3F65D84E",
    x"3F65DB12",
    x"3F65DDD6",
    x"3F65E09A",
    x"3F65E35E",
    x"3F65E621",
    x"3F65E8E5",
    x"3F65EBA8",
    x"3F65EE6C",
    x"3F65F12F",
    x"3F65F3F2",
    x"3F65F6B4",
    x"3F65F977",
    x"3F65FC3A",
    x"3F65FEFC",
    x"3F6601BE",
    x"3F660480",
    x"3F660742",
    x"3F660A04",
    x"3F660CC6",
    x"3F660F88",
    x"3F661249",
    x"3F66150A",
    x"3F6617CC",
    x"3F661A8D",
    x"3F661D4D",
    x"3F66200E",
    x"3F6622CF",
    x"3F66258F",
    x"3F662850",
    x"3F662B10",
    x"3F662DD0",
    x"3F663090",
    x"3F663350",
    x"3F66360F",
    x"3F6638CF",
    x"3F663B8E",
    x"3F663E4D",
    x"3F66410C",
    x"3F6643CB",
    x"3F66468A",
    x"3F664949",
    x"3F664C07",
    x"3F664EC6",
    x"3F665184",
    x"3F665442",
    x"3F665700",
    x"3F6659BE",
    x"3F665C7C",
    x"3F665F39",
    x"3F6661F7",
    x"3F6664B4",
    x"3F666771",
    x"3F666A2E",
    x"3F666CEB",
    x"3F666FA8",
    x"3F667264",
    x"3F667521",
    x"3F6677DD",
    x"3F667A99",
    x"3F667D55",
    x"3F668011",
    x"3F6682CD",
    x"3F668588",
    x"3F668844",
    x"3F668AFF",
    x"3F668DBA",
    x"3F669076",
    x"3F669330",
    x"3F6695EB",
    x"3F6698A6",
    x"3F669B60",
    x"3F669E1B",
    x"3F66A0D5",
    x"3F66A38F",
    x"3F66A649",
    x"3F66A903",
    x"3F66ABBC",
    x"3F66AE76",
    x"3F66B12F",
    x"3F66B3E9",
    x"3F66B6A2",
    x"3F66B95B",
    x"3F66BC14",
    x"3F66BECC",
    x"3F66C185",
    x"3F66C43D",
    x"3F66C6F6",
    x"3F66C9AE",
    x"3F66CC66",
    x"3F66CF1E",
    x"3F66D1D5",
    x"3F66D48D",
    x"3F66D744",
    x"3F66D9FC",
    x"3F66DCB3",
    x"3F66DF6A",
    x"3F66E221",
    x"3F66E4D7",
    x"3F66E78E",
    x"3F66EA45",
    x"3F66ECFB",
    x"3F66EFB1",
    x"3F66F267",
    x"3F66F51D",
    x"3F66F7D3",
    x"3F66FA88",
    x"3F66FD3E",
    x"3F66FFF3",
    x"3F6702A9",
    x"3F67055E",
    x"3F670813",
    x"3F670AC7",
    x"3F670D7C",
    x"3F671031",
    x"3F6712E5",
    x"3F671599",
    x"3F67184D",
    x"3F671B01",
    x"3F671DB5",
    x"3F672069",
    x"3F67231C",
    x"3F6725D0",
    x"3F672883",
    x"3F672B36",
    x"3F672DE9",
    x"3F67309C",
    x"3F67334F",
    x"3F673601",
    x"3F6738B4",
    x"3F673B66",
    x"3F673E18",
    x"3F6740CA",
    x"3F67437C",
    x"3F67462E",
    x"3F6748DF",
    x"3F674B91",
    x"3F674E42",
    x"3F6750F3",
    x"3F6753A5",
    x"3F675655",
    x"3F675906",
    x"3F675BB7",
    x"3F675E67",
    x"3F676118",
    x"3F6763C8",
    x"3F676678",
    x"3F676928",
    x"3F676BD8",
    x"3F676E87",
    x"3F677137",
    x"3F6773E6",
    x"3F677695",
    x"3F677944",
    x"3F677BF3",
    x"3F677EA2",
    x"3F678151",
    x"3F6783FF",
    x"3F6786AE",
    x"3F67895C",
    x"3F678C0A",
    x"3F678EB8",
    x"3F679166",
    x"3F679414",
    x"3F6796C1",
    x"3F67996F",
    x"3F679C1C",
    x"3F679EC9",
    x"3F67A176",
    x"3F67A423",
    x"3F67A6D0",
    x"3F67A97C",
    x"3F67AC29",
    x"3F67AED5",
    x"3F67B181",
    x"3F67B42D",
    x"3F67B6D9",
    x"3F67B985",
    x"3F67BC30",
    x"3F67BEDC",
    x"3F67C187",
    x"3F67C432",
    x"3F67C6DE",
    x"3F67C988",
    x"3F67CC33",
    x"3F67CEDE",
    x"3F67D188",
    x"3F67D433",
    x"3F67D6DD",
    x"3F67D987",
    x"3F67DC31",
    x"3F67DEDB",
    x"3F67E184",
    x"3F67E42E",
    x"3F67E6D7",
    x"3F67E980",
    x"3F67EC29",
    x"3F67EED2",
    x"3F67F17B",
    x"3F67F424",
    x"3F67F6CC",
    x"3F67F975",
    x"3F67FC1D",
    x"3F67FEC5",
    x"3F68016D",
    x"3F680415",
    x"3F6806BD",
    x"3F680964",
    x"3F680C0C",
    x"3F680EB3",
    x"3F68115A",
    x"3F681401",
    x"3F6816A8",
    x"3F68194F",
    x"3F681BF5",
    x"3F681E9C",
    x"3F682142",
    x"3F6823E8",
    x"3F68268E",
    x"3F682934",
    x"3F682BDA",
    x"3F682E7F",
    x"3F683125",
    x"3F6833CA",
    x"3F68366F",
    x"3F683914",
    x"3F683BB9",
    x"3F683E5E",
    x"3F684103",
    x"3F6843A7",
    x"3F68464B",
    x"3F6848F0",
    x"3F684B94",
    x"3F684E38",
    x"3F6850DB",
    x"3F68537F",
    x"3F685623",
    x"3F6858C6",
    x"3F685B69",
    x"3F685E0C",
    x"3F6860AF",
    x"3F686352",
    x"3F6865F5",
    x"3F686897",
    x"3F686B39",
    x"3F686DDC",
    x"3F68707E",
    x"3F687320",
    x"3F6875C2",
    x"3F687863",
    x"3F687B05",
    x"3F687DA6",
    x"3F688047",
    x"3F6882E9",
    x"3F68858A",
    x"3F68882A",
    x"3F688ACB",
    x"3F688D6C",
    x"3F68900C",
    x"3F6892AC",
    x"3F68954C",
    x"3F6897EC",
    x"3F689A8C",
    x"3F689D2C",
    x"3F689FCC",
    x"3F68A26B",
    x"3F68A50A",
    x"3F68A7AA",
    x"3F68AA49",
    x"3F68ACE7",
    x"3F68AF86",
    x"3F68B225",
    x"3F68B4C3",
    x"3F68B762",
    x"3F68BA00",
    x"3F68BC9E",
    x"3F68BF3C",
    x"3F68C1D9",
    x"3F68C477",
    x"3F68C714",
    x"3F68C9B2",
    x"3F68CC4F",
    x"3F68CEEC",
    x"3F68D189",
    x"3F68D426",
    x"3F68D6C2",
    x"3F68D95F",
    x"3F68DBFB",
    x"3F68DE97",
    x"3F68E134",
    x"3F68E3CF",
    x"3F68E66B",
    x"3F68E907",
    x"3F68EBA2",
    x"3F68EE3E",
    x"3F68F0D9",
    x"3F68F374",
    x"3F68F60F",
    x"3F68F8AA",
    x"3F68FB45",
    x"3F68FDDF",
    x"3F690079",
    x"3F690314",
    x"3F6905AE",
    x"3F690848",
    x"3F690AE2",
    x"3F690D7B",
    x"3F691015",
    x"3F6912AE",
    x"3F691547",
    x"3F6917E1",
    x"3F691A7A",
    x"3F691D12",
    x"3F691FAB",
    x"3F692244",
    x"3F6924DC",
    x"3F692774",
    x"3F692A0D",
    x"3F692CA5",
    x"3F692F3C",
    x"3F6931D4",
    x"3F69346C",
    x"3F693703",
    x"3F69399A",
    x"3F693C32",
    x"3F693EC9",
    x"3F694160",
    x"3F6943F6",
    x"3F69468D",
    x"3F694923",
    x"3F694BBA",
    x"3F694E50",
    x"3F6950E6",
    x"3F69537C",
    x"3F695611",
    x"3F6958A7",
    x"3F695B3D",
    x"3F695DD2",
    x"3F696067",
    x"3F6962FC",
    x"3F696591",
    x"3F696826",
    x"3F696ABA",
    x"3F696D4F",
    x"3F696FE3",
    x"3F697277",
    x"3F69750C",
    x"3F69779F",
    x"3F697A33",
    x"3F697CC7",
    x"3F697F5A",
    x"3F6981EE",
    x"3F698481",
    x"3F698714",
    x"3F6989A7",
    x"3F698C3A",
    x"3F698ECC",
    x"3F69915F",
    x"3F6993F1",
    x"3F699684",
    x"3F699916",
    x"3F699BA8",
    x"3F699E39",
    x"3F69A0CB",
    x"3F69A35D",
    x"3F69A5EE",
    x"3F69A87F",
    x"3F69AB10",
    x"3F69ADA1",
    x"3F69B032",
    x"3F69B2C3",
    x"3F69B553",
    x"3F69B7E4",
    x"3F69BA74",
    x"3F69BD04",
    x"3F69BF94",
    x"3F69C224",
    x"3F69C4B4",
    x"3F69C743",
    x"3F69C9D3",
    x"3F69CC62",
    x"3F69CEF1",
    x"3F69D180",
    x"3F69D40F",
    x"3F69D69E",
    x"3F69D92C",
    x"3F69DBBB",
    x"3F69DE49",
    x"3F69E0D7",
    x"3F69E365",
    x"3F69E5F3",
    x"3F69E881",
    x"3F69EB0E",
    x"3F69ED9C",
    x"3F69F029",
    x"3F69F2B6",
    x"3F69F543",
    x"3F69F7D0",
    x"3F69FA5D",
    x"3F69FCEA",
    x"3F69FF76",
    x"3F6A0202",
    x"3F6A048F",
    x"3F6A071B",
    x"3F6A09A7",
    x"3F6A0C32",
    x"3F6A0EBE",
    x"3F6A1149",
    x"3F6A13D5",
    x"3F6A1660",
    x"3F6A18EB",
    x"3F6A1B76",
    x"3F6A1E01",
    x"3F6A208B",
    x"3F6A2316",
    x"3F6A25A0",
    x"3F6A282A",
    x"3F6A2AB4",
    x"3F6A2D3E",
    x"3F6A2FC8",
    x"3F6A3252",
    x"3F6A34DB",
    x"3F6A3765",
    x"3F6A39EE",
    x"3F6A3C77",
    x"3F6A3F00",
    x"3F6A4189",
    x"3F6A4411",
    x"3F6A469A",
    x"3F6A4922",
    x"3F6A4BAA",
    x"3F6A4E33",
    x"3F6A50BA",
    x"3F6A5342",
    x"3F6A55CA",
    x"3F6A5851",
    x"3F6A5AD9",
    x"3F6A5D60",
    x"3F6A5FE7",
    x"3F6A626E",
    x"3F6A64F5",
    x"3F6A677C",
    x"3F6A6A02",
    x"3F6A6C89",
    x"3F6A6F0F",
    x"3F6A7195",
    x"3F6A741B",
    x"3F6A76A1",
    x"3F6A7926",
    x"3F6A7BAC",
    x"3F6A7E31",
    x"3F6A80B7",
    x"3F6A833C",
    x"3F6A85C1",
    x"3F6A8846",
    x"3F6A8ACA",
    x"3F6A8D4F",
    x"3F6A8FD3",
    x"3F6A9258",
    x"3F6A94DC",
    x"3F6A9760",
    x"3F6A99E4",
    x"3F6A9C67",
    x"3F6A9EEB",
    x"3F6AA16E",
    x"3F6AA3F2",
    x"3F6AA675",
    x"3F6AA8F8",
    x"3F6AAB7B",
    x"3F6AADFD",
    x"3F6AB080",
    x"3F6AB302",
    x"3F6AB585",
    x"3F6AB807",
    x"3F6ABA89",
    x"3F6ABD0B",
    x"3F6ABF8C",
    x"3F6AC20E",
    x"3F6AC48F",
    x"3F6AC711",
    x"3F6AC992",
    x"3F6ACC13",
    x"3F6ACE94",
    x"3F6AD115",
    x"3F6AD395",
    x"3F6AD616",
    x"3F6AD896",
    x"3F6ADB16",
    x"3F6ADD96",
    x"3F6AE016",
    x"3F6AE296",
    x"3F6AE515",
    x"3F6AE795",
    x"3F6AEA14",
    x"3F6AEC93",
    x"3F6AEF12",
    x"3F6AF191",
    x"3F6AF410",
    x"3F6AF68F",
    x"3F6AF90D",
    x"3F6AFB8C",
    x"3F6AFE0A",
    x"3F6B0088",
    x"3F6B0306",
    x"3F6B0584",
    x"3F6B0801",
    x"3F6B0A7F",
    x"3F6B0CFC",
    x"3F6B0F79",
    x"3F6B11F6",
    x"3F6B1473",
    x"3F6B16F0",
    x"3F6B196D",
    x"3F6B1BE9",
    x"3F6B1E65",
    x"3F6B20E2",
    x"3F6B235E",
    x"3F6B25DA",
    x"3F6B2855",
    x"3F6B2AD1",
    x"3F6B2D4D",
    x"3F6B2FC8",
    x"3F6B3243",
    x"3F6B34BE",
    x"3F6B3739",
    x"3F6B39B4",
    x"3F6B3C2F",
    x"3F6B3EA9",
    x"3F6B4124",
    x"3F6B439E",
    x"3F6B4618",
    x"3F6B4892",
    x"3F6B4B0C",
    x"3F6B4D85",
    x"3F6B4FFF",
    x"3F6B5278",
    x"3F6B54F1",
    x"3F6B576B",
    x"3F6B59E3",
    x"3F6B5C5C",
    x"3F6B5ED5",
    x"3F6B614D",
    x"3F6B63C6",
    x"3F6B663E",
    x"3F6B68B6",
    x"3F6B6B2E",
    x"3F6B6DA6",
    x"3F6B701E",
    x"3F6B7295",
    x"3F6B750D",
    x"3F6B7784",
    x"3F6B79FB",
    x"3F6B7C72",
    x"3F6B7EE9",
    x"3F6B815F",
    x"3F6B83D6",
    x"3F6B864C",
    x"3F6B88C3",
    x"3F6B8B39",
    x"3F6B8DAF",
    x"3F6B9025",
    x"3F6B929A",
    x"3F6B9510",
    x"3F6B9785",
    x"3F6B99FB",
    x"3F6B9C70",
    x"3F6B9EE5",
    x"3F6BA159",
    x"3F6BA3CE",
    x"3F6BA643",
    x"3F6BA8B7",
    x"3F6BAB2B",
    x"3F6BADA0",
    x"3F6BB014",
    x"3F6BB287",
    x"3F6BB4FB",
    x"3F6BB76F",
    x"3F6BB9E2",
    x"3F6BBC55",
    x"3F6BBEC8",
    x"3F6BC13B",
    x"3F6BC3AE",
    x"3F6BC621",
    x"3F6BC894",
    x"3F6BCB06",
    x"3F6BCD78",
    x"3F6BCFEA",
    x"3F6BD25C",
    x"3F6BD4CE",
    x"3F6BD740",
    x"3F6BD9B2",
    x"3F6BDC23",
    x"3F6BDE94",
    x"3F6BE105",
    x"3F6BE376",
    x"3F6BE5E7",
    x"3F6BE858",
    x"3F6BEAC9",
    x"3F6BED39",
    x"3F6BEFA9",
    x"3F6BF21A",
    x"3F6BF48A",
    x"3F6BF6F9",
    x"3F6BF969",
    x"3F6BFBD9",
    x"3F6BFE48",
    x"3F6C00B7",
    x"3F6C0327",
    x"3F6C0596",
    x"3F6C0805",
    x"3F6C0A73",
    x"3F6C0CE2",
    x"3F6C0F50",
    x"3F6C11BF",
    x"3F6C142D",
    x"3F6C169B",
    x"3F6C1909",
    x"3F6C1B76",
    x"3F6C1DE4",
    x"3F6C2051",
    x"3F6C22BF",
    x"3F6C252C",
    x"3F6C2799",
    x"3F6C2A06",
    x"3F6C2C73",
    x"3F6C2EDF",
    x"3F6C314C",
    x"3F6C33B8",
    x"3F6C3624",
    x"3F6C3890",
    x"3F6C3AFC",
    x"3F6C3D68",
    x"3F6C3FD3",
    x"3F6C423F",
    x"3F6C44AA",
    x"3F6C4715",
    x"3F6C4980",
    x"3F6C4BEB",
    x"3F6C4E56",
    x"3F6C50C1",
    x"3F6C532B",
    x"3F6C5595",
    x"3F6C5800",
    x"3F6C5A6A",
    x"3F6C5CD4",
    x"3F6C5F3D",
    x"3F6C61A7",
    x"3F6C6410",
    x"3F6C667A",
    x"3F6C68E3",
    x"3F6C6B4C",
    x"3F6C6DB5",
    x"3F6C701E",
    x"3F6C7286",
    x"3F6C74EF",
    x"3F6C7757",
    x"3F6C79BF",
    x"3F6C7C27",
    x"3F6C7E8F",
    x"3F6C80F7",
    x"3F6C835E",
    x"3F6C85C6",
    x"3F6C882D",
    x"3F6C8A94",
    x"3F6C8CFC",
    x"3F6C8F62",
    x"3F6C91C9",
    x"3F6C9430",
    x"3F6C9696",
    x"3F6C98FD",
    x"3F6C9B63",
    x"3F6C9DC9",
    x"3F6CA02F",
    x"3F6CA295",
    x"3F6CA4FA",
    x"3F6CA760",
    x"3F6CA9C5",
    x"3F6CAC2A",
    x"3F6CAE8F",
    x"3F6CB0F4",
    x"3F6CB359",
    x"3F6CB5BD",
    x"3F6CB822",
    x"3F6CBA86",
    x"3F6CBCEA",
    x"3F6CBF4F",
    x"3F6CC1B2",
    x"3F6CC416",
    x"3F6CC67A",
    x"3F6CC8DD",
    x"3F6CCB41",
    x"3F6CCDA4",
    x"3F6CD007",
    x"3F6CD26A",
    x"3F6CD4CD",
    x"3F6CD72F",
    x"3F6CD992",
    x"3F6CDBF4",
    x"3F6CDE56",
    x"3F6CE0B8",
    x"3F6CE31A",
    x"3F6CE57C",
    x"3F6CE7DE",
    x"3F6CEA3F",
    x"3F6CECA0",
    x"3F6CEF02",
    x"3F6CF163",
    x"3F6CF3C4",
    x"3F6CF624",
    x"3F6CF885",
    x"3F6CFAE5",
    x"3F6CFD46",
    x"3F6CFFA6",
    x"3F6D0206",
    x"3F6D0466",
    x"3F6D06C6",
    x"3F6D0925",
    x"3F6D0B85",
    x"3F6D0DE4",
    x"3F6D1043",
    x"3F6D12A2",
    x"3F6D1501",
    x"3F6D1760",
    x"3F6D19BF",
    x"3F6D1C1D",
    x"3F6D1E7C",
    x"3F6D20DA",
    x"3F6D2338",
    x"3F6D2596",
    x"3F6D27F4",
    x"3F6D2A51",
    x"3F6D2CAF",
    x"3F6D2F0C",
    x"3F6D3169",
    x"3F6D33C6",
    x"3F6D3623",
    x"3F6D3880",
    x"3F6D3ADD",
    x"3F6D3D39",
    x"3F6D3F95",
    x"3F6D41F2",
    x"3F6D444E",
    x"3F6D46AA",
    x"3F6D4905",
    x"3F6D4B61",
    x"3F6D4DBC",
    x"3F6D5018",
    x"3F6D5273",
    x"3F6D54CE",
    x"3F6D5729",
    x"3F6D5984",
    x"3F6D5BDE",
    x"3F6D5E39",
    x"3F6D6093",
    x"3F6D62ED",
    x"3F6D6547",
    x"3F6D67A1",
    x"3F6D69FB",
    x"3F6D6C55",
    x"3F6D6EAE",
    x"3F6D7108",
    x"3F6D7361",
    x"3F6D75BA",
    x"3F6D7813",
    x"3F6D7A6C",
    x"3F6D7CC4",
    x"3F6D7F1D",
    x"3F6D8175",
    x"3F6D83CD",
    x"3F6D8625",
    x"3F6D887D",
    x"3F6D8AD5",
    x"3F6D8D2D",
    x"3F6D8F84",
    x"3F6D91DB",
    x"3F6D9433",
    x"3F6D968A",
    x"3F6D98E1",
    x"3F6D9B37",
    x"3F6D9D8E",
    x"3F6D9FE4",
    x"3F6DA23B",
    x"3F6DA491",
    x"3F6DA6E7",
    x"3F6DA93D",
    x"3F6DAB93",
    x"3F6DADE8",
    x"3F6DB03E",
    x"3F6DB293",
    x"3F6DB4E8",
    x"3F6DB73D",
    x"3F6DB992",
    x"3F6DBBE7",
    x"3F6DBE3C",
    x"3F6DC090",
    x"3F6DC2E4",
    x"3F6DC539",
    x"3F6DC78D",
    x"3F6DC9E1",
    x"3F6DCC34",
    x"3F6DCE88",
    x"3F6DD0DB",
    x"3F6DD32F",
    x"3F6DD582",
    x"3F6DD7D5",
    x"3F6DDA28",
    x"3F6DDC7B",
    x"3F6DDECD",
    x"3F6DE120",
    x"3F6DE372",
    x"3F6DE5C4",
    x"3F6DE816",
    x"3F6DEA68",
    x"3F6DECBA",
    x"3F6DEF0B",
    x"3F6DF15D",
    x"3F6DF3AE",
    x"3F6DF5FF",
    x"3F6DF850",
    x"3F6DFAA1",
    x"3F6DFCF2",
    x"3F6DFF43",
    x"3F6E0193",
    x"3F6E03E3",
    x"3F6E0634",
    x"3F6E0884",
    x"3F6E0AD4",
    x"3F6E0D23",
    x"3F6E0F73",
    x"3F6E11C2",
    x"3F6E1412",
    x"3F6E1661",
    x"3F6E18B0",
    x"3F6E1AFF",
    x"3F6E1D4E",
    x"3F6E1F9C",
    x"3F6E21EB",
    x"3F6E2439",
    x"3F6E2687",
    x"3F6E28D5",
    x"3F6E2B23",
    x"3F6E2D71",
    x"3F6E2FBE",
    x"3F6E320C",
    x"3F6E3459",
    x"3F6E36A6",
    x"3F6E38F3",
    x"3F6E3B40",
    x"3F6E3D8D",
    x"3F6E3FD9",
    x"3F6E4226",
    x"3F6E4472",
    x"3F6E46BE",
    x"3F6E490A",
    x"3F6E4B56",
    x"3F6E4DA2",
    x"3F6E4FEE",
    x"3F6E5239",
    x"3F6E5484",
    x"3F6E56CF",
    x"3F6E591A",
    x"3F6E5B65",
    x"3F6E5DB0",
    x"3F6E5FFB",
    x"3F6E6245",
    x"3F6E648F",
    x"3F6E66D9",
    x"3F6E6924",
    x"3F6E6B6D",
    x"3F6E6DB7",
    x"3F6E7001",
    x"3F6E724A",
    x"3F6E7493",
    x"3F6E76DD",
    x"3F6E7926",
    x"3F6E7B6E",
    x"3F6E7DB7",
    x"3F6E8000",
    x"3F6E8248",
    x"3F6E8490",
    x"3F6E86D8",
    x"3F6E8920",
    x"3F6E8B68",
    x"3F6E8DB0",
    x"3F6E8FF8",
    x"3F6E923F",
    x"3F6E9486",
    x"3F6E96CD",
    x"3F6E9914",
    x"3F6E9B5B",
    x"3F6E9DA2",
    x"3F6E9FE9",
    x"3F6EA22F",
    x"3F6EA475",
    x"3F6EA6BB",
    x"3F6EA901",
    x"3F6EAB47",
    x"3F6EAD8D",
    x"3F6EAFD2",
    x"3F6EB218",
    x"3F6EB45D",
    x"3F6EB6A2",
    x"3F6EB8E7",
    x"3F6EBB2C",
    x"3F6EBD71",
    x"3F6EBFB5",
    x"3F6EC1FA",
    x"3F6EC43E",
    x"3F6EC682",
    x"3F6EC8C6",
    x"3F6ECB0A",
    x"3F6ECD4D",
    x"3F6ECF91",
    x"3F6ED1D4",
    x"3F6ED418",
    x"3F6ED65B",
    x"3F6ED89E",
    x"3F6EDAE1",
    x"3F6EDD23",
    x"3F6EDF66",
    x"3F6EE1A8",
    x"3F6EE3EA",
    x"3F6EE62C",
    x"3F6EE86E",
    x"3F6EEAB0",
    x"3F6EECF2",
    x"3F6EEF33",
    x"3F6EF175",
    x"3F6EF3B6",
    x"3F6EF5F7",
    x"3F6EF838",
    x"3F6EFA79",
    x"3F6EFCBA",
    x"3F6EFEFA",
    x"3F6F013A",
    x"3F6F037B",
    x"3F6F05BB",
    x"3F6F07FB",
    x"3F6F0A3A",
    x"3F6F0C7A",
    x"3F6F0EBA",
    x"3F6F10F9",
    x"3F6F1338",
    x"3F6F1577",
    x"3F6F17B6",
    x"3F6F19F5",
    x"3F6F1C34",
    x"3F6F1E72",
    x"3F6F20B0",
    x"3F6F22EF",
    x"3F6F252D",
    x"3F6F276B",
    x"3F6F29A8",
    x"3F6F2BE6",
    x"3F6F2E24",
    x"3F6F3061",
    x"3F6F329E",
    x"3F6F34DB",
    x"3F6F3718",
    x"3F6F3955",
    x"3F6F3B92",
    x"3F6F3DCE",
    x"3F6F400A",
    x"3F6F4247",
    x"3F6F4483",
    x"3F6F46BE",
    x"3F6F48FA",
    x"3F6F4B36",
    x"3F6F4D71",
    x"3F6F4FAD",
    x"3F6F51E8",
    x"3F6F5423",
    x"3F6F565E",
    x"3F6F5899",
    x"3F6F5AD3",
    x"3F6F5D0E",
    x"3F6F5F48",
    x"3F6F6182",
    x"3F6F63BC",
    x"3F6F65F6",
    x"3F6F6830",
    x"3F6F6A69",
    x"3F6F6CA3",
    x"3F6F6EDC",
    x"3F6F7115",
    x"3F6F734E",
    x"3F6F7587",
    x"3F6F77C0",
    x"3F6F79F8",
    x"3F6F7C31",
    x"3F6F7E69",
    x"3F6F80A1",
    x"3F6F82D9",
    x"3F6F8511",
    x"3F6F8749",
    x"3F6F8981",
    x"3F6F8BB8",
    x"3F6F8DEF",
    x"3F6F9026",
    x"3F6F925D",
    x"3F6F9494",
    x"3F6F96CB",
    x"3F6F9902",
    x"3F6F9B38",
    x"3F6F9D6E",
    x"3F6F9FA4",
    x"3F6FA1DA",
    x"3F6FA410",
    x"3F6FA646",
    x"3F6FA87C",
    x"3F6FAAB1",
    x"3F6FACE6",
    x"3F6FAF1B",
    x"3F6FB150",
    x"3F6FB385",
    x"3F6FB5BA",
    x"3F6FB7EE",
    x"3F6FBA23",
    x"3F6FBC57",
    x"3F6FBE8B",
    x"3F6FC0BF",
    x"3F6FC2F3",
    x"3F6FC527",
    x"3F6FC75A",
    x"3F6FC98E",
    x"3F6FCBC1",
    x"3F6FCDF4",
    x"3F6FD027",
    x"3F6FD25A",
    x"3F6FD48C",
    x"3F6FD6BF",
    x"3F6FD8F1",
    x"3F6FDB24",
    x"3F6FDD56",
    x"3F6FDF88",
    x"3F6FE1B9",
    x"3F6FE3EB",
    x"3F6FE61D",
    x"3F6FE84E",
    x"3F6FEA7F",
    x"3F6FECB0",
    x"3F6FEEE1",
    x"3F6FF112",
    x"3F6FF343",
    x"3F6FF573",
    x"3F6FF7A3",
    x"3F6FF9D4",
    x"3F6FFC04",
    x"3F6FFE34",
    x"3F700063",
    x"3F700293",
    x"3F7004C3",
    x"3F7006F2",
    x"3F700921",
    x"3F700B50",
    x"3F700D7F",
    x"3F700FAE",
    x"3F7011DC",
    x"3F70140B",
    x"3F701639",
    x"3F701867",
    x"3F701A95",
    x"3F701CC3",
    x"3F701EF1",
    x"3F70211F",
    x"3F70234C",
    x"3F70257A",
    x"3F7027A7",
    x"3F7029D4",
    x"3F702C01",
    x"3F702E2D",
    x"3F70305A",
    x"3F703286",
    x"3F7034B3",
    x"3F7036DF",
    x"3F70390B",
    x"3F703B37",
    x"3F703D63",
    x"3F703F8E",
    x"3F7041BA",
    x"3F7043E5",
    x"3F704610",
    x"3F70483B",
    x"3F704A66",
    x"3F704C91",
    x"3F704EBB",
    x"3F7050E6",
    x"3F705310",
    x"3F70553A",
    x"3F705764",
    x"3F70598E",
    x"3F705BB8",
    x"3F705DE1",
    x"3F70600A",
    x"3F706234",
    x"3F70645D",
    x"3F706686",
    x"3F7068AF",
    x"3F706AD7",
    x"3F706D00",
    x"3F706F28",
    x"3F707151",
    x"3F707379",
    x"3F7075A1",
    x"3F7077C8",
    x"3F7079F0",
    x"3F707C18",
    x"3F707E3F",
    x"3F708066",
    x"3F70828D",
    x"3F7084B4",
    x"3F7086DB",
    x"3F708902",
    x"3F708B28",
    x"3F708D4F",
    x"3F708F75",
    x"3F70919B",
    x"3F7093C1",
    x"3F7095E7",
    x"3F70980C",
    x"3F709A32",
    x"3F709C57",
    x"3F709E7C",
    x"3F70A0A2",
    x"3F70A2C6",
    x"3F70A4EB",
    x"3F70A710",
    x"3F70A934",
    x"3F70AB59",
    x"3F70AD7D",
    x"3F70AFA1",
    x"3F70B1C5",
    x"3F70B3E9",
    x"3F70B60C",
    x"3F70B830",
    x"3F70BA53",
    x"3F70BC76",
    x"3F70BE99",
    x"3F70C0BC",
    x"3F70C2DF",
    x"3F70C501",
    x"3F70C724",
    x"3F70C946",
    x"3F70CB68",
    x"3F70CD8A",
    x"3F70CFAC",
    x"3F70D1CE",
    x"3F70D3F0",
    x"3F70D611",
    x"3F70D832",
    x"3F70DA54",
    x"3F70DC75",
    x"3F70DE95",
    x"3F70E0B6",
    x"3F70E2D7",
    x"3F70E4F7",
    x"3F70E717",
    x"3F70E938",
    x"3F70EB58",
    x"3F70ED77",
    x"3F70EF97",
    x"3F70F1B7",
    x"3F70F3D6",
    x"3F70F5F5",
    x"3F70F814",
    x"3F70FA33",
    x"3F70FC52",
    x"3F70FE71",
    x"3F71008F",
    x"3F7102AE",
    x"3F7104CC",
    x"3F7106EA",
    x"3F710908",
    x"3F710B26",
    x"3F710D44",
    x"3F710F61",
    x"3F71117F",
    x"3F71139C",
    x"3F7115B9",
    x"3F7117D6",
    x"3F7119F3",
    x"3F711C0F",
    x"3F711E2C",
    x"3F712048",
    x"3F712264",
    x"3F712480",
    x"3F71269C",
    x"3F7128B8",
    x"3F712AD4",
    x"3F712CEF",
    x"3F712F0B",
    x"3F713126",
    x"3F713341",
    x"3F71355C",
    x"3F713776",
    x"3F713991",
    x"3F713BAC",
    x"3F713DC6",
    x"3F713FE0",
    x"3F7141FA",
    x"3F714414",
    x"3F71462E",
    x"3F714847",
    x"3F714A61",
    x"3F714C7A",
    x"3F714E93",
    x"3F7150AC",
    x"3F7152C5",
    x"3F7154DE",
    x"3F7156F6",
    x"3F71590F",
    x"3F715B27",
    x"3F715D3F",
    x"3F715F57",
    x"3F71616F",
    x"3F716387",
    x"3F71659F",
    x"3F7167B6",
    x"3F7169CD",
    x"3F716BE4",
    x"3F716DFB",
    x"3F717012",
    x"3F717229",
    x"3F71743F",
    x"3F717656",
    x"3F71786C",
    x"3F717A82",
    x"3F717C98",
    x"3F717EAE",
    x"3F7180C4",
    x"3F7182D9",
    x"3F7184EF",
    x"3F718704",
    x"3F718919",
    x"3F718B2E",
    x"3F718D43",
    x"3F718F57",
    x"3F71916C",
    x"3F719380",
    x"3F719594",
    x"3F7197A8",
    x"3F7199BC",
    x"3F719BD0",
    x"3F719DE4",
    x"3F719FF7",
    x"3F71A20B",
    x"3F71A41E",
    x"3F71A631",
    x"3F71A844",
    x"3F71AA57",
    x"3F71AC69",
    x"3F71AE7C",
    x"3F71B08E",
    x"3F71B2A0",
    x"3F71B4B2",
    x"3F71B6C4",
    x"3F71B8D6",
    x"3F71BAE7",
    x"3F71BCF9",
    x"3F71BF0A",
    x"3F71C11B",
    x"3F71C32C",
    x"3F71C53D",
    x"3F71C74E",
    x"3F71C95F",
    x"3F71CB6F",
    x"3F71CD7F",
    x"3F71CF8F",
    x"3F71D19F",
    x"3F71D3AF",
    x"3F71D5BF",
    x"3F71D7CF",
    x"3F71D9DE",
    x"3F71DBED",
    x"3F71DDFC",
    x"3F71E00B",
    x"3F71E21A",
    x"3F71E429",
    x"3F71E637",
    x"3F71E846",
    x"3F71EA54",
    x"3F71EC62",
    x"3F71EE70",
    x"3F71F07E",
    x"3F71F28C",
    x"3F71F499",
    x"3F71F6A6",
    x"3F71F8B4",
    x"3F71FAC1",
    x"3F71FCCE",
    x"3F71FEDA",
    x"3F7200E7",
    x"3F7202F4",
    x"3F720500",
    x"3F72070C",
    x"3F720918",
    x"3F720B24",
    x"3F720D30",
    x"3F720F3C",
    x"3F721147",
    x"3F721352",
    x"3F72155E",
    x"3F721769",
    x"3F721973",
    x"3F721B7E",
    x"3F721D89",
    x"3F721F93",
    x"3F72219E",
    x"3F7223A8",
    x"3F7225B2",
    x"3F7227BC",
    x"3F7229C5",
    x"3F722BCF",
    x"3F722DD8",
    x"3F722FE2",
    x"3F7231EB",
    x"3F7233F4",
    x"3F7235FD",
    x"3F723805",
    x"3F723A0E",
    x"3F723C16",
    x"3F723E1F",
    x"3F724027",
    x"3F72422F",
    x"3F724437",
    x"3F72463E",
    x"3F724846",
    x"3F724A4D",
    x"3F724C54",
    x"3F724E5C",
    x"3F725063",
    x"3F725269",
    x"3F725470",
    x"3F725677",
    x"3F72587D",
    x"3F725A83",
    x"3F725C89",
    x"3F725E8F",
    x"3F726095",
    x"3F72629B",
    x"3F7264A0",
    x"3F7266A5",
    x"3F7268AB",
    x"3F726AB0",
    x"3F726CB5",
    x"3F726EB9",
    x"3F7270BE",
    x"3F7272C2",
    x"3F7274C7",
    x"3F7276CB",
    x"3F7278CF",
    x"3F727AD3",
    x"3F727CD7",
    x"3F727EDA",
    x"3F7280DE",
    x"3F7282E1",
    x"3F7284E4",
    x"3F7286E7",
    x"3F7288EA",
    x"3F728AED",
    x"3F728CEF",
    x"3F728EF2",
    x"3F7290F4",
    x"3F7292F6",
    x"3F7294F8",
    x"3F7296FA",
    x"3F7298FC",
    x"3F729AFD",
    x"3F729CFF",
    x"3F729F00",
    x"3F72A101",
    x"3F72A302",
    x"3F72A503",
    x"3F72A703",
    x"3F72A904",
    x"3F72AB04",
    x"3F72AD05",
    x"3F72AF05",
    x"3F72B105",
    x"3F72B304",
    x"3F72B504",
    x"3F72B704",
    x"3F72B903",
    x"3F72BB02",
    x"3F72BD01",
    x"3F72BF00",
    x"3F72C0FF",
    x"3F72C2FE",
    x"3F72C4FC",
    x"3F72C6FA",
    x"3F72C8F9",
    x"3F72CAF7",
    x"3F72CCF5",
    x"3F72CEF2",
    x"3F72D0F0",
    x"3F72D2ED",
    x"3F72D4EB",
    x"3F72D6E8",
    x"3F72D8E5",
    x"3F72DAE2",
    x"3F72DCDE",
    x"3F72DEDB",
    x"3F72E0D7",
    x"3F72E2D4",
    x"3F72E4D0",
    x"3F72E6CC",
    x"3F72E8C8",
    x"3F72EAC3",
    x"3F72ECBF",
    x"3F72EEBA",
    x"3F72F0B6",
    x"3F72F2B1",
    x"3F72F4AC",
    x"3F72F6A7",
    x"3F72F8A1",
    x"3F72FA9C",
    x"3F72FC96",
    x"3F72FE90",
    x"3F73008B",
    x"3F730284",
    x"3F73047E",
    x"3F730678",
    x"3F730871",
    x"3F730A6B",
    x"3F730C64",
    x"3F730E5D",
    x"3F731056",
    x"3F73124F",
    x"3F731447",
    x"3F731640",
    x"3F731838",
    x"3F731A30",
    x"3F731C28",
    x"3F731E20",
    x"3F732018",
    x"3F732210",
    x"3F732407",
    x"3F7325FE",
    x"3F7327F6",
    x"3F7329ED",
    x"3F732BE4",
    x"3F732DDA",
    x"3F732FD1",
    x"3F7331C7",
    x"3F7333BE",
    x"3F7335B4",
    x"3F7337AA",
    x"3F7339A0",
    x"3F733B95",
    x"3F733D8B",
    x"3F733F80",
    x"3F734175",
    x"3F73436B",
    x"3F734560",
    x"3F734754",
    x"3F734949",
    x"3F734B3E",
    x"3F734D32",
    x"3F734F26",
    x"3F73511A",
    x"3F73530E",
    x"3F735502",
    x"3F7356F6",
    x"3F7358E9",
    x"3F735ADC",
    x"3F735CD0",
    x"3F735EC3",
    x"3F7360B6",
    x"3F7362A8",
    x"3F73649B",
    x"3F73668E",
    x"3F736880",
    x"3F736A72",
    x"3F736C64",
    x"3F736E56",
    x"3F737048",
    x"3F737239",
    x"3F73742B",
    x"3F73761C",
    x"3F73780D",
    x"3F7379FE",
    x"3F737BEF",
    x"3F737DE0",
    x"3F737FD0",
    x"3F7381C1",
    x"3F7383B1",
    x"3F7385A1",
    x"3F738791",
    x"3F738981",
    x"3F738B71",
    x"3F738D60",
    x"3F738F50",
    x"3F73913F",
    x"3F73932E",
    x"3F73951D",
    x"3F73970C",
    x"3F7398FA",
    x"3F739AE9",
    x"3F739CD7",
    x"3F739EC5",
    x"3F73A0B4",
    x"3F73A2A1",
    x"3F73A48F",
    x"3F73A67D",
    x"3F73A86A",
    x"3F73AA58",
    x"3F73AC45",
    x"3F73AE32",
    x"3F73B01F",
    x"3F73B20C",
    x"3F73B3F8",
    x"3F73B5E5",
    x"3F73B7D1",
    x"3F73B9BD",
    x"3F73BBA9",
    x"3F73BD95",
    x"3F73BF81",
    x"3F73C16C",
    x"3F73C358",
    x"3F73C543",
    x"3F73C72E",
    x"3F73C919",
    x"3F73CB04",
    x"3F73CCEF",
    x"3F73CED9",
    x"3F73D0C4",
    x"3F73D2AE",
    x"3F73D498",
    x"3F73D682",
    x"3F73D86C",
    x"3F73DA56",
    x"3F73DC3F",
    x"3F73DE28",
    x"3F73E012",
    x"3F73E1FB",
    x"3F73E3E4",
    x"3F73E5CC",
    x"3F73E7B5",
    x"3F73E99E",
    x"3F73EB86",
    x"3F73ED6E",
    x"3F73EF56",
    x"3F73F13E",
    x"3F73F326",
    x"3F73F50D",
    x"3F73F6F5",
    x"3F73F8DC",
    x"3F73FAC3",
    x"3F73FCAA",
    x"3F73FE91",
    x"3F740078",
    x"3F74025F",
    x"3F740445",
    x"3F74062B",
    x"3F740812",
    x"3F7409F8",
    x"3F740BDD",
    x"3F740DC3",
    x"3F740FA9",
    x"3F74118E",
    x"3F741373",
    x"3F741558",
    x"3F74173D",
    x"3F741922",
    x"3F741B07",
    x"3F741CEB",
    x"3F741ED0",
    x"3F7420B4",
    x"3F742298",
    x"3F74247C",
    x"3F742660",
    x"3F742843",
    x"3F742A27",
    x"3F742C0A",
    x"3F742DED",
    x"3F742FD1",
    x"3F7431B3",
    x"3F743396",
    x"3F743579",
    x"3F74375B",
    x"3F74393E",
    x"3F743B20",
    x"3F743D02",
    x"3F743EE4",
    x"3F7440C5",
    x"3F7442A7",
    x"3F744488",
    x"3F74466A",
    x"3F74484B",
    x"3F744A2C",
    x"3F744C0D",
    x"3F744DED",
    x"3F744FCE",
    x"3F7451AE",
    x"3F74538F",
    x"3F74556F",
    x"3F74574F",
    x"3F74592F",
    x"3F745B0E",
    x"3F745CEE",
    x"3F745ECD",
    x"3F7460AC",
    x"3F74628B",
    x"3F74646A",
    x"3F746649",
    x"3F746828",
    x"3F746A06",
    x"3F746BE5",
    x"3F746DC3",
    x"3F746FA1",
    x"3F74717F",
    x"3F74735D",
    x"3F74753A",
    x"3F747718",
    x"3F7478F5",
    x"3F747AD2",
    x"3F747CAF",
    x"3F747E8C",
    x"3F748069",
    x"3F748245",
    x"3F748422",
    x"3F7485FE",
    x"3F7487DA",
    x"3F7489B6",
    x"3F748B92",
    x"3F748D6E",
    x"3F748F49",
    x"3F749125",
    x"3F749300",
    x"3F7494DB",
    x"3F7496B6",
    x"3F749891",
    x"3F749A6B",
    x"3F749C46",
    x"3F749E20",
    x"3F749FFA",
    x"3F74A1D5",
    x"3F74A3AE",
    x"3F74A588",
    x"3F74A762",
    x"3F74A93B",
    x"3F74AB15",
    x"3F74ACEE",
    x"3F74AEC7",
    x"3F74B0A0",
    x"3F74B279",
    x"3F74B451",
    x"3F74B62A",
    x"3F74B802",
    x"3F74B9DA",
    x"3F74BBB2",
    x"3F74BD8A",
    x"3F74BF62",
    x"3F74C139",
    x"3F74C311",
    x"3F74C4E8",
    x"3F74C6BF",
    x"3F74C896",
    x"3F74CA6D",
    x"3F74CC44",
    x"3F74CE1A",
    x"3F74CFF0",
    x"3F74D1C7",
    x"3F74D39D",
    x"3F74D573",
    x"3F74D749",
    x"3F74D91E",
    x"3F74DAF4",
    x"3F74DCC9",
    x"3F74DE9E",
    x"3F74E073",
    x"3F74E248",
    x"3F74E41D",
    x"3F74E5F2",
    x"3F74E7C6",
    x"3F74E99A",
    x"3F74EB6F",
    x"3F74ED43",
    x"3F74EF17",
    x"3F74F0EA",
    x"3F74F2BE",
    x"3F74F491",
    x"3F74F665",
    x"3F74F838",
    x"3F74FA0B",
    x"3F74FBDE",
    x"3F74FDB0",
    x"3F74FF83",
    x"3F750155",
    x"3F750327",
    x"3F7504FA",
    x"3F7506CC",
    x"3F75089D",
    x"3F750A6F",
    x"3F750C41",
    x"3F750E12",
    x"3F750FE3",
    x"3F7511B4",
    x"3F751385",
    x"3F751556",
    x"3F751727",
    x"3F7518F7",
    x"3F751AC7",
    x"3F751C98",
    x"3F751E68",
    x"3F752038",
    x"3F752207",
    x"3F7523D7",
    x"3F7525A6",
    x"3F752776",
    x"3F752945",
    x"3F752B14",
    x"3F752CE3",
    x"3F752EB1",
    x"3F753080",
    x"3F75324E",
    x"3F75341D",
    x"3F7535EB",
    x"3F7537B9",
    x"3F753987",
    x"3F753B54",
    x"3F753D22",
    x"3F753EEF",
    x"3F7540BC",
    x"3F754289",
    x"3F754456",
    x"3F754623",
    x"3F7547F0",
    x"3F7549BC",
    x"3F754B89",
    x"3F754D55",
    x"3F754F21",
    x"3F7550ED",
    x"3F7552B9",
    x"3F755484",
    x"3F755650",
    x"3F75581B",
    x"3F7559E6",
    x"3F755BB1",
    x"3F755D7C",
    x"3F755F47",
    x"3F756111",
    x"3F7562DC",
    x"3F7564A6",
    x"3F756670",
    x"3F75683A",
    x"3F756A04",
    x"3F756BCE",
    x"3F756D97",
    x"3F756F61",
    x"3F75712A",
    x"3F7572F3",
    x"3F7574BC",
    x"3F757685",
    x"3F75784D",
    x"3F757A16",
    x"3F757BDE",
    x"3F757DA7",
    x"3F757F6F",
    x"3F758136",
    x"3F7582FE",
    x"3F7584C6",
    x"3F75868D",
    x"3F758855",
    x"3F758A1C",
    x"3F758BE3",
    x"3F758DAA",
    x"3F758F70",
    x"3F759137",
    x"3F7592FE",
    x"3F7594C4",
    x"3F75968A",
    x"3F759850",
    x"3F759A16",
    x"3F759BDB",
    x"3F759DA1",
    x"3F759F66",
    x"3F75A12C",
    x"3F75A2F1",
    x"3F75A4B6",
    x"3F75A67B",
    x"3F75A83F",
    x"3F75AA04",
    x"3F75ABC8",
    x"3F75AD8C",
    x"3F75AF50",
    x"3F75B114",
    x"3F75B2D8",
    x"3F75B49C",
    x"3F75B65F",
    x"3F75B822",
    x"3F75B9E6",
    x"3F75BBA9",
    x"3F75BD6C",
    x"3F75BF2E",
    x"3F75C0F1",
    x"3F75C2B3",
    x"3F75C476",
    x"3F75C638",
    x"3F75C7FA",
    x"3F75C9BC",
    x"3F75CB7D",
    x"3F75CD3F",
    x"3F75CF00",
    x"3F75D0C2",
    x"3F75D283",
    x"3F75D444",
    x"3F75D604",
    x"3F75D7C5",
    x"3F75D986",
    x"3F75DB46",
    x"3F75DD06",
    x"3F75DEC6",
    x"3F75E086",
    x"3F75E246",
    x"3F75E406",
    x"3F75E5C5",
    x"3F75E784",
    x"3F75E944",
    x"3F75EB03",
    x"3F75ECC2",
    x"3F75EE80",
    x"3F75F03F",
    x"3F75F1FD",
    x"3F75F3BC",
    x"3F75F57A",
    x"3F75F738",
    x"3F75F8F6",
    x"3F75FAB3",
    x"3F75FC71",
    x"3F75FE2E",
    x"3F75FFEB",
    x"3F7601A9",
    x"3F760366",
    x"3F760522",
    x"3F7606DF",
    x"3F76089C",
    x"3F760A58",
    x"3F760C14",
    x"3F760DD0",
    x"3F760F8C",
    x"3F761148",
    x"3F761304",
    x"3F7614BF",
    x"3F76167A",
    x"3F761836",
    x"3F7619F1",
    x"3F761BAB",
    x"3F761D66",
    x"3F761F21",
    x"3F7620DB",
    x"3F762296",
    x"3F762450",
    x"3F76260A",
    x"3F7627C3",
    x"3F76297D",
    x"3F762B37",
    x"3F762CF0",
    x"3F762EA9",
    x"3F763063",
    x"3F76321B",
    x"3F7633D4",
    x"3F76358D",
    x"3F763745",
    x"3F7638FE",
    x"3F763AB6",
    x"3F763C6E",
    x"3F763E26",
    x"3F763FDE",
    x"3F764195",
    x"3F76434D",
    x"3F764504",
    x"3F7646BB",
    x"3F764872",
    x"3F764A29",
    x"3F764BE0",
    x"3F764D97",
    x"3F764F4D",
    x"3F765103",
    x"3F7652B9",
    x"3F76546F",
    x"3F765625",
    x"3F7657DB",
    x"3F765991",
    x"3F765B46",
    x"3F765CFB",
    x"3F765EB0",
    x"3F766065",
    x"3F76621A",
    x"3F7663CF",
    x"3F766583",
    x"3F766738",
    x"3F7668EC",
    x"3F766AA0",
    x"3F766C54",
    x"3F766E08",
    x"3F766FBB",
    x"3F76716F",
    x"3F767322",
    x"3F7674D5",
    x"3F767688",
    x"3F76783B",
    x"3F7679EE",
    x"3F767BA0",
    x"3F767D53",
    x"3F767F05",
    x"3F7680B7",
    x"3F768269",
    x"3F76841B",
    x"3F7685CD",
    x"3F76877E",
    x"3F768930",
    x"3F768AE1",
    x"3F768C92",
    x"3F768E43",
    x"3F768FF4",
    x"3F7691A4",
    x"3F769355",
    x"3F769505",
    x"3F7696B5",
    x"3F769865",
    x"3F769A15",
    x"3F769BC5",
    x"3F769D75",
    x"3F769F24",
    x"3F76A0D3",
    x"3F76A283",
    x"3F76A432",
    x"3F76A5E0",
    x"3F76A78F",
    x"3F76A93E",
    x"3F76AAEC",
    x"3F76AC9A",
    x"3F76AE49",
    x"3F76AFF7",
    x"3F76B1A4",
    x"3F76B352",
    x"3F76B500",
    x"3F76B6AD",
    x"3F76B85A",
    x"3F76BA07",
    x"3F76BBB4",
    x"3F76BD61",
    x"3F76BF0E",
    x"3F76C0BA",
    x"3F76C266",
    x"3F76C413",
    x"3F76C5BF",
    x"3F76C76B",
    x"3F76C916",
    x"3F76CAC2",
    x"3F76CC6D",
    x"3F76CE19",
    x"3F76CFC4",
    x"3F76D16F",
    x"3F76D31A",
    x"3F76D4C4",
    x"3F76D66F",
    x"3F76D819",
    x"3F76D9C4",
    x"3F76DB6E",
    x"3F76DD18",
    x"3F76DEC1",
    x"3F76E06B",
    x"3F76E215",
    x"3F76E3BE",
    x"3F76E567",
    x"3F76E710",
    x"3F76E8B9",
    x"3F76EA62",
    x"3F76EC0B",
    x"3F76EDB3",
    x"3F76EF5B",
    x"3F76F103",
    x"3F76F2AC",
    x"3F76F453",
    x"3F76F5FB",
    x"3F76F7A3",
    x"3F76F94A",
    x"3F76FAF1",
    x"3F76FC99",
    x"3F76FE40",
    x"3F76FFE6",
    x"3F77018D",
    x"3F770334",
    x"3F7704DA",
    x"3F770680",
    x"3F770826",
    x"3F7709CC",
    x"3F770B72",
    x"3F770D18",
    x"3F770EBD",
    x"3F771063",
    x"3F771208",
    x"3F7713AD",
    x"3F771552",
    x"3F7716F6",
    x"3F77189B",
    x"3F771A3F",
    x"3F771BE4",
    x"3F771D88",
    x"3F771F2C",
    x"3F7720D0",
    x"3F772274",
    x"3F772417",
    x"3F7725BA",
    x"3F77275E",
    x"3F772901",
    x"3F772AA4",
    x"3F772C47",
    x"3F772DE9",
    x"3F772F8C",
    x"3F77312E",
    x"3F7732D0",
    x"3F773472",
    x"3F773614",
    x"3F7737B6",
    x"3F773958",
    x"3F773AF9",
    x"3F773C9B",
    x"3F773E3C",
    x"3F773FDD",
    x"3F77417E",
    x"3F77431E",
    x"3F7744BF",
    x"3F77465F",
    x"3F774800",
    x"3F7749A0",
    x"3F774B40",
    x"3F774CE0",
    x"3F774E7F",
    x"3F77501F",
    x"3F7751BE",
    x"3F77535E",
    x"3F7754FD",
    x"3F77569C",
    x"3F77583A",
    x"3F7759D9",
    x"3F775B78",
    x"3F775D16",
    x"3F775EB4",
    x"3F776052",
    x"3F7761F0",
    x"3F77638E",
    x"3F77652B",
    x"3F7766C9",
    x"3F776866",
    x"3F776A03",
    x"3F776BA0",
    x"3F776D3D",
    x"3F776EDA",
    x"3F777076",
    x"3F777213",
    x"3F7773AF",
    x"3F77754B",
    x"3F7776E7",
    x"3F777883",
    x"3F777A1F",
    x"3F777BBA",
    x"3F777D56",
    x"3F777EF1",
    x"3F77808C",
    x"3F778227",
    x"3F7783C2",
    x"3F77855C",
    x"3F7786F7",
    x"3F778891",
    x"3F778A2B",
    x"3F778BC5",
    x"3F778D5F",
    x"3F778EF9",
    x"3F779092",
    x"3F77922C",
    x"3F7793C5",
    x"3F77955E",
    x"3F7796F7",
    x"3F779890",
    x"3F779A29",
    x"3F779BC1",
    x"3F779D5A",
    x"3F779EF2",
    x"3F77A08A",
    x"3F77A222",
    x"3F77A3BA",
    x"3F77A551",
    x"3F77A6E9",
    x"3F77A880",
    x"3F77AA17",
    x"3F77ABAE",
    x"3F77AD45",
    x"3F77AEDC",
    x"3F77B073",
    x"3F77B209",
    x"3F77B39F",
    x"3F77B535",
    x"3F77B6CB",
    x"3F77B861",
    x"3F77B9F7",
    x"3F77BB8D",
    x"3F77BD22",
    x"3F77BEB7",
    x"3F77C04C",
    x"3F77C1E1",
    x"3F77C376",
    x"3F77C50B",
    x"3F77C69F",
    x"3F77C834",
    x"3F77C9C8",
    x"3F77CB5C",
    x"3F77CCF0",
    x"3F77CE83",
    x"3F77D017",
    x"3F77D1AB",
    x"3F77D33E",
    x"3F77D4D1",
    x"3F77D664",
    x"3F77D7F7",
    x"3F77D98A",
    x"3F77DB1C",
    x"3F77DCAF",
    x"3F77DE41",
    x"3F77DFD3",
    x"3F77E165",
    x"3F77E2F7",
    x"3F77E488",
    x"3F77E61A",
    x"3F77E7AB",
    x"3F77E93D",
    x"3F77EACE",
    x"3F77EC5F",
    x"3F77EDEF",
    x"3F77EF80",
    x"3F77F110",
    x"3F77F2A1",
    x"3F77F431",
    x"3F77F5C1",
    x"3F77F751",
    x"3F77F8E1",
    x"3F77FA70",
    x"3F77FC00",
    x"3F77FD8F",
    x"3F77FF1E",
    x"3F7800AD",
    x"3F78023C",
    x"3F7803CA",
    x"3F780559",
    x"3F7806E7",
    x"3F780876",
    x"3F780A04",
    x"3F780B92",
    x"3F780D1F",
    x"3F780EAD",
    x"3F78103A",
    x"3F7811C8",
    x"3F781355",
    x"3F7814E2",
    x"3F78166F",
    x"3F7817FC",
    x"3F781988",
    x"3F781B15",
    x"3F781CA1",
    x"3F781E2D",
    x"3F781FB9",
    x"3F782145",
    x"3F7822D1",
    x"3F78245C",
    x"3F7825E8",
    x"3F782773",
    x"3F7828FE",
    x"3F782A89",
    x"3F782C14",
    x"3F782D9E",
    x"3F782F29",
    x"3F7830B3",
    x"3F78323D",
    x"3F7833C7",
    x"3F783551",
    x"3F7836DB",
    x"3F783865",
    x"3F7839EE",
    x"3F783B77",
    x"3F783D01",
    x"3F783E8A",
    x"3F784012",
    x"3F78419B",
    x"3F784324",
    x"3F7844AC",
    x"3F784634",
    x"3F7847BC",
    x"3F784944",
    x"3F784ACC",
    x"3F784C54",
    x"3F784DDB",
    x"3F784F63",
    x"3F7850EA",
    x"3F785271",
    x"3F7853F8",
    x"3F78557F",
    x"3F785705",
    x"3F78588C",
    x"3F785A12",
    x"3F785B98",
    x"3F785D1E",
    x"3F785EA4",
    x"3F78602A",
    x"3F7861AF",
    x"3F786335",
    x"3F7864BA",
    x"3F78663F",
    x"3F7867C4",
    x"3F786949",
    x"3F786ACE",
    x"3F786C52",
    x"3F786DD6",
    x"3F786F5B",
    x"3F7870DF",
    x"3F787263",
    x"3F7873E6",
    x"3F78756A",
    x"3F7876ED",
    x"3F787871",
    x"3F7879F4",
    x"3F787B77",
    x"3F787CFA",
    x"3F787E7D",
    x"3F787FFF",
    x"3F788182",
    x"3F788304",
    x"3F788486",
    x"3F788608",
    x"3F78878A",
    x"3F78890B",
    x"3F788A8D",
    x"3F788C0E",
    x"3F788D8F",
    x"3F788F11",
    x"3F789091",
    x"3F789212",
    x"3F789393",
    x"3F789513",
    x"3F789694",
    x"3F789814",
    x"3F789994",
    x"3F789B14",
    x"3F789C93",
    x"3F789E13",
    x"3F789F92",
    x"3F78A112",
    x"3F78A291",
    x"3F78A410",
    x"3F78A58F",
    x"3F78A70D",
    x"3F78A88C",
    x"3F78AA0A",
    x"3F78AB88",
    x"3F78AD06",
    x"3F78AE84",
    x"3F78B002",
    x"3F78B180",
    x"3F78B2FD",
    x"3F78B47B",
    x"3F78B5F8",
    x"3F78B775",
    x"3F78B8F2",
    x"3F78BA6E",
    x"3F78BBEB",
    x"3F78BD67",
    x"3F78BEE4",
    x"3F78C060",
    x"3F78C1DC",
    x"3F78C358",
    x"3F78C4D3",
    x"3F78C64F",
    x"3F78C7CA",
    x"3F78C945",
    x"3F78CAC1",
    x"3F78CC3B",
    x"3F78CDB6",
    x"3F78CF31",
    x"3F78D0AB",
    x"3F78D226",
    x"3F78D3A0",
    x"3F78D51A",
    x"3F78D694",
    x"3F78D80E",
    x"3F78D987",
    x"3F78DB01",
    x"3F78DC7A",
    x"3F78DDF3",
    x"3F78DF6C",
    x"3F78E0E5",
    x"3F78E25D",
    x"3F78E3D6",
    x"3F78E54E",
    x"3F78E6C7",
    x"3F78E83F",
    x"3F78E9B7",
    x"3F78EB2E",
    x"3F78ECA6",
    x"3F78EE1D",
    x"3F78EF95",
    x"3F78F10C",
    x"3F78F283",
    x"3F78F3FA",
    x"3F78F571",
    x"3F78F6E7",
    x"3F78F85E",
    x"3F78F9D4",
    x"3F78FB4A",
    x"3F78FCC0",
    x"3F78FE36",
    x"3F78FFAC",
    x"3F790121",
    x"3F790296",
    x"3F79040C",
    x"3F790581",
    x"3F7906F6",
    x"3F79086A",
    x"3F7909DF",
    x"3F790B54",
    x"3F790CC8",
    x"3F790E3C",
    x"3F790FB0",
    x"3F791124",
    x"3F791298",
    x"3F79140B",
    x"3F79157F",
    x"3F7916F2",
    x"3F791865",
    x"3F7919D8",
    x"3F791B4B",
    x"3F791CBE",
    x"3F791E30",
    x"3F791FA3",
    x"3F792115",
    x"3F792287",
    x"3F7923F9",
    x"3F79256B",
    x"3F7926DC",
    x"3F79284E",
    x"3F7929BF",
    x"3F792B30",
    x"3F792CA1",
    x"3F792E12",
    x"3F792F83",
    x"3F7930F3",
    x"3F793264",
    x"3F7933D4",
    x"3F793544",
    x"3F7936B4",
    x"3F793824",
    x"3F793994",
    x"3F793B03",
    x"3F793C73",
    x"3F793DE2",
    x"3F793F51",
    x"3F7940C0",
    x"3F79422F",
    x"3F79439D",
    x"3F79450C",
    x"3F79467A",
    x"3F7947E8",
    x"3F794956",
    x"3F794AC4",
    x"3F794C32",
    x"3F794D9F",
    x"3F794F0D",
    x"3F79507A",
    x"3F7951E7",
    x"3F795354",
    x"3F7954C1",
    x"3F79562E",
    x"3F79579A",
    x"3F795907",
    x"3F795A73",
    x"3F795BDF",
    x"3F795D4B",
    x"3F795EB7",
    x"3F796022",
    x"3F79618E",
    x"3F7962F9",
    x"3F796464",
    x"3F7965CF",
    x"3F79673A",
    x"3F7968A5",
    x"3F796A0F",
    x"3F796B7A",
    x"3F796CE4",
    x"3F796E4E",
    x"3F796FB8",
    x"3F797122",
    x"3F79728C",
    x"3F7973F5",
    x"3F79755F",
    x"3F7976C8",
    x"3F797831",
    x"3F79799A",
    x"3F797B03",
    x"3F797C6B",
    x"3F797DD4",
    x"3F797F3C",
    x"3F7980A4",
    x"3F79820C",
    x"3F798374",
    x"3F7984DC",
    x"3F798643",
    x"3F7987AB",
    x"3F798912",
    x"3F798A79",
    x"3F798BE0",
    x"3F798D47",
    x"3F798EAE",
    x"3F799014",
    x"3F79917A",
    x"3F7992E1",
    x"3F799447",
    x"3F7995AD",
    x"3F799712",
    x"3F799878",
    x"3F7999DE",
    x"3F799B43",
    x"3F799CA8",
    x"3F799E0D",
    x"3F799F72",
    x"3F79A0D7",
    x"3F79A23B",
    x"3F79A3A0",
    x"3F79A504",
    x"3F79A668",
    x"3F79A7CC",
    x"3F79A930",
    x"3F79AA93",
    x"3F79ABF7",
    x"3F79AD5A",
    x"3F79AEBD",
    x"3F79B020",
    x"3F79B183",
    x"3F79B2E6",
    x"3F79B449",
    x"3F79B5AB",
    x"3F79B70D",
    x"3F79B870",
    x"3F79B9D2",
    x"3F79BB33",
    x"3F79BC95",
    x"3F79BDF7",
    x"3F79BF58",
    x"3F79C0B9",
    x"3F79C21A",
    x"3F79C37B",
    x"3F79C4DC",
    x"3F79C63D",
    x"3F79C79D",
    x"3F79C8FE",
    x"3F79CA5E",
    x"3F79CBBE",
    x"3F79CD1E",
    x"3F79CE7E",
    x"3F79CFDD",
    x"3F79D13D",
    x"3F79D29C",
    x"3F79D3FB",
    x"3F79D55A",
    x"3F79D6B9",
    x"3F79D818",
    x"3F79D976",
    x"3F79DAD5",
    x"3F79DC33",
    x"3F79DD91",
    x"3F79DEEF",
    x"3F79E04D",
    x"3F79E1AA",
    x"3F79E308",
    x"3F79E465",
    x"3F79E5C2",
    x"3F79E71F",
    x"3F79E87C",
    x"3F79E9D9",
    x"3F79EB36",
    x"3F79EC92",
    x"3F79EDEE",
    x"3F79EF4A",
    x"3F79F0A6",
    x"3F79F202",
    x"3F79F35E",
    x"3F79F4B9",
    x"3F79F615",
    x"3F79F770",
    x"3F79F8CB",
    x"3F79FA26",
    x"3F79FB81",
    x"3F79FCDB",
    x"3F79FE36",
    x"3F79FF90",
    x"3F7A00EA",
    x"3F7A0244",
    x"3F7A039E",
    x"3F7A04F8",
    x"3F7A0652",
    x"3F7A07AB",
    x"3F7A0904",
    x"3F7A0A5D",
    x"3F7A0BB6",
    x"3F7A0D0F",
    x"3F7A0E68",
    x"3F7A0FC0",
    x"3F7A1119",
    x"3F7A1271",
    x"3F7A13C9",
    x"3F7A1521",
    x"3F7A1679",
    x"3F7A17D0",
    x"3F7A1928",
    x"3F7A1A7F",
    x"3F7A1BD6",
    x"3F7A1D2D",
    x"3F7A1E84",
    x"3F7A1FDB",
    x"3F7A2131",
    x"3F7A2288",
    x"3F7A23DE",
    x"3F7A2534",
    x"3F7A268A",
    x"3F7A27E0",
    x"3F7A2936",
    x"3F7A2A8B",
    x"3F7A2BE1",
    x"3F7A2D36",
    x"3F7A2E8B",
    x"3F7A2FE0",
    x"3F7A3134",
    x"3F7A3289",
    x"3F7A33DD",
    x"3F7A3532",
    x"3F7A3686",
    x"3F7A37DA",
    x"3F7A392E",
    x"3F7A3A81",
    x"3F7A3BD5",
    x"3F7A3D28",
    x"3F7A3E7C",
    x"3F7A3FCF",
    x"3F7A4122",
    x"3F7A4275",
    x"3F7A43C7",
    x"3F7A451A",
    x"3F7A466C",
    x"3F7A47BE",
    x"3F7A4910",
    x"3F7A4A62",
    x"3F7A4BB4",
    x"3F7A4D05",
    x"3F7A4E57",
    x"3F7A4FA8",
    x"3F7A50F9",
    x"3F7A524A",
    x"3F7A539B",
    x"3F7A54EC",
    x"3F7A563C",
    x"3F7A578D",
    x"3F7A58DD",
    x"3F7A5A2D",
    x"3F7A5B7D",
    x"3F7A5CCD",
    x"3F7A5E1C",
    x"3F7A5F6C",
    x"3F7A60BB",
    x"3F7A620A",
    x"3F7A6359",
    x"3F7A64A8",
    x"3F7A65F7",
    x"3F7A6745",
    x"3F7A6894",
    x"3F7A69E2",
    x"3F7A6B30",
    x"3F7A6C7E",
    x"3F7A6DCC",
    x"3F7A6F1A",
    x"3F7A7067",
    x"3F7A71B5",
    x"3F7A7302",
    x"3F7A744F",
    x"3F7A759C",
    x"3F7A76E9",
    x"3F7A7835",
    x"3F7A7982",
    x"3F7A7ACE",
    x"3F7A7C1A",
    x"3F7A7D66",
    x"3F7A7EB2",
    x"3F7A7FFE",
    x"3F7A8149",
    x"3F7A8295",
    x"3F7A83E0",
    x"3F7A852B",
    x"3F7A8676",
    x"3F7A87C1",
    x"3F7A890B",
    x"3F7A8A56",
    x"3F7A8BA0",
    x"3F7A8CEA",
    x"3F7A8E34",
    x"3F7A8F7E",
    x"3F7A90C8",
    x"3F7A9212",
    x"3F7A935B",
    x"3F7A94A4",
    x"3F7A95EE",
    x"3F7A9737",
    x"3F7A987F",
    x"3F7A99C8",
    x"3F7A9B11",
    x"3F7A9C59",
    x"3F7A9DA1",
    x"3F7A9EE9",
    x"3F7AA031",
    x"3F7AA179",
    x"3F7AA2C1",
    x"3F7AA408",
    x"3F7AA54F",
    x"3F7AA697",
    x"3F7AA7DE",
    x"3F7AA925",
    x"3F7AAA6B",
    x"3F7AABB2",
    x"3F7AACF8",
    x"3F7AAE3F",
    x"3F7AAF85",
    x"3F7AB0CB",
    x"3F7AB210",
    x"3F7AB356",
    x"3F7AB49C",
    x"3F7AB5E1",
    x"3F7AB726",
    x"3F7AB86B",
    x"3F7AB9B0",
    x"3F7ABAF5",
    x"3F7ABC3A",
    x"3F7ABD7E",
    x"3F7ABEC2",
    x"3F7AC006",
    x"3F7AC14A",
    x"3F7AC28E",
    x"3F7AC3D2",
    x"3F7AC516",
    x"3F7AC659",
    x"3F7AC79C",
    x"3F7AC8DF",
    x"3F7ACA22",
    x"3F7ACB65",
    x"3F7ACCA8",
    x"3F7ACDEA",
    x"3F7ACF2D",
    x"3F7AD06F",
    x"3F7AD1B1",
    x"3F7AD2F3",
    x"3F7AD434",
    x"3F7AD576",
    x"3F7AD6B7",
    x"3F7AD7F9",
    x"3F7AD93A",
    x"3F7ADA7B",
    x"3F7ADBBC",
    x"3F7ADCFC",
    x"3F7ADE3D",
    x"3F7ADF7D",
    x"3F7AE0BD",
    x"3F7AE1FE",
    x"3F7AE33D",
    x"3F7AE47D",
    x"3F7AE5BD",
    x"3F7AE6FC",
    x"3F7AE83C",
    x"3F7AE97B",
    x"3F7AEABA",
    x"3F7AEBF9",
    x"3F7AED37",
    x"3F7AEE76",
    x"3F7AEFB4",
    x"3F7AF0F3",
    x"3F7AF231",
    x"3F7AF36F",
    x"3F7AF4AD",
    x"3F7AF5EA",
    x"3F7AF728",
    x"3F7AF865",
    x"3F7AF9A2",
    x"3F7AFADF",
    x"3F7AFC1C",
    x"3F7AFD59",
    x"3F7AFE96",
    x"3F7AFFD2",
    x"3F7B010E",
    x"3F7B024A",
    x"3F7B0386",
    x"3F7B04C2",
    x"3F7B05FE",
    x"3F7B073A",
    x"3F7B0875",
    x"3F7B09B0",
    x"3F7B0AEB",
    x"3F7B0C26",
    x"3F7B0D61",
    x"3F7B0E9C",
    x"3F7B0FD6",
    x"3F7B1110",
    x"3F7B124B",
    x"3F7B1385",
    x"3F7B14BE",
    x"3F7B15F8",
    x"3F7B1732",
    x"3F7B186B",
    x"3F7B19A4",
    x"3F7B1ADE",
    x"3F7B1C17",
    x"3F7B1D4F",
    x"3F7B1E88",
    x"3F7B1FC1",
    x"3F7B20F9",
    x"3F7B2231",
    x"3F7B2369",
    x"3F7B24A1",
    x"3F7B25D9",
    x"3F7B2711",
    x"3F7B2848",
    x"3F7B297F",
    x"3F7B2AB6",
    x"3F7B2BED",
    x"3F7B2D24",
    x"3F7B2E5B",
    x"3F7B2F92",
    x"3F7B30C8",
    x"3F7B31FE",
    x"3F7B3334",
    x"3F7B346A",
    x"3F7B35A0",
    x"3F7B36D6",
    x"3F7B380B",
    x"3F7B3940",
    x"3F7B3A76",
    x"3F7B3BAB",
    x"3F7B3CE0",
    x"3F7B3E14",
    x"3F7B3F49",
    x"3F7B407D",
    x"3F7B41B2",
    x"3F7B42E6",
    x"3F7B441A",
    x"3F7B454E",
    x"3F7B4681",
    x"3F7B47B5",
    x"3F7B48E8",
    x"3F7B4A1B",
    x"3F7B4B4E",
    x"3F7B4C81",
    x"3F7B4DB4",
    x"3F7B4EE7",
    x"3F7B5019",
    x"3F7B514B",
    x"3F7B527E",
    x"3F7B53B0",
    x"3F7B54E1",
    x"3F7B5613",
    x"3F7B5745",
    x"3F7B5876",
    x"3F7B59A7",
    x"3F7B5AD9",
    x"3F7B5C09",
    x"3F7B5D3A",
    x"3F7B5E6B",
    x"3F7B5F9B",
    x"3F7B60CC",
    x"3F7B61FC",
    x"3F7B632C",
    x"3F7B645C",
    x"3F7B658C",
    x"3F7B66BB",
    x"3F7B67EB",
    x"3F7B691A",
    x"3F7B6A49",
    x"3F7B6B78",
    x"3F7B6CA7",
    x"3F7B6DD6",
    x"3F7B6F04",
    x"3F7B7032",
    x"3F7B7161",
    x"3F7B728F",
    x"3F7B73BD",
    x"3F7B74EA",
    x"3F7B7618",
    x"3F7B7745",
    x"3F7B7873",
    x"3F7B79A0",
    x"3F7B7ACD",
    x"3F7B7BFA",
    x"3F7B7D27",
    x"3F7B7E53",
    x"3F7B7F80",
    x"3F7B80AC",
    x"3F7B81D8",
    x"3F7B8304",
    x"3F7B8430",
    x"3F7B855B",
    x"3F7B8687",
    x"3F7B87B2",
    x"3F7B88DD",
    x"3F7B8A08",
    x"3F7B8B33",
    x"3F7B8C5E",
    x"3F7B8D89",
    x"3F7B8EB3",
    x"3F7B8FDD",
    x"3F7B9107",
    x"3F7B9231",
    x"3F7B935B",
    x"3F7B9485",
    x"3F7B95AE",
    x"3F7B96D8",
    x"3F7B9801",
    x"3F7B992A",
    x"3F7B9A53",
    x"3F7B9B7C",
    x"3F7B9CA4",
    x"3F7B9DCD",
    x"3F7B9EF5",
    x"3F7BA01D",
    x"3F7BA145",
    x"3F7BA26D",
    x"3F7BA395",
    x"3F7BA4BC",
    x"3F7BA5E4",
    x"3F7BA70B",
    x"3F7BA832",
    x"3F7BA959",
    x"3F7BAA80",
    x"3F7BABA7",
    x"3F7BACCD",
    x"3F7BADF3",
    x"3F7BAF1A",
    x"3F7BB040",
    x"3F7BB166",
    x"3F7BB28B",
    x"3F7BB3B1",
    x"3F7BB4D6",
    x"3F7BB5FC",
    x"3F7BB721",
    x"3F7BB846",
    x"3F7BB96B",
    x"3F7BBA8F",
    x"3F7BBBB4",
    x"3F7BBCD8",
    x"3F7BBDFC",
    x"3F7BBF20",
    x"3F7BC044",
    x"3F7BC168",
    x"3F7BC28C",
    x"3F7BC3AF",
    x"3F7BC4D2",
    x"3F7BC5F6",
    x"3F7BC719",
    x"3F7BC83B",
    x"3F7BC95E",
    x"3F7BCA81",
    x"3F7BCBA3",
    x"3F7BCCC5",
    x"3F7BCDE7",
    x"3F7BCF09",
    x"3F7BD02B",
    x"3F7BD14D",
    x"3F7BD26E",
    x"3F7BD390",
    x"3F7BD4B1",
    x"3F7BD5D2",
    x"3F7BD6F3",
    x"3F7BD814",
    x"3F7BD934",
    x"3F7BDA55",
    x"3F7BDB75",
    x"3F7BDC95",
    x"3F7BDDB5",
    x"3F7BDED5",
    x"3F7BDFF4",
    x"3F7BE114",
    x"3F7BE233",
    x"3F7BE353",
    x"3F7BE472",
    x"3F7BE590",
    x"3F7BE6AF",
    x"3F7BE7CE",
    x"3F7BE8EC",
    x"3F7BEA0B",
    x"3F7BEB29",
    x"3F7BEC47",
    x"3F7BED65",
    x"3F7BEE82",
    x"3F7BEFA0",
    x"3F7BF0BD",
    x"3F7BF1DA",
    x"3F7BF2F8",
    x"3F7BF415",
    x"3F7BF531",
    x"3F7BF64E",
    x"3F7BF76A",
    x"3F7BF887",
    x"3F7BF9A3",
    x"3F7BFABF",
    x"3F7BFBDB",
    x"3F7BFCF7",
    x"3F7BFE12",
    x"3F7BFF2E",
    x"3F7C0049",
    x"3F7C0164",
    x"3F7C027F",
    x"3F7C039A",
    x"3F7C04B4",
    x"3F7C05CF",
    x"3F7C06E9",
    x"3F7C0803",
    x"3F7C091E",
    x"3F7C0A37",
    x"3F7C0B51",
    x"3F7C0C6B",
    x"3F7C0D84",
    x"3F7C0E9D",
    x"3F7C0FB7",
    x"3F7C10D0",
    x"3F7C11E8",
    x"3F7C1301",
    x"3F7C141A",
    x"3F7C1532",
    x"3F7C164A",
    x"3F7C1762",
    x"3F7C187A",
    x"3F7C1992",
    x"3F7C1AAA",
    x"3F7C1BC1",
    x"3F7C1CD9",
    x"3F7C1DF0",
    x"3F7C1F07",
    x"3F7C201E",
    x"3F7C2134",
    x"3F7C224B",
    x"3F7C2361",
    x"3F7C2478",
    x"3F7C258E",
    x"3F7C26A4",
    x"3F7C27B9",
    x"3F7C28CF",
    x"3F7C29E5",
    x"3F7C2AFA",
    x"3F7C2C0F",
    x"3F7C2D24",
    x"3F7C2E39",
    x"3F7C2F4E",
    x"3F7C3062",
    x"3F7C3177",
    x"3F7C328B",
    x"3F7C339F",
    x"3F7C34B3",
    x"3F7C35C7",
    x"3F7C36DB",
    x"3F7C37EE",
    x"3F7C3902",
    x"3F7C3A15",
    x"3F7C3B28",
    x"3F7C3C3B",
    x"3F7C3D4E",
    x"3F7C3E60",
    x"3F7C3F73",
    x"3F7C4085",
    x"3F7C4197",
    x"3F7C42A9",
    x"3F7C43BB",
    x"3F7C44CD",
    x"3F7C45DE",
    x"3F7C46F0",
    x"3F7C4801",
    x"3F7C4912",
    x"3F7C4A23",
    x"3F7C4B34",
    x"3F7C4C44",
    x"3F7C4D55",
    x"3F7C4E65",
    x"3F7C4F75",
    x"3F7C5085",
    x"3F7C5195",
    x"3F7C52A5",
    x"3F7C53B4",
    x"3F7C54C4",
    x"3F7C55D3",
    x"3F7C56E2",
    x"3F7C57F1",
    x"3F7C5900",
    x"3F7C5A0F",
    x"3F7C5B1D",
    x"3F7C5C2C",
    x"3F7C5D3A",
    x"3F7C5E48",
    x"3F7C5F56",
    x"3F7C6063",
    x"3F7C6171",
    x"3F7C627E",
    x"3F7C638C",
    x"3F7C6499",
    x"3F7C65A6",
    x"3F7C66B3",
    x"3F7C67BF",
    x"3F7C68CC",
    x"3F7C69D8",
    x"3F7C6AE5",
    x"3F7C6BF1",
    x"3F7C6CFD",
    x"3F7C6E08",
    x"3F7C6F14",
    x"3F7C701F",
    x"3F7C712B",
    x"3F7C7236",
    x"3F7C7341",
    x"3F7C744C",
    x"3F7C7556",
    x"3F7C7661",
    x"3F7C776B",
    x"3F7C7876",
    x"3F7C7980",
    x"3F7C7A8A",
    x"3F7C7B94",
    x"3F7C7C9D",
    x"3F7C7DA7",
    x"3F7C7EB0",
    x"3F7C7FB9",
    x"3F7C80C2",
    x"3F7C81CB",
    x"3F7C82D4",
    x"3F7C83DC",
    x"3F7C84E5",
    x"3F7C85ED",
    x"3F7C86F5",
    x"3F7C87FD",
    x"3F7C8905",
    x"3F7C8A0D",
    x"3F7C8B14",
    x"3F7C8C1C",
    x"3F7C8D23",
    x"3F7C8E2A",
    x"3F7C8F31",
    x"3F7C9037",
    x"3F7C913E",
    x"3F7C9245",
    x"3F7C934B",
    x"3F7C9451",
    x"3F7C9557",
    x"3F7C965D",
    x"3F7C9762",
    x"3F7C9868",
    x"3F7C996D",
    x"3F7C9A73",
    x"3F7C9B78",
    x"3F7C9C7D",
    x"3F7C9D81",
    x"3F7C9E86",
    x"3F7C9F8A",
    x"3F7CA08F",
    x"3F7CA193",
    x"3F7CA297",
    x"3F7CA39B",
    x"3F7CA49F",
    x"3F7CA5A2",
    x"3F7CA6A6",
    x"3F7CA7A9",
    x"3F7CA8AC",
    x"3F7CA9AF",
    x"3F7CAAB2",
    x"3F7CABB4",
    x"3F7CACB7",
    x"3F7CADB9",
    x"3F7CAEBB",
    x"3F7CAFBD",
    x"3F7CB0BF",
    x"3F7CB1C1",
    x"3F7CB2C2",
    x"3F7CB3C4",
    x"3F7CB4C5",
    x"3F7CB5C6",
    x"3F7CB6C7",
    x"3F7CB7C8",
    x"3F7CB8C9",
    x"3F7CB9C9",
    x"3F7CBACA",
    x"3F7CBBCA",
    x"3F7CBCCA",
    x"3F7CBDCA",
    x"3F7CBECA",
    x"3F7CBFC9",
    x"3F7CC0C9",
    x"3F7CC1C8",
    x"3F7CC2C7",
    x"3F7CC3C6",
    x"3F7CC4C5",
    x"3F7CC5C4",
    x"3F7CC6C2",
    x"3F7CC7C0",
    x"3F7CC8BF",
    x"3F7CC9BD",
    x"3F7CCABB",
    x"3F7CCBB8",
    x"3F7CCCB6",
    x"3F7CCDB4",
    x"3F7CCEB1",
    x"3F7CCFAE",
    x"3F7CD0AB",
    x"3F7CD1A8",
    x"3F7CD2A5",
    x"3F7CD3A1",
    x"3F7CD49E",
    x"3F7CD59A",
    x"3F7CD696",
    x"3F7CD792",
    x"3F7CD88E",
    x"3F7CD989",
    x"3F7CDA85",
    x"3F7CDB80",
    x"3F7CDC7B",
    x"3F7CDD76",
    x"3F7CDE71",
    x"3F7CDF6C",
    x"3F7CE066",
    x"3F7CE161",
    x"3F7CE25B",
    x"3F7CE355",
    x"3F7CE44F",
    x"3F7CE549",
    x"3F7CE643",
    x"3F7CE73C",
    x"3F7CE836",
    x"3F7CE92F",
    x"3F7CEA28",
    x"3F7CEB21",
    x"3F7CEC19",
    x"3F7CED12",
    x"3F7CEE0B",
    x"3F7CEF03",
    x"3F7CEFFB",
    x"3F7CF0F3",
    x"3F7CF1EB",
    x"3F7CF2E2",
    x"3F7CF3DA",
    x"3F7CF4D1",
    x"3F7CF5C9",
    x"3F7CF6C0",
    x"3F7CF7B7",
    x"3F7CF8AD",
    x"3F7CF9A4",
    x"3F7CFA9A",
    x"3F7CFB91",
    x"3F7CFC87",
    x"3F7CFD7D",
    x"3F7CFE73",
    x"3F7CFF68",
    x"3F7D005E",
    x"3F7D0153",
    x"3F7D0249",
    x"3F7D033E",
    x"3F7D0433",
    x"3F7D0527",
    x"3F7D061C",
    x"3F7D0710",
    x"3F7D0805",
    x"3F7D08F9",
    x"3F7D09ED",
    x"3F7D0AE1",
    x"3F7D0BD5",
    x"3F7D0CC8",
    x"3F7D0DBC",
    x"3F7D0EAF",
    x"3F7D0FA2",
    x"3F7D1095",
    x"3F7D1188",
    x"3F7D127A",
    x"3F7D136D",
    x"3F7D145F",
    x"3F7D1551",
    x"3F7D1643",
    x"3F7D1735",
    x"3F7D1827",
    x"3F7D1919",
    x"3F7D1A0A",
    x"3F7D1AFB",
    x"3F7D1BEC",
    x"3F7D1CDD",
    x"3F7D1DCE",
    x"3F7D1EBF",
    x"3F7D1FAF",
    x"3F7D20A0",
    x"3F7D2190",
    x"3F7D2280",
    x"3F7D2370",
    x"3F7D2460",
    x"3F7D254F",
    x"3F7D263F",
    x"3F7D272E",
    x"3F7D281D",
    x"3F7D290C",
    x"3F7D29FB",
    x"3F7D2AEA",
    x"3F7D2BD8",
    x"3F7D2CC7",
    x"3F7D2DB5",
    x"3F7D2EA3",
    x"3F7D2F91",
    x"3F7D307F",
    x"3F7D316C",
    x"3F7D325A",
    x"3F7D3347",
    x"3F7D3434",
    x"3F7D3521",
    x"3F7D360E",
    x"3F7D36FB",
    x"3F7D37E7",
    x"3F7D38D4",
    x"3F7D39C0",
    x"3F7D3AAC",
    x"3F7D3B98",
    x"3F7D3C84",
    x"3F7D3D6F",
    x"3F7D3E5B",
    x"3F7D3F46",
    x"3F7D4031",
    x"3F7D411C",
    x"3F7D4207",
    x"3F7D42F2",
    x"3F7D43DC",
    x"3F7D44C7",
    x"3F7D45B1",
    x"3F7D469B",
    x"3F7D4785",
    x"3F7D486F",
    x"3F7D4959",
    x"3F7D4A42",
    x"3F7D4B2C",
    x"3F7D4C15",
    x"3F7D4CFE",
    x"3F7D4DE7",
    x"3F7D4ECF",
    x"3F7D4FB8",
    x"3F7D50A0",
    x"3F7D5189",
    x"3F7D5271",
    x"3F7D5359",
    x"3F7D5441",
    x"3F7D5528",
    x"3F7D5610",
    x"3F7D56F7",
    x"3F7D57DE",
    x"3F7D58C5",
    x"3F7D59AC",
    x"3F7D5A93",
    x"3F7D5B7A",
    x"3F7D5C60",
    x"3F7D5D46",
    x"3F7D5E2D",
    x"3F7D5F13",
    x"3F7D5FF8",
    x"3F7D60DE",
    x"3F7D61C4",
    x"3F7D62A9",
    x"3F7D638E",
    x"3F7D6473",
    x"3F7D6558",
    x"3F7D663D",
    x"3F7D6722",
    x"3F7D6806",
    x"3F7D68EA",
    x"3F7D69CE",
    x"3F7D6AB2",
    x"3F7D6B96",
    x"3F7D6C7A",
    x"3F7D6D5E",
    x"3F7D6E41",
    x"3F7D6F24",
    x"3F7D7007",
    x"3F7D70EA",
    x"3F7D71CD",
    x"3F7D72B0",
    x"3F7D7392",
    x"3F7D7474",
    x"3F7D7557",
    x"3F7D7639",
    x"3F7D771B",
    x"3F7D77FC",
    x"3F7D78DE",
    x"3F7D79BF",
    x"3F7D7AA0",
    x"3F7D7B82",
    x"3F7D7C62",
    x"3F7D7D43",
    x"3F7D7E24",
    x"3F7D7F04",
    x"3F7D7FE5",
    x"3F7D80C5",
    x"3F7D81A5",
    x"3F7D8285",
    x"3F7D8365",
    x"3F7D8444",
    x"3F7D8524",
    x"3F7D8603",
    x"3F7D86E2",
    x"3F7D87C1",
    x"3F7D88A0",
    x"3F7D897E",
    x"3F7D8A5D",
    x"3F7D8B3B",
    x"3F7D8C19",
    x"3F7D8CF8",
    x"3F7D8DD5",
    x"3F7D8EB3",
    x"3F7D8F91",
    x"3F7D906E",
    x"3F7D914B",
    x"3F7D9229",
    x"3F7D9306",
    x"3F7D93E2",
    x"3F7D94BF",
    x"3F7D959C",
    x"3F7D9678",
    x"3F7D9754",
    x"3F7D9830",
    x"3F7D990C",
    x"3F7D99E8",
    x"3F7D9AC4",
    x"3F7D9B9F",
    x"3F7D9C7A",
    x"3F7D9D55",
    x"3F7D9E30",
    x"3F7D9F0B",
    x"3F7D9FE6",
    x"3F7DA0C0",
    x"3F7DA19B",
    x"3F7DA275",
    x"3F7DA34F",
    x"3F7DA429",
    x"3F7DA503",
    x"3F7DA5DC",
    x"3F7DA6B6",
    x"3F7DA78F",
    x"3F7DA868",
    x"3F7DA941",
    x"3F7DAA1A",
    x"3F7DAAF3",
    x"3F7DABCC",
    x"3F7DACA4",
    x"3F7DAD7C",
    x"3F7DAE54",
    x"3F7DAF2C",
    x"3F7DB004",
    x"3F7DB0DC",
    x"3F7DB1B3",
    x"3F7DB28A",
    x"3F7DB362",
    x"3F7DB439",
    x"3F7DB510",
    x"3F7DB5E6",
    x"3F7DB6BD",
    x"3F7DB793",
    x"3F7DB869",
    x"3F7DB940",
    x"3F7DBA15",
    x"3F7DBAEB",
    x"3F7DBBC1",
    x"3F7DBC96",
    x"3F7DBD6C",
    x"3F7DBE41",
    x"3F7DBF16",
    x"3F7DBFEB",
    x"3F7DC0C0",
    x"3F7DC194",
    x"3F7DC269",
    x"3F7DC33D",
    x"3F7DC411",
    x"3F7DC4E5",
    x"3F7DC5B9",
    x"3F7DC68C",
    x"3F7DC760",
    x"3F7DC833",
    x"3F7DC906",
    x"3F7DC9DA",
    x"3F7DCAAC",
    x"3F7DCB7F",
    x"3F7DCC52",
    x"3F7DCD24",
    x"3F7DCDF6",
    x"3F7DCEC9",
    x"3F7DCF9B",
    x"3F7DD06C",
    x"3F7DD13E",
    x"3F7DD210",
    x"3F7DD2E1",
    x"3F7DD3B2",
    x"3F7DD483",
    x"3F7DD554",
    x"3F7DD625",
    x"3F7DD6F5",
    x"3F7DD7C6",
    x"3F7DD896",
    x"3F7DD966",
    x"3F7DDA36",
    x"3F7DDB06",
    x"3F7DDBD6",
    x"3F7DDCA5",
    x"3F7DDD75",
    x"3F7DDE44",
    x"3F7DDF13",
    x"3F7DDFE2",
    x"3F7DE0B1",
    x"3F7DE17F",
    x"3F7DE24E",
    x"3F7DE31C",
    x"3F7DE3EA",
    x"3F7DE4B8",
    x"3F7DE586",
    x"3F7DE654",
    x"3F7DE721",
    x"3F7DE7EF",
    x"3F7DE8BC",
    x"3F7DE989",
    x"3F7DEA56",
    x"3F7DEB23",
    x"3F7DEBEF",
    x"3F7DECBC",
    x"3F7DED88",
    x"3F7DEE54",
    x"3F7DEF20",
    x"3F7DEFEC",
    x"3F7DF0B8",
    x"3F7DF183",
    x"3F7DF24F",
    x"3F7DF31A",
    x"3F7DF3E5",
    x"3F7DF4B0",
    x"3F7DF57B",
    x"3F7DF646",
    x"3F7DF710",
    x"3F7DF7DA",
    x"3F7DF8A5",
    x"3F7DF96F",
    x"3F7DFA38",
    x"3F7DFB02",
    x"3F7DFBCC",
    x"3F7DFC95",
    x"3F7DFD5E",
    x"3F7DFE28",
    x"3F7DFEF0",
    x"3F7DFFB9",
    x"3F7E0082",
    x"3F7E014A",
    x"3F7E0213",
    x"3F7E02DB",
    x"3F7E03A3",
    x"3F7E046B",
    x"3F7E0533",
    x"3F7E05FA",
    x"3F7E06C2",
    x"3F7E0789",
    x"3F7E0850",
    x"3F7E0917",
    x"3F7E09DE",
    x"3F7E0AA4",
    x"3F7E0B6B",
    x"3F7E0C31",
    x"3F7E0CF7",
    x"3F7E0DBD",
    x"3F7E0E83",
    x"3F7E0F49",
    x"3F7E100F",
    x"3F7E10D4",
    x"3F7E1199",
    x"3F7E125F",
    x"3F7E1324",
    x"3F7E13E8",
    x"3F7E14AD",
    x"3F7E1572",
    x"3F7E1636",
    x"3F7E16FA",
    x"3F7E17BE",
    x"3F7E1882",
    x"3F7E1946",
    x"3F7E1A09",
    x"3F7E1ACD",
    x"3F7E1B90",
    x"3F7E1C53",
    x"3F7E1D16",
    x"3F7E1DD9",
    x"3F7E1E9C",
    x"3F7E1F5E",
    x"3F7E2021",
    x"3F7E20E3",
    x"3F7E21A5",
    x"3F7E2267",
    x"3F7E2329",
    x"3F7E23EA",
    x"3F7E24AC",
    x"3F7E256D",
    x"3F7E262E",
    x"3F7E26EF",
    x"3F7E27B0",
    x"3F7E2871",
    x"3F7E2931",
    x"3F7E29F2",
    x"3F7E2AB2",
    x"3F7E2B72",
    x"3F7E2C32",
    x"3F7E2CF2",
    x"3F7E2DB1",
    x"3F7E2E71",
    x"3F7E2F30",
    x"3F7E2FEF",
    x"3F7E30AE",
    x"3F7E316D",
    x"3F7E322C",
    x"3F7E32EA",
    x"3F7E33A9",
    x"3F7E3467",
    x"3F7E3525",
    x"3F7E35E3",
    x"3F7E36A1",
    x"3F7E375E",
    x"3F7E381C",
    x"3F7E38D9",
    x"3F7E3996",
    x"3F7E3A53",
    x"3F7E3B10",
    x"3F7E3BCD",
    x"3F7E3C89",
    x"3F7E3D46",
    x"3F7E3E02",
    x"3F7E3EBE",
    x"3F7E3F7A",
    x"3F7E4036",
    x"3F7E40F1",
    x"3F7E41AD",
    x"3F7E4268",
    x"3F7E4323",
    x"3F7E43DE",
    x"3F7E4499",
    x"3F7E4554",
    x"3F7E460F",
    x"3F7E46C9",
    x"3F7E4783",
    x"3F7E483D",
    x"3F7E48F7",
    x"3F7E49B1",
    x"3F7E4A6B",
    x"3F7E4B24",
    x"3F7E4BDE",
    x"3F7E4C97",
    x"3F7E4D50",
    x"3F7E4E09",
    x"3F7E4EC1",
    x"3F7E4F7A",
    x"3F7E5032",
    x"3F7E50EB",
    x"3F7E51A3",
    x"3F7E525B",
    x"3F7E5312",
    x"3F7E53CA",
    x"3F7E5482",
    x"3F7E5539",
    x"3F7E55F0",
    x"3F7E56A7",
    x"3F7E575E",
    x"3F7E5815",
    x"3F7E58CB",
    x"3F7E5982",
    x"3F7E5A38",
    x"3F7E5AEE",
    x"3F7E5BA4",
    x"3F7E5C5A",
    x"3F7E5D10",
    x"3F7E5DC5",
    x"3F7E5E7B",
    x"3F7E5F30",
    x"3F7E5FE5",
    x"3F7E609A",
    x"3F7E614E",
    x"3F7E6203",
    x"3F7E62B7",
    x"3F7E636C",
    x"3F7E6420",
    x"3F7E64D4",
    x"3F7E6588",
    x"3F7E663B",
    x"3F7E66EF",
    x"3F7E67A2",
    x"3F7E6855",
    x"3F7E6908",
    x"3F7E69BB",
    x"3F7E6A6E",
    x"3F7E6B21",
    x"3F7E6BD3",
    x"3F7E6C85",
    x"3F7E6D38",
    x"3F7E6DEA",
    x"3F7E6E9B",
    x"3F7E6F4D",
    x"3F7E6FFF",
    x"3F7E70B0",
    x"3F7E7161",
    x"3F7E7212",
    x"3F7E72C3",
    x"3F7E7374",
    x"3F7E7424",
    x"3F7E74D5",
    x"3F7E7585",
    x"3F7E7635",
    x"3F7E76E5",
    x"3F7E7795",
    x"3F7E7845",
    x"3F7E78F4",
    x"3F7E79A4",
    x"3F7E7A53",
    x"3F7E7B02",
    x"3F7E7BB1",
    x"3F7E7C60",
    x"3F7E7D0E",
    x"3F7E7DBD",
    x"3F7E7E6B",
    x"3F7E7F19",
    x"3F7E7FC7",
    x"3F7E8075",
    x"3F7E8123",
    x"3F7E81D0",
    x"3F7E827E",
    x"3F7E832B",
    x"3F7E83D8",
    x"3F7E8485",
    x"3F7E8532",
    x"3F7E85DE",
    x"3F7E868B",
    x"3F7E8737",
    x"3F7E87E3",
    x"3F7E888F",
    x"3F7E893B",
    x"3F7E89E7",
    x"3F7E8A92",
    x"3F7E8B3E",
    x"3F7E8BE9",
    x"3F7E8C94",
    x"3F7E8D3F",
    x"3F7E8DEA",
    x"3F7E8E94",
    x"3F7E8F3F",
    x"3F7E8FE9",
    x"3F7E9093",
    x"3F7E913D",
    x"3F7E91E7",
    x"3F7E9291",
    x"3F7E933A",
    x"3F7E93E4",
    x"3F7E948D",
    x"3F7E9536",
    x"3F7E95DF",
    x"3F7E9688",
    x"3F7E9731",
    x"3F7E97D9",
    x"3F7E9881",
    x"3F7E9929",
    x"3F7E99D2",
    x"3F7E9A79",
    x"3F7E9B21",
    x"3F7E9BC9",
    x"3F7E9C70",
    x"3F7E9D17",
    x"3F7E9DBE",
    x"3F7E9E65",
    x"3F7E9F0C",
    x"3F7E9FB3",
    x"3F7EA059",
    x"3F7EA100",
    x"3F7EA1A6",
    x"3F7EA24C",
    x"3F7EA2F2",
    x"3F7EA397",
    x"3F7EA43D",
    x"3F7EA4E2",
    x"3F7EA588",
    x"3F7EA62D",
    x"3F7EA6D2",
    x"3F7EA776",
    x"3F7EA81B",
    x"3F7EA8C0",
    x"3F7EA964",
    x"3F7EAA08",
    x"3F7EAAAC",
    x"3F7EAB50",
    x"3F7EABF4",
    x"3F7EAC97",
    x"3F7EAD3B",
    x"3F7EADDE",
    x"3F7EAE81",
    x"3F7EAF24",
    x"3F7EAFC7",
    x"3F7EB069",
    x"3F7EB10C",
    x"3F7EB1AE",
    x"3F7EB250",
    x"3F7EB2F2",
    x"3F7EB394",
    x"3F7EB436",
    x"3F7EB4D8",
    x"3F7EB579",
    x"3F7EB61A",
    x"3F7EB6BB",
    x"3F7EB75C",
    x"3F7EB7FD",
    x"3F7EB89E",
    x"3F7EB93E",
    x"3F7EB9DF",
    x"3F7EBA7F",
    x"3F7EBB1F",
    x"3F7EBBBF",
    x"3F7EBC5F",
    x"3F7EBCFE",
    x"3F7EBD9E",
    x"3F7EBE3D",
    x"3F7EBEDC",
    x"3F7EBF7B",
    x"3F7EC01A",
    x"3F7EC0B8",
    x"3F7EC157",
    x"3F7EC1F5",
    x"3F7EC293",
    x"3F7EC331",
    x"3F7EC3CF",
    x"3F7EC46D",
    x"3F7EC50B",
    x"3F7EC5A8",
    x"3F7EC645",
    x"3F7EC6E3",
    x"3F7EC780",
    x"3F7EC81C",
    x"3F7EC8B9",
    x"3F7EC955",
    x"3F7EC9F2",
    x"3F7ECA8E",
    x"3F7ECB2A",
    x"3F7ECBC6",
    x"3F7ECC62",
    x"3F7ECCFD",
    x"3F7ECD99",
    x"3F7ECE34",
    x"3F7ECECF",
    x"3F7ECF6A",
    x"3F7ED005",
    x"3F7ED0A0",
    x"3F7ED13A",
    x"3F7ED1D4",
    x"3F7ED26F",
    x"3F7ED309",
    x"3F7ED3A3",
    x"3F7ED43C",
    x"3F7ED4D6",
    x"3F7ED56F",
    x"3F7ED609",
    x"3F7ED6A2",
    x"3F7ED73B",
    x"3F7ED7D4",
    x"3F7ED86C",
    x"3F7ED905",
    x"3F7ED99D",
    x"3F7EDA35",
    x"3F7EDACD",
    x"3F7EDB65",
    x"3F7EDBFD",
    x"3F7EDC95",
    x"3F7EDD2C",
    x"3F7EDDC3",
    x"3F7EDE5B",
    x"3F7EDEF2",
    x"3F7EDF88",
    x"3F7EE01F",
    x"3F7EE0B6",
    x"3F7EE14C",
    x"3F7EE1E2",
    x"3F7EE278",
    x"3F7EE30E",
    x"3F7EE3A4",
    x"3F7EE43A",
    x"3F7EE4CF",
    x"3F7EE564",
    x"3F7EE5F9",
    x"3F7EE68E",
    x"3F7EE723",
    x"3F7EE7B8",
    x"3F7EE84C",
    x"3F7EE8E1",
    x"3F7EE975",
    x"3F7EEA09",
    x"3F7EEA9D",
    x"3F7EEB31",
    x"3F7EEBC4",
    x"3F7EEC58",
    x"3F7EECEB",
    x"3F7EED7E",
    x"3F7EEE11",
    x"3F7EEEA4",
    x"3F7EEF37",
    x"3F7EEFC9",
    x"3F7EF05C",
    x"3F7EF0EE",
    x"3F7EF180",
    x"3F7EF212",
    x"3F7EF2A4",
    x"3F7EF335",
    x"3F7EF3C7",
    x"3F7EF458",
    x"3F7EF4E9",
    x"3F7EF57A",
    x"3F7EF60B",
    x"3F7EF69C",
    x"3F7EF72C",
    x"3F7EF7BD",
    x"3F7EF84D",
    x"3F7EF8DD",
    x"3F7EF96D",
    x"3F7EF9FD",
    x"3F7EFA8C",
    x"3F7EFB1C",
    x"3F7EFBAB",
    x"3F7EFC3A",
    x"3F7EFCC9",
    x"3F7EFD58",
    x"3F7EFDE7",
    x"3F7EFE75",
    x"3F7EFF04",
    x"3F7EFF92",
    x"3F7F0020",
    x"3F7F00AE",
    x"3F7F013C",
    x"3F7F01C9",
    x"3F7F0257",
    x"3F7F02E4",
    x"3F7F0371",
    x"3F7F03FE",
    x"3F7F048B",
    x"3F7F0518",
    x"3F7F05A4",
    x"3F7F0631",
    x"3F7F06BD",
    x"3F7F0749",
    x"3F7F07D5",
    x"3F7F0861",
    x"3F7F08EC",
    x"3F7F0978",
    x"3F7F0A03",
    x"3F7F0A8E",
    x"3F7F0B19",
    x"3F7F0BA4",
    x"3F7F0C2F",
    x"3F7F0CB9",
    x"3F7F0D44",
    x"3F7F0DCE",
    x"3F7F0E58",
    x"3F7F0EE2",
    x"3F7F0F6C",
    x"3F7F0FF5",
    x"3F7F107F",
    x"3F7F1108",
    x"3F7F1191",
    x"3F7F121A",
    x"3F7F12A3",
    x"3F7F132C",
    x"3F7F13B4",
    x"3F7F143D",
    x"3F7F14C5",
    x"3F7F154D",
    x"3F7F15D5",
    x"3F7F165D",
    x"3F7F16E4",
    x"3F7F176C",
    x"3F7F17F3",
    x"3F7F187A",
    x"3F7F1901",
    x"3F7F1988",
    x"3F7F1A0F",
    x"3F7F1A95",
    x"3F7F1B1C",
    x"3F7F1BA2",
    x"3F7F1C28",
    x"3F7F1CAE",
    x"3F7F1D34",
    x"3F7F1DB9",
    x"3F7F1E3F",
    x"3F7F1EC4",
    x"3F7F1F49",
    x"3F7F1FCE",
    x"3F7F2053",
    x"3F7F20D8",
    x"3F7F215C",
    x"3F7F21E1",
    x"3F7F2265",
    x"3F7F22E9",
    x"3F7F236D",
    x"3F7F23F1",
    x"3F7F2475",
    x"3F7F24F8",
    x"3F7F257B",
    x"3F7F25FF",
    x"3F7F2682",
    x"3F7F2704",
    x"3F7F2787",
    x"3F7F280A",
    x"3F7F288C",
    x"3F7F290E",
    x"3F7F2990",
    x"3F7F2A12",
    x"3F7F2A94",
    x"3F7F2B16",
    x"3F7F2B97",
    x"3F7F2C19",
    x"3F7F2C9A",
    x"3F7F2D1B",
    x"3F7F2D9C",
    x"3F7F2E1C",
    x"3F7F2E9D",
    x"3F7F2F1D",
    x"3F7F2F9D",
    x"3F7F301E",
    x"3F7F309E",
    x"3F7F311D",
    x"3F7F319D",
    x"3F7F321C",
    x"3F7F329C",
    x"3F7F331B",
    x"3F7F339A",
    x"3F7F3419",
    x"3F7F3497",
    x"3F7F3516",
    x"3F7F3594",
    x"3F7F3613",
    x"3F7F3691",
    x"3F7F370F",
    x"3F7F378C",
    x"3F7F380A",
    x"3F7F3888",
    x"3F7F3905",
    x"3F7F3982",
    x"3F7F39FF",
    x"3F7F3A7C",
    x"3F7F3AF9",
    x"3F7F3B75",
    x"3F7F3BF2",
    x"3F7F3C6E",
    x"3F7F3CEA",
    x"3F7F3D66",
    x"3F7F3DE2",
    x"3F7F3E5D",
    x"3F7F3ED9",
    x"3F7F3F54",
    x"3F7F3FCF",
    x"3F7F404A",
    x"3F7F40C5",
    x"3F7F4140",
    x"3F7F41BA",
    x"3F7F4235",
    x"3F7F42AF",
    x"3F7F4329",
    x"3F7F43A3",
    x"3F7F441D",
    x"3F7F4497",
    x"3F7F4510",
    x"3F7F4589",
    x"3F7F4603",
    x"3F7F467C",
    x"3F7F46F4",
    x"3F7F476D",
    x"3F7F47E6",
    x"3F7F485E",
    x"3F7F48D6",
    x"3F7F494E",
    x"3F7F49C6",
    x"3F7F4A3E",
    x"3F7F4AB6",
    x"3F7F4B2D",
    x"3F7F4BA5",
    x"3F7F4C1C",
    x"3F7F4C93",
    x"3F7F4D0A",
    x"3F7F4D80",
    x"3F7F4DF7",
    x"3F7F4E6D",
    x"3F7F4EE4",
    x"3F7F4F5A",
    x"3F7F4FD0",
    x"3F7F5045",
    x"3F7F50BB",
    x"3F7F5131",
    x"3F7F51A6",
    x"3F7F521B",
    x"3F7F5290",
    x"3F7F5305",
    x"3F7F537A",
    x"3F7F53EE",
    x"3F7F5463",
    x"3F7F54D7",
    x"3F7F554B",
    x"3F7F55BF",
    x"3F7F5633",
    x"3F7F56A6",
    x"3F7F571A",
    x"3F7F578D",
    x"3F7F5800",
    x"3F7F5873",
    x"3F7F58E6",
    x"3F7F5959",
    x"3F7F59CC",
    x"3F7F5A3E",
    x"3F7F5AB0",
    x"3F7F5B22",
    x"3F7F5B94",
    x"3F7F5C06",
    x"3F7F5C78",
    x"3F7F5CE9",
    x"3F7F5D5A",
    x"3F7F5DCC",
    x"3F7F5E3D",
    x"3F7F5EAE",
    x"3F7F5F1E",
    x"3F7F5F8F",
    x"3F7F5FFF",
    x"3F7F606F",
    x"3F7F60E0",
    x"3F7F6150",
    x"3F7F61BF",
    x"3F7F622F",
    x"3F7F629E",
    x"3F7F630E",
    x"3F7F637D",
    x"3F7F63EC",
    x"3F7F645B",
    x"3F7F64CA",
    x"3F7F6538",
    x"3F7F65A7",
    x"3F7F6615",
    x"3F7F6683",
    x"3F7F66F1",
    x"3F7F675F",
    x"3F7F67CC",
    x"3F7F683A",
    x"3F7F68A7",
    x"3F7F6914",
    x"3F7F6981",
    x"3F7F69EE",
    x"3F7F6A5B",
    x"3F7F6AC7",
    x"3F7F6B34",
    x"3F7F6BA0",
    x"3F7F6C0C",
    x"3F7F6C78",
    x"3F7F6CE4",
    x"3F7F6D50",
    x"3F7F6DBB",
    x"3F7F6E26",
    x"3F7F6E92",
    x"3F7F6EFD",
    x"3F7F6F67",
    x"3F7F6FD2",
    x"3F7F703D",
    x"3F7F70A7",
    x"3F7F7111",
    x"3F7F717B",
    x"3F7F71E5",
    x"3F7F724F",
    x"3F7F72B9",
    x"3F7F7322",
    x"3F7F738C",
    x"3F7F73F5",
    x"3F7F745E",
    x"3F7F74C7",
    x"3F7F752F",
    x"3F7F7598",
    x"3F7F7600",
    x"3F7F7669",
    x"3F7F76D1",
    x"3F7F7739",
    x"3F7F77A0",
    x"3F7F7808",
    x"3F7F7870",
    x"3F7F78D7",
    x"3F7F793E",
    x"3F7F79A5",
    x"3F7F7A0C",
    x"3F7F7A73",
    x"3F7F7AD9",
    x"3F7F7B40",
    x"3F7F7BA6",
    x"3F7F7C0C",
    x"3F7F7C72",
    x"3F7F7CD8",
    x"3F7F7D3D",
    x"3F7F7DA3",
    x"3F7F7E08",
    x"3F7F7E6D",
    x"3F7F7ED2",
    x"3F7F7F37",
    x"3F7F7F9C",
    x"3F7F8000",
    x"3F7F8065",
    x"3F7F80C9",
    x"3F7F812D",
    x"3F7F8191",
    x"3F7F81F5",
    x"3F7F8259",
    x"3F7F82BC",
    x"3F7F831F",
    x"3F7F8383",
    x"3F7F83E6",
    x"3F7F8448",
    x"3F7F84AB",
    x"3F7F850E",
    x"3F7F8570",
    x"3F7F85D2",
    x"3F7F8634",
    x"3F7F8696",
    x"3F7F86F8",
    x"3F7F875A",
    x"3F7F87BB",
    x"3F7F881D",
    x"3F7F887E",
    x"3F7F88DF",
    x"3F7F8940",
    x"3F7F89A0",
    x"3F7F8A01",
    x"3F7F8A61",
    x"3F7F8AC2",
    x"3F7F8B22",
    x"3F7F8B82",
    x"3F7F8BE1",
    x"3F7F8C41",
    x"3F7F8CA1",
    x"3F7F8D00",
    x"3F7F8D5F",
    x"3F7F8DBE",
    x"3F7F8E1D",
    x"3F7F8E7C",
    x"3F7F8EDA",
    x"3F7F8F39",
    x"3F7F8F97",
    x"3F7F8FF5",
    x"3F7F9053",
    x"3F7F90B1",
    x"3F7F910E",
    x"3F7F916C",
    x"3F7F91C9",
    x"3F7F9226",
    x"3F7F9283",
    x"3F7F92E0",
    x"3F7F933D",
    x"3F7F9399",
    x"3F7F93F6",
    x"3F7F9452",
    x"3F7F94AE",
    x"3F7F950A",
    x"3F7F9566",
    x"3F7F95C1",
    x"3F7F961D",
    x"3F7F9678",
    x"3F7F96D3",
    x"3F7F972E",
    x"3F7F9789",
    x"3F7F97E4",
    x"3F7F983F",
    x"3F7F9899",
    x"3F7F98F3",
    x"3F7F994D",
    x"3F7F99A7",
    x"3F7F9A01",
    x"3F7F9A5B",
    x"3F7F9AB4",
    x"3F7F9B0D",
    x"3F7F9B67",
    x"3F7F9BC0",
    x"3F7F9C18",
    x"3F7F9C71",
    x"3F7F9CCA",
    x"3F7F9D22",
    x"3F7F9D7A",
    x"3F7F9DD2",
    x"3F7F9E2A",
    x"3F7F9E82",
    x"3F7F9EDA",
    x"3F7F9F31",
    x"3F7F9F89",
    x"3F7F9FE0",
    x"3F7FA037",
    x"3F7FA08E",
    x"3F7FA0E4",
    x"3F7FA13B",
    x"3F7FA191",
    x"3F7FA1E8",
    x"3F7FA23E",
    x"3F7FA294",
    x"3F7FA2E9",
    x"3F7FA33F",
    x"3F7FA394",
    x"3F7FA3EA",
    x"3F7FA43F",
    x"3F7FA494",
    x"3F7FA4E9",
    x"3F7FA53D",
    x"3F7FA592",
    x"3F7FA5E6",
    x"3F7FA63B",
    x"3F7FA68F",
    x"3F7FA6E3",
    x"3F7FA736",
    x"3F7FA78A",
    x"3F7FA7DE",
    x"3F7FA831",
    x"3F7FA884",
    x"3F7FA8D7",
    x"3F7FA92A",
    x"3F7FA97D",
    x"3F7FA9CF",
    x"3F7FAA21",
    x"3F7FAA74",
    x"3F7FAAC6",
    x"3F7FAB18",
    x"3F7FAB6A",
    x"3F7FABBB",
    x"3F7FAC0D",
    x"3F7FAC5E",
    x"3F7FACAF",
    x"3F7FAD00",
    x"3F7FAD51",
    x"3F7FADA2",
    x"3F7FADF2",
    x"3F7FAE43",
    x"3F7FAE93",
    x"3F7FAEE3",
    x"3F7FAF33",
    x"3F7FAF83",
    x"3F7FAFD2",
    x"3F7FB022",
    x"3F7FB071",
    x"3F7FB0C0",
    x"3F7FB10F",
    x"3F7FB15E",
    x"3F7FB1AD",
    x"3F7FB1FB",
    x"3F7FB24A",
    x"3F7FB298",
    x"3F7FB2E6",
    x"3F7FB334",
    x"3F7FB382",
    x"3F7FB3CF",
    x"3F7FB41D",
    x"3F7FB46A",
    x"3F7FB4B7",
    x"3F7FB504",
    x"3F7FB551",
    x"3F7FB59E",
    x"3F7FB5EA",
    x"3F7FB637",
    x"3F7FB683",
    x"3F7FB6CF",
    x"3F7FB71B",
    x"3F7FB767",
    x"3F7FB7B2",
    x"3F7FB7FE",
    x"3F7FB849",
    x"3F7FB894",
    x"3F7FB8DF",
    x"3F7FB92A",
    x"3F7FB975",
    x"3F7FB9BF",
    x"3F7FBA0A",
    x"3F7FBA54",
    x"3F7FBA9E",
    x"3F7FBAE8",
    x"3F7FBB32",
    x"3F7FBB7B",
    x"3F7FBBC5",
    x"3F7FBC0E",
    x"3F7FBC57",
    x"3F7FBCA0",
    x"3F7FBCE9",
    x"3F7FBD32",
    x"3F7FBD7A",
    x"3F7FBDC2",
    x"3F7FBE0B",
    x"3F7FBE53",
    x"3F7FBE9B",
    x"3F7FBEE2",
    x"3F7FBF2A",
    x"3F7FBF72",
    x"3F7FBFB9",
    x"3F7FC000",
    x"3F7FC047",
    x"3F7FC08E",
    x"3F7FC0D4",
    x"3F7FC11B",
    x"3F7FC161",
    x"3F7FC1A8",
    x"3F7FC1EE",
    x"3F7FC234",
    x"3F7FC279",
    x"3F7FC2BF",
    x"3F7FC304",
    x"3F7FC34A",
    x"3F7FC38F",
    x"3F7FC3D4",
    x"3F7FC419",
    x"3F7FC45D",
    x"3F7FC4A2",
    x"3F7FC4E6",
    x"3F7FC52A",
    x"3F7FC56F",
    x"3F7FC5B2",
    x"3F7FC5F6",
    x"3F7FC63A",
    x"3F7FC67D",
    x"3F7FC6C1",
    x"3F7FC704",
    x"3F7FC747",
    x"3F7FC789",
    x"3F7FC7CC",
    x"3F7FC80F",
    x"3F7FC851",
    x"3F7FC893",
    x"3F7FC8D5",
    x"3F7FC917",
    x"3F7FC959",
    x"3F7FC99B",
    x"3F7FC9DC",
    x"3F7FCA1D",
    x"3F7FCA5E",
    x"3F7FCA9F",
    x"3F7FCAE0",
    x"3F7FCB21",
    x"3F7FCB61",
    x"3F7FCBA2",
    x"3F7FCBE2",
    x"3F7FCC22",
    x"3F7FCC62",
    x"3F7FCCA2",
    x"3F7FCCE1",
    x"3F7FCD21",
    x"3F7FCD60",
    x"3F7FCD9F",
    x"3F7FCDDE",
    x"3F7FCE1D",
    x"3F7FCE5C",
    x"3F7FCE9A",
    x"3F7FCED9",
    x"3F7FCF17",
    x"3F7FCF55",
    x"3F7FCF93",
    x"3F7FCFD1",
    x"3F7FD00E",
    x"3F7FD04C",
    x"3F7FD089",
    x"3F7FD0C6",
    x"3F7FD103",
    x"3F7FD140",
    x"3F7FD17C",
    x"3F7FD1B9",
    x"3F7FD1F5",
    x"3F7FD232",
    x"3F7FD26E",
    x"3F7FD2A9",
    x"3F7FD2E5",
    x"3F7FD321",
    x"3F7FD35C",
    x"3F7FD397",
    x"3F7FD3D3",
    x"3F7FD40E",
    x"3F7FD448",
    x"3F7FD483",
    x"3F7FD4BE",
    x"3F7FD4F8",
    x"3F7FD532",
    x"3F7FD56C",
    x"3F7FD5A6",
    x"3F7FD5E0",
    x"3F7FD619",
    x"3F7FD653",
    x"3F7FD68C",
    x"3F7FD6C5",
    x"3F7FD6FE",
    x"3F7FD737",
    x"3F7FD770",
    x"3F7FD7A8",
    x"3F7FD7E1",
    x"3F7FD819",
    x"3F7FD851",
    x"3F7FD889",
    x"3F7FD8C0",
    x"3F7FD8F8",
    x"3F7FD92F",
    x"3F7FD967",
    x"3F7FD99E",
    x"3F7FD9D5",
    x"3F7FDA0C",
    x"3F7FDA42",
    x"3F7FDA79",
    x"3F7FDAAF",
    x"3F7FDAE5",
    x"3F7FDB1B",
    x"3F7FDB51",
    x"3F7FDB87",
    x"3F7FDBBD",
    x"3F7FDBF2",
    x"3F7FDC27",
    x"3F7FDC5C",
    x"3F7FDC91",
    x"3F7FDCC6",
    x"3F7FDCFB",
    x"3F7FDD2F",
    x"3F7FDD64",
    x"3F7FDD98",
    x"3F7FDDCC",
    x"3F7FDE00",
    x"3F7FDE33",
    x"3F7FDE67",
    x"3F7FDE9A",
    x"3F7FDECE",
    x"3F7FDF01",
    x"3F7FDF34",
    x"3F7FDF67",
    x"3F7FDF99",
    x"3F7FDFCC",
    x"3F7FDFFE",
    x"3F7FE030",
    x"3F7FE062",
    x"3F7FE094",
    x"3F7FE0C6",
    x"3F7FE0F8",
    x"3F7FE129",
    x"3F7FE15A",
    x"3F7FE18B",
    x"3F7FE1BC",
    x"3F7FE1ED",
    x"3F7FE21E",
    x"3F7FE24E",
    x"3F7FE27F",
    x"3F7FE2AF",
    x"3F7FE2DF",
    x"3F7FE30F",
    x"3F7FE33E",
    x"3F7FE36E",
    x"3F7FE39D",
    x"3F7FE3CD",
    x"3F7FE3FC",
    x"3F7FE42B",
    x"3F7FE459",
    x"3F7FE488",
    x"3F7FE4B7",
    x"3F7FE4E5",
    x"3F7FE513",
    x"3F7FE541",
    x"3F7FE56F",
    x"3F7FE59D",
    x"3F7FE5CA",
    x"3F7FE5F8",
    x"3F7FE625",
    x"3F7FE652",
    x"3F7FE67F",
    x"3F7FE6AC",
    x"3F7FE6D8",
    x"3F7FE705",
    x"3F7FE731",
    x"3F7FE75D",
    x"3F7FE789",
    x"3F7FE7B5",
    x"3F7FE7E1",
    x"3F7FE80D",
    x"3F7FE838",
    x"3F7FE863",
    x"3F7FE88E",
    x"3F7FE8B9",
    x"3F7FE8E4",
    x"3F7FE90F",
    x"3F7FE939",
    x"3F7FE964",
    x"3F7FE98E",
    x"3F7FE9B8",
    x"3F7FE9E2",
    x"3F7FEA0B",
    x"3F7FEA35",
    x"3F7FEA5E",
    x"3F7FEA87",
    x"3F7FEAB1",
    x"3F7FEADA",
    x"3F7FEB02",
    x"3F7FEB2B",
    x"3F7FEB53",
    x"3F7FEB7C",
    x"3F7FEBA4",
    x"3F7FEBCC",
    x"3F7FEBF4",
    x"3F7FEC1B",
    x"3F7FEC43",
    x"3F7FEC6A",
    x"3F7FEC92",
    x"3F7FECB9",
    x"3F7FECE0",
    x"3F7FED06",
    x"3F7FED2D",
    x"3F7FED54",
    x"3F7FED7A",
    x"3F7FEDA0",
    x"3F7FEDC6",
    x"3F7FEDEC",
    x"3F7FEE12",
    x"3F7FEE37",
    x"3F7FEE5D",
    x"3F7FEE82",
    x"3F7FEEA7",
    x"3F7FEECC",
    x"3F7FEEF1",
    x"3F7FEF15",
    x"3F7FEF3A",
    x"3F7FEF5E",
    x"3F7FEF82",
    x"3F7FEFA6",
    x"3F7FEFCA",
    x"3F7FEFEE",
    x"3F7FF011",
    x"3F7FF035",
    x"3F7FF058",
    x"3F7FF07B",
    x"3F7FF09E",
    x"3F7FF0C1",
    x"3F7FF0E3",
    x"3F7FF106",
    x"3F7FF128",
    x"3F7FF14A",
    x"3F7FF16C",
    x"3F7FF18E",
    x"3F7FF1B0",
    x"3F7FF1D1",
    x"3F7FF1F3",
    x"3F7FF214",
    x"3F7FF235",
    x"3F7FF256",
    x"3F7FF277",
    x"3F7FF297",
    x"3F7FF2B8",
    x"3F7FF2D8",
    x"3F7FF2F8",
    x"3F7FF318",
    x"3F7FF338",
    x"3F7FF358",
    x"3F7FF377",
    x"3F7FF397",
    x"3F7FF3B6",
    x"3F7FF3D5",
    x"3F7FF3F4",
    x"3F7FF413",
    x"3F7FF431",
    x"3F7FF450",
    x"3F7FF46E",
    x"3F7FF48C",
    x"3F7FF4AA",
    x"3F7FF4C8",
    x"3F7FF4E6",
    x"3F7FF503",
    x"3F7FF521",
    x"3F7FF53E",
    x"3F7FF55B",
    x"3F7FF578",
    x"3F7FF595",
    x"3F7FF5B1",
    x"3F7FF5CE",
    x"3F7FF5EA",
    x"3F7FF606",
    x"3F7FF622",
    x"3F7FF63E",
    x"3F7FF659",
    x"3F7FF675",
    x"3F7FF690",
    x"3F7FF6AC",
    x"3F7FF6C7",
    x"3F7FF6E2",
    x"3F7FF6FC",
    x"3F7FF717",
    x"3F7FF731",
    x"3F7FF74C",
    x"3F7FF766",
    x"3F7FF780",
    x"3F7FF79A",
    x"3F7FF7B3",
    x"3F7FF7CD",
    x"3F7FF7E6",
    x"3F7FF7FF",
    x"3F7FF818",
    x"3F7FF831",
    x"3F7FF84A",
    x"3F7FF863",
    x"3F7FF87B",
    x"3F7FF893",
    x"3F7FF8AC",
    x"3F7FF8C4",
    x"3F7FF8DB",
    x"3F7FF8F3",
    x"3F7FF90B",
    x"3F7FF922",
    x"3F7FF939",
    x"3F7FF950",
    x"3F7FF967",
    x"3F7FF97E",
    x"3F7FF994",
    x"3F7FF9AB",
    x"3F7FF9C1",
    x"3F7FF9D7",
    x"3F7FF9ED",
    x"3F7FFA03",
    x"3F7FFA19",
    x"3F7FFA2E",
    x"3F7FFA44",
    x"3F7FFA59",
    x"3F7FFA6E",
    x"3F7FFA83",
    x"3F7FFA97",
    x"3F7FFAAC",
    x"3F7FFAC1",
    x"3F7FFAD5",
    x"3F7FFAE9",
    x"3F7FFAFD",
    x"3F7FFB11",
    x"3F7FFB24",
    x"3F7FFB38",
    x"3F7FFB4B",
    x"3F7FFB5E",
    x"3F7FFB71",
    x"3F7FFB84",
    x"3F7FFB97",
    x"3F7FFBAA",
    x"3F7FFBBC",
    x"3F7FFBCE",
    x"3F7FFBE1",
    x"3F7FFBF2",
    x"3F7FFC04",
    x"3F7FFC16",
    x"3F7FFC27",
    x"3F7FFC39",
    x"3F7FFC4A",
    x"3F7FFC5B",
    x"3F7FFC6C",
    x"3F7FFC7D",
    x"3F7FFC8D",
    x"3F7FFC9E",
    x"3F7FFCAE",
    x"3F7FFCBE",
    x"3F7FFCCE",
    x"3F7FFCDE",
    x"3F7FFCED",
    x"3F7FFCFD",
    x"3F7FFD0C",
    x"3F7FFD1B",
    x"3F7FFD2B",
    x"3F7FFD39",
    x"3F7FFD48",
    x"3F7FFD57",
    x"3F7FFD65",
    x"3F7FFD73",
    x"3F7FFD81",
    x"3F7FFD8F",
    x"3F7FFD9D",
    x"3F7FFDAB",
    x"3F7FFDB8",
    x"3F7FFDC6",
    x"3F7FFDD3",
    x"3F7FFDE0",
    x"3F7FFDED",
    x"3F7FFDFA",
    x"3F7FFE06",
    x"3F7FFE13",
    x"3F7FFE1F",
    x"3F7FFE2B",
    x"3F7FFE37",
    x"3F7FFE43",
    x"3F7FFE4E",
    x"3F7FFE5A",
    x"3F7FFE65",
    x"3F7FFE70",
    x"3F7FFE7B",
    x"3F7FFE86",
    x"3F7FFE91",
    x"3F7FFE9B",
    x"3F7FFEA6",
    x"3F7FFEB0",
    x"3F7FFEBA",
    x"3F7FFEC4",
    x"3F7FFECE",
    x"3F7FFED8",
    x"3F7FFEE1",
    x"3F7FFEEA",
    x"3F7FFEF4",
    x"3F7FFEFD",
    x"3F7FFF05",
    x"3F7FFF0E",
    x"3F7FFF17",
    x"3F7FFF1F",
    x"3F7FFF27",
    x"3F7FFF30",
    x"3F7FFF37",
    x"3F7FFF3F",
    x"3F7FFF47",
    x"3F7FFF4E",
    x"3F7FFF56",
    x"3F7FFF5D",
    x"3F7FFF64",
    x"3F7FFF6B",
    x"3F7FFF71",
    x"3F7FFF78",
    x"3F7FFF7E",
    x"3F7FFF85",
    x"3F7FFF8B",
    x"3F7FFF91",
    x"3F7FFF96",
    x"3F7FFF9C",
    x"3F7FFFA2",
    x"3F7FFFA7",
    x"3F7FFFAC",
    x"3F7FFFB1",
    x"3F7FFFB6",
    x"3F7FFFBB",
    x"3F7FFFBF",
    x"3F7FFFC4",
    x"3F7FFFC8",
    x"3F7FFFCC",
    x"3F7FFFD0",
    x"3F7FFFD4",
    x"3F7FFFD7",
    x"3F7FFFDB",
    x"3F7FFFDE",
    x"3F7FFFE1",
    x"3F7FFFE4",
    x"3F7FFFE7",
    x"3F7FFFEA",
    x"3F7FFFEC",
    x"3F7FFFEF",
    x"3F7FFFF1",
    x"3F7FFFF3",
    x"3F7FFFF5",
    x"3F7FFFF7",
    x"3F7FFFF8",
    x"3F7FFFFA",
    x"3F7FFFFB",
    x"3F7FFFFC",
    x"3F7FFFFD",
    x"3F7FFFFE",
    x"3F7FFFFF",
    x"3F7FFFFF",
    x"3F800000",
    x"3F800000"
  );

begin

  p_mem_read : process (clk) begin
    if rising_edge(clk) then
      data_out <= mem(to_integer(unsigned(address)));
    end if;
  end process;

end architecture;
